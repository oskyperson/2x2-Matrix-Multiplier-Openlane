VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO matrix_multiplier
  CLASS BLOCK ;
  FOREIGN matrix_multiplier ;
  ORIGIN 0.000 0.000 ;
  SIZE 236.440 BY 247.160 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 234.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 234.160 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 234.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 234.160 ;
    END
  END VPWR
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 128.890 243.160 129.170 247.160 ;
    END
  END cs
  PIN hz100
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END hz100
  PIN miso
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 232.440 190.440 236.440 191.040 ;
    END
  END miso
  PIN mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 243.160 116.290 247.160 ;
    END
  END mosi
  PIN ready
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END ready
  PIN spi_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 206.170 243.160 206.450 247.160 ;
    END
  END spi_clk
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 231.110 234.005 ;
      LAYER li1 ;
        RECT 5.520 10.795 230.920 234.005 ;
      LAYER met1 ;
        RECT 0.530 10.640 230.920 234.160 ;
      LAYER met2 ;
        RECT 0.550 242.880 115.730 243.850 ;
        RECT 116.570 242.880 128.610 243.850 ;
        RECT 129.450 242.880 205.890 243.850 ;
        RECT 206.730 242.880 229.910 243.850 ;
        RECT 0.550 4.280 229.910 242.880 ;
        RECT 0.550 4.000 131.830 4.280 ;
        RECT 132.670 4.000 229.910 4.280 ;
      LAYER met3 ;
        RECT 0.525 215.240 232.440 234.085 ;
        RECT 4.400 213.840 232.440 215.240 ;
        RECT 0.525 191.440 232.440 213.840 ;
        RECT 0.525 190.040 232.040 191.440 ;
        RECT 0.525 10.715 232.440 190.040 ;
      LAYER met4 ;
        RECT 65.615 47.775 174.240 210.625 ;
        RECT 176.640 47.775 177.540 210.625 ;
        RECT 179.940 47.775 226.945 210.625 ;
  END
END matrix_multiplier
END LIBRARY


magic
tech sky130A
magscale 1 2
timestamp 1726721562
<< viali >>
rect 13001 28713 13035 28747
rect 13553 28713 13587 28747
rect 14381 28713 14415 28747
rect 15025 28713 15059 28747
rect 15669 28713 15703 28747
rect 16773 28713 16807 28747
rect 17877 28713 17911 28747
rect 18521 28713 18555 28747
rect 19901 28713 19935 28747
rect 21097 28713 21131 28747
rect 23121 28713 23155 28747
rect 23673 28713 23707 28747
rect 24593 28713 24627 28747
rect 25697 28713 25731 28747
rect 26157 28713 26191 28747
rect 27169 28713 27203 28747
rect 17509 28645 17543 28679
rect 19533 28645 19567 28679
rect 20729 28645 20763 28679
rect 22109 28645 22143 28679
rect 22661 28645 22695 28679
rect 25237 28645 25271 28679
rect 15301 28509 15335 28543
rect 17325 28509 17359 28543
rect 27077 28509 27111 28543
rect 13277 28441 13311 28475
rect 13829 28441 13863 28475
rect 14657 28441 14691 28475
rect 15945 28441 15979 28475
rect 17049 28441 17083 28475
rect 18153 28441 18187 28475
rect 18429 28441 18463 28475
rect 19349 28441 19383 28475
rect 20177 28441 20211 28475
rect 20453 28441 20487 28475
rect 21005 28441 21039 28475
rect 21925 28441 21959 28475
rect 22477 28441 22511 28475
rect 23029 28441 23063 28475
rect 23581 28441 23615 28475
rect 24501 28441 24535 28475
rect 25053 28441 25087 28475
rect 25605 28441 25639 28475
rect 26433 28441 26467 28475
rect 18061 28169 18095 28203
rect 19073 28169 19107 28203
rect 20085 28169 20119 28203
rect 20177 28169 20211 28203
rect 22385 28169 22419 28203
rect 27353 28169 27387 28203
rect 19241 28101 19275 28135
rect 19441 28101 19475 28135
rect 19533 28101 19567 28135
rect 20329 28101 20363 28135
rect 20545 28101 20579 28135
rect 22201 28101 22235 28135
rect 25973 28101 26007 28135
rect 27261 28101 27295 28135
rect 6837 28033 6871 28067
rect 7021 28033 7055 28067
rect 10977 28033 11011 28067
rect 11804 28033 11838 28067
rect 11897 28033 11931 28067
rect 17969 28033 18003 28067
rect 18153 28033 18187 28067
rect 19717 28033 19751 28067
rect 19809 28033 19843 28067
rect 19901 28033 19935 28067
rect 21097 28033 21131 28067
rect 21189 28033 21223 28067
rect 22017 28033 22051 28067
rect 22109 28033 22143 28067
rect 24685 28033 24719 28067
rect 25145 28033 25179 28067
rect 25881 28033 25915 28067
rect 26065 28033 26099 28067
rect 26433 28033 26467 28067
rect 26801 28033 26835 28067
rect 11253 27965 11287 27999
rect 25053 27965 25087 27999
rect 21833 27897 21867 27931
rect 7021 27829 7055 27863
rect 10793 27829 10827 27863
rect 11161 27829 11195 27863
rect 11713 27829 11747 27863
rect 19257 27829 19291 27863
rect 20361 27829 20395 27863
rect 24869 27829 24903 27863
rect 25329 27829 25363 27863
rect 5641 27625 5675 27659
rect 10425 27625 10459 27659
rect 11069 27625 11103 27659
rect 17233 27625 17267 27659
rect 18245 27625 18279 27659
rect 18981 27625 19015 27659
rect 19441 27625 19475 27659
rect 20821 27625 20855 27659
rect 21281 27625 21315 27659
rect 21925 27625 21959 27659
rect 22109 27625 22143 27659
rect 23489 27625 23523 27659
rect 24869 27625 24903 27659
rect 25145 27625 25179 27659
rect 25697 27625 25731 27659
rect 26341 27625 26375 27659
rect 10333 27557 10367 27591
rect 17509 27557 17543 27591
rect 17785 27557 17819 27591
rect 19257 27557 19291 27591
rect 19993 27557 20027 27591
rect 21465 27557 21499 27591
rect 23029 27557 23063 27591
rect 24225 27557 24259 27591
rect 27721 27557 27755 27591
rect 5089 27489 5123 27523
rect 7021 27489 7055 27523
rect 7389 27489 7423 27523
rect 9689 27489 9723 27523
rect 9965 27489 9999 27523
rect 10793 27489 10827 27523
rect 19533 27489 19567 27523
rect 22753 27489 22787 27523
rect 3801 27421 3835 27455
rect 3985 27421 4019 27455
rect 4997 27421 5031 27455
rect 6101 27421 6135 27455
rect 6285 27421 6319 27455
rect 6469 27421 6503 27455
rect 6653 27421 6687 27455
rect 6929 27421 6963 27455
rect 7573 27421 7607 27455
rect 7849 27421 7883 27455
rect 8033 27421 8067 27455
rect 9597 27421 9631 27455
rect 10609 27421 10643 27455
rect 10701 27421 10735 27455
rect 10885 27421 10919 27455
rect 11161 27421 11195 27455
rect 11345 27421 11379 27455
rect 11529 27421 11563 27455
rect 11805 27421 11839 27455
rect 11897 27421 11931 27455
rect 12081 27421 12115 27455
rect 12295 27421 12329 27455
rect 12449 27421 12483 27455
rect 17233 27421 17267 27455
rect 17417 27421 17451 27455
rect 17509 27421 17543 27455
rect 17693 27421 17727 27455
rect 17785 27421 17819 27455
rect 17969 27421 18003 27455
rect 18061 27421 18095 27455
rect 18245 27421 18279 27455
rect 18613 27421 18647 27455
rect 18797 27421 18831 27455
rect 19073 27421 19107 27455
rect 19441 27421 19475 27455
rect 20269 27421 20303 27455
rect 20637 27421 20671 27455
rect 20821 27421 20855 27455
rect 20913 27421 20947 27455
rect 21557 27421 21591 27455
rect 22385 27421 22419 27455
rect 23213 27421 23247 27455
rect 23305 27421 23339 27455
rect 24041 27421 24075 27455
rect 24225 27421 24259 27455
rect 24501 27421 24535 27455
rect 24593 27421 24627 27455
rect 24961 27421 24995 27455
rect 25329 27421 25363 27455
rect 25421 27421 25455 27455
rect 25789 27421 25823 27455
rect 26065 27421 26099 27455
rect 26249 27421 26283 27455
rect 26341 27421 26375 27455
rect 26525 27421 26559 27455
rect 27445 27421 27479 27455
rect 5457 27353 5491 27387
rect 12541 27353 12575 27387
rect 12725 27353 12759 27387
rect 12909 27353 12943 27387
rect 19901 27353 19935 27387
rect 20545 27353 20579 27387
rect 21925 27353 21959 27387
rect 22870 27353 22904 27387
rect 26893 27353 26927 27387
rect 27261 27353 27295 27387
rect 3893 27285 3927 27319
rect 5365 27285 5399 27319
rect 5657 27285 5691 27319
rect 5825 27285 5859 27319
rect 6101 27285 6135 27319
rect 6561 27285 6595 27319
rect 7297 27285 7331 27319
rect 9229 27285 9263 27319
rect 18429 27285 18463 27319
rect 20177 27285 20211 27319
rect 20361 27285 20395 27319
rect 21281 27285 21315 27319
rect 22661 27285 22695 27319
rect 25973 27285 26007 27319
rect 26157 27285 26191 27319
rect 3525 27081 3559 27115
rect 5273 27081 5307 27115
rect 6377 27081 6411 27115
rect 7941 27081 7975 27115
rect 10701 27081 10735 27115
rect 11529 27081 11563 27115
rect 12173 27081 12207 27115
rect 17877 27081 17911 27115
rect 18337 27081 18371 27115
rect 20269 27081 20303 27115
rect 22017 27081 22051 27115
rect 22201 27081 22235 27115
rect 24869 27081 24903 27115
rect 25053 27081 25087 27115
rect 25789 27081 25823 27115
rect 26065 27081 26099 27115
rect 26341 27081 26375 27115
rect 3157 27013 3191 27047
rect 3357 27013 3391 27047
rect 3893 27013 3927 27047
rect 7297 27013 7331 27047
rect 11161 27013 11195 27047
rect 12325 27013 12359 27047
rect 12541 27013 12575 27047
rect 12817 27013 12851 27047
rect 18889 27013 18923 27047
rect 19901 27013 19935 27047
rect 21189 27013 21223 27047
rect 22753 27013 22787 27047
rect 22937 27013 22971 27047
rect 23153 27013 23187 27047
rect 23397 27013 23431 27047
rect 23581 27013 23615 27047
rect 2421 26945 2455 26979
rect 3617 26945 3651 26979
rect 3709 26945 3743 26979
rect 4077 26945 4111 26979
rect 4445 26945 4479 26979
rect 5181 26945 5215 26979
rect 5365 26945 5399 26979
rect 5548 26945 5582 26979
rect 6561 26945 6595 26979
rect 6653 26945 6687 26979
rect 6929 26945 6963 26979
rect 7389 26945 7423 26979
rect 7481 26945 7515 26979
rect 7757 26945 7791 26979
rect 8033 26945 8067 26979
rect 8217 26945 8251 26979
rect 10057 26945 10091 26979
rect 10977 26945 11011 26979
rect 11253 26945 11287 26979
rect 11713 26945 11747 26979
rect 12081 26945 12115 26979
rect 12633 26945 12667 26979
rect 17785 26945 17819 26979
rect 17969 26945 18003 26979
rect 18245 26945 18279 26979
rect 18429 26945 18463 26979
rect 19164 26945 19198 26979
rect 19257 26945 19291 26979
rect 19533 26945 19567 26979
rect 20361 26945 20395 26979
rect 20545 26945 20579 26979
rect 20729 26945 20763 26979
rect 21005 26945 21039 26979
rect 21556 26945 21590 26979
rect 21649 26945 21683 26979
rect 24225 26945 24259 26979
rect 24685 26945 24719 26979
rect 24961 26945 24995 26979
rect 25145 26945 25179 26979
rect 25697 26945 25731 26979
rect 25881 26945 25915 26979
rect 25973 26945 26007 26979
rect 26157 26945 26191 26979
rect 26249 26945 26283 26979
rect 26433 26945 26467 26979
rect 27537 26945 27571 26979
rect 2329 26877 2363 26911
rect 2789 26877 2823 26911
rect 5089 26877 5123 26911
rect 5641 26877 5675 26911
rect 5733 26877 5767 26911
rect 5825 26877 5859 26911
rect 6377 26877 6411 26911
rect 7205 26877 7239 26911
rect 7573 26877 7607 26911
rect 10241 26877 10275 26911
rect 10333 26877 10367 26911
rect 21281 26877 21315 26911
rect 22293 26877 22327 26911
rect 24501 26877 24535 26911
rect 20085 26809 20119 26843
rect 20821 26809 20855 26843
rect 20913 26809 20947 26843
rect 22753 26809 22787 26843
rect 3341 26741 3375 26775
rect 3893 26741 3927 26775
rect 6009 26741 6043 26775
rect 7067 26741 7101 26775
rect 7481 26741 7515 26775
rect 8125 26741 8159 26775
rect 10793 26741 10827 26775
rect 11989 26741 12023 26775
rect 12357 26741 12391 26775
rect 13001 26741 13035 26775
rect 19901 26741 19935 26775
rect 23121 26741 23155 26775
rect 23305 26741 23339 26775
rect 24317 26741 24351 26775
rect 27721 26741 27755 26775
rect 3249 26537 3283 26571
rect 3985 26537 4019 26571
rect 4261 26537 4295 26571
rect 6929 26537 6963 26571
rect 9505 26537 9539 26571
rect 12081 26537 12115 26571
rect 19717 26537 19751 26571
rect 20177 26537 20211 26571
rect 20361 26537 20395 26571
rect 22385 26537 22419 26571
rect 26801 26537 26835 26571
rect 5549 26469 5583 26503
rect 12817 26469 12851 26503
rect 22845 26469 22879 26503
rect 23581 26469 23615 26503
rect 27721 26469 27755 26503
rect 6469 26401 6503 26435
rect 12725 26401 12759 26435
rect 19993 26401 20027 26435
rect 20729 26401 20763 26435
rect 23213 26401 23247 26435
rect 23305 26401 23339 26435
rect 25262 26401 25296 26435
rect 26065 26401 26099 26435
rect 1869 26333 1903 26367
rect 3341 26333 3375 26367
rect 4261 26333 4295 26367
rect 4445 26333 4479 26367
rect 4997 26333 5031 26367
rect 5181 26333 5215 26367
rect 5273 26333 5307 26367
rect 5365 26333 5399 26367
rect 5549 26333 5583 26367
rect 5825 26333 5859 26367
rect 5917 26333 5951 26367
rect 6377 26333 6411 26367
rect 6837 26333 6871 26367
rect 9045 26333 9079 26367
rect 9137 26333 9171 26367
rect 9321 26333 9355 26367
rect 9597 26333 9631 26367
rect 9689 26333 9723 26367
rect 9873 26333 9907 26367
rect 10609 26333 10643 26367
rect 10793 26333 10827 26367
rect 10885 26333 10919 26367
rect 11989 26333 12023 26367
rect 12265 26333 12299 26367
rect 12541 26333 12575 26367
rect 13093 26333 13127 26367
rect 13185 26333 13219 26367
rect 13369 26333 13403 26367
rect 20269 26333 20303 26367
rect 20545 26333 20579 26367
rect 22477 26333 22511 26367
rect 22661 26333 22695 26367
rect 22845 26333 22879 26367
rect 22937 26333 22971 26367
rect 24777 26333 24811 26367
rect 25145 26333 25179 26367
rect 25697 26333 25731 26367
rect 26341 26333 26375 26367
rect 26709 26333 26743 26367
rect 27537 26333 27571 26367
rect 2881 26265 2915 26299
rect 5089 26265 5123 26299
rect 6101 26265 6135 26299
rect 12817 26265 12851 26299
rect 13277 26265 13311 26299
rect 23422 26265 23456 26299
rect 25053 26265 25087 26299
rect 26525 26265 26559 26299
rect 6745 26197 6779 26231
rect 9781 26197 9815 26231
rect 10885 26197 10919 26231
rect 12357 26197 12391 26231
rect 13001 26197 13035 26231
rect 25421 26197 25455 26231
rect 12449 25993 12483 26027
rect 12909 25993 12943 26027
rect 26173 25993 26207 26027
rect 26341 25993 26375 26027
rect 8217 25925 8251 25959
rect 8401 25925 8435 25959
rect 8585 25925 8619 25959
rect 12633 25925 12667 25959
rect 12817 25925 12851 25959
rect 23029 25925 23063 25959
rect 25513 25925 25547 25959
rect 25605 25925 25639 25959
rect 25973 25925 26007 25959
rect 2789 25857 2823 25891
rect 3157 25857 3191 25891
rect 6745 25857 6779 25891
rect 7941 25857 7975 25891
rect 8135 25857 8169 25891
rect 8677 25857 8711 25891
rect 8861 25857 8895 25891
rect 12265 25857 12299 25891
rect 12541 25857 12575 25891
rect 12909 25857 12943 25891
rect 20453 25857 20487 25891
rect 22661 25857 22695 25891
rect 22845 25857 22879 25891
rect 25421 25857 25455 25891
rect 26433 25857 26467 25891
rect 2513 25789 2547 25823
rect 6837 25789 6871 25823
rect 7205 25789 7239 25823
rect 8033 25789 8067 25823
rect 25789 25789 25823 25823
rect 7481 25721 7515 25755
rect 25237 25721 25271 25755
rect 26525 25721 26559 25755
rect 7021 25653 7055 25687
rect 7665 25653 7699 25687
rect 8769 25653 8803 25687
rect 12081 25653 12115 25687
rect 20545 25653 20579 25687
rect 26157 25653 26191 25687
rect 13001 25449 13035 25483
rect 15945 25449 15979 25483
rect 16957 25449 16991 25483
rect 25697 25449 25731 25483
rect 26525 25449 26559 25483
rect 9689 25245 9723 25279
rect 9873 25245 9907 25279
rect 10241 25245 10275 25279
rect 10395 25245 10429 25279
rect 10701 25245 10735 25279
rect 10885 25245 10919 25279
rect 12357 25245 12391 25279
rect 12449 25245 12483 25279
rect 12633 25245 12667 25279
rect 12725 25245 12759 25279
rect 15577 25245 15611 25279
rect 15669 25245 15703 25279
rect 15761 25245 15795 25279
rect 22017 25245 22051 25279
rect 25605 25245 25639 25279
rect 25881 25245 25915 25279
rect 27537 25245 27571 25279
rect 12909 25177 12943 25211
rect 16773 25177 16807 25211
rect 22201 25177 22235 25211
rect 26065 25177 26099 25211
rect 26157 25177 26191 25211
rect 26341 25177 26375 25211
rect 27169 25177 27203 25211
rect 9873 25109 9907 25143
rect 10609 25109 10643 25143
rect 10885 25109 10919 25143
rect 12173 25109 12207 25143
rect 16973 25109 17007 25143
rect 17141 25109 17175 25143
rect 27077 25109 27111 25143
rect 27721 25109 27755 25143
rect 14933 24905 14967 24939
rect 16865 24905 16899 24939
rect 17417 24905 17451 24939
rect 21557 24905 21591 24939
rect 25881 24905 25915 24939
rect 27185 24905 27219 24939
rect 10149 24837 10183 24871
rect 11805 24837 11839 24871
rect 12021 24837 12055 24871
rect 16221 24837 16255 24871
rect 16405 24837 16439 24871
rect 26985 24837 27019 24871
rect 1409 24769 1443 24803
rect 2513 24769 2547 24803
rect 2697 24769 2731 24803
rect 2789 24769 2823 24803
rect 2973 24769 3007 24803
rect 3157 24769 3191 24803
rect 4445 24769 4479 24803
rect 4629 24769 4663 24803
rect 5089 24769 5123 24803
rect 5273 24769 5307 24803
rect 5365 24769 5399 24803
rect 5457 24769 5491 24803
rect 8217 24769 8251 24803
rect 8401 24769 8435 24803
rect 8677 24769 8711 24803
rect 9045 24769 9079 24803
rect 10333 24769 10367 24803
rect 10609 24769 10643 24803
rect 10793 24769 10827 24803
rect 10885 24769 10919 24803
rect 10977 24769 11011 24803
rect 14841 24769 14875 24803
rect 15117 24769 15151 24803
rect 15393 24769 15427 24803
rect 15838 24769 15872 24803
rect 16129 24769 16163 24803
rect 16681 24769 16715 24803
rect 16773 24769 16807 24803
rect 17141 24769 17175 24803
rect 17325 24769 17359 24803
rect 17601 24769 17635 24803
rect 21465 24769 21499 24803
rect 22017 24769 22051 24803
rect 22293 24769 22327 24803
rect 22569 24769 22603 24803
rect 22937 24769 22971 24803
rect 23121 24769 23155 24803
rect 23213 24769 23247 24803
rect 25789 24769 25823 24803
rect 25881 24769 25915 24803
rect 25973 24769 26007 24803
rect 26433 24769 26467 24803
rect 27537 24769 27571 24803
rect 2605 24701 2639 24735
rect 4169 24701 4203 24735
rect 9137 24701 9171 24735
rect 9229 24701 9263 24735
rect 15761 24701 15795 24735
rect 22845 24701 22879 24735
rect 25605 24701 25639 24735
rect 26249 24701 26283 24735
rect 5181 24633 5215 24667
rect 15301 24633 15335 24667
rect 16313 24633 16347 24667
rect 22937 24633 22971 24667
rect 27353 24633 27387 24667
rect 1593 24565 1627 24599
rect 2973 24565 3007 24599
rect 4537 24565 4571 24599
rect 8861 24565 8895 24599
rect 9413 24565 9447 24599
rect 10517 24565 10551 24599
rect 11253 24565 11287 24599
rect 11989 24565 12023 24599
rect 12173 24565 12207 24599
rect 16037 24565 16071 24599
rect 17049 24565 17083 24599
rect 17141 24565 17175 24599
rect 17785 24565 17819 24599
rect 21833 24565 21867 24599
rect 22201 24565 22235 24599
rect 22385 24565 22419 24599
rect 22753 24565 22787 24599
rect 26065 24565 26099 24599
rect 26617 24565 26651 24599
rect 27169 24565 27203 24599
rect 27721 24565 27755 24599
rect 3433 24361 3467 24395
rect 7849 24361 7883 24395
rect 10241 24361 10275 24395
rect 21465 24361 21499 24395
rect 23305 24361 23339 24395
rect 23489 24361 23523 24395
rect 25881 24361 25915 24395
rect 26893 24361 26927 24395
rect 4721 24293 4755 24327
rect 9597 24293 9631 24327
rect 12633 24293 12667 24327
rect 13001 24293 13035 24327
rect 17417 24293 17451 24327
rect 26433 24293 26467 24327
rect 4261 24225 4295 24259
rect 4445 24225 4479 24259
rect 5089 24225 5123 24259
rect 10609 24225 10643 24259
rect 10701 24225 10735 24259
rect 11713 24225 11747 24259
rect 15117 24225 15151 24259
rect 15485 24225 15519 24259
rect 18061 24225 18095 24259
rect 21097 24225 21131 24259
rect 21833 24225 21867 24259
rect 24777 24225 24811 24259
rect 25881 24225 25915 24259
rect 26249 24225 26283 24259
rect 26801 24225 26835 24259
rect 2421 24157 2455 24191
rect 2513 24157 2547 24191
rect 4353 24157 4387 24191
rect 4537 24157 4571 24191
rect 7481 24157 7515 24191
rect 7665 24157 7699 24191
rect 9413 24157 9447 24191
rect 9689 24157 9723 24191
rect 9781 24157 9815 24191
rect 9965 24157 9999 24191
rect 10057 24157 10091 24191
rect 10333 24157 10367 24191
rect 10425 24157 10459 24191
rect 11989 24157 12023 24191
rect 12541 24157 12575 24191
rect 12817 24157 12851 24191
rect 13001 24157 13035 24191
rect 14289 24157 14323 24191
rect 15301 24157 15335 24191
rect 15669 24157 15703 24191
rect 17969 24157 18003 24191
rect 21281 24157 21315 24191
rect 21465 24157 21499 24191
rect 21557 24157 21591 24191
rect 23673 24157 23707 24191
rect 23765 24157 23799 24191
rect 24685 24157 24719 24191
rect 25145 24157 25179 24191
rect 26893 24157 26927 24191
rect 27077 24157 27111 24191
rect 27537 24157 27571 24191
rect 1501 24089 1535 24123
rect 3525 24089 3559 24123
rect 5641 24089 5675 24123
rect 9229 24089 9263 24123
rect 10793 24089 10827 24123
rect 15945 24089 15979 24123
rect 20821 24089 20855 24123
rect 25053 24089 25087 24123
rect 1777 24021 1811 24055
rect 3065 24021 3099 24055
rect 14197 24021 14231 24055
rect 17601 24021 17635 24055
rect 19349 24021 19383 24055
rect 24501 24021 24535 24055
rect 24869 24021 24903 24055
rect 26065 24021 26099 24055
rect 26341 24021 26375 24055
rect 27721 24021 27755 24055
rect 9229 23817 9263 23851
rect 18061 23817 18095 23851
rect 18889 23817 18923 23851
rect 26249 23817 26283 23851
rect 2513 23749 2547 23783
rect 9413 23749 9447 23783
rect 9781 23749 9815 23783
rect 10057 23749 10091 23783
rect 13553 23749 13587 23783
rect 17509 23749 17543 23783
rect 18153 23749 18187 23783
rect 18489 23749 18523 23783
rect 18705 23749 18739 23783
rect 19165 23749 19199 23783
rect 21373 23749 21407 23783
rect 25881 23749 25915 23783
rect 25973 23749 26007 23783
rect 4537 23681 4571 23715
rect 4721 23681 4755 23715
rect 5549 23681 5583 23715
rect 5951 23681 5985 23715
rect 7297 23681 7331 23715
rect 9137 23681 9171 23715
rect 9321 23681 9355 23715
rect 9597 23681 9631 23715
rect 10241 23681 10275 23715
rect 12265 23681 12299 23715
rect 12909 23681 12943 23715
rect 13277 23681 13311 23715
rect 15945 23681 15979 23715
rect 16129 23681 16163 23715
rect 16773 23681 16807 23715
rect 17141 23681 17175 23715
rect 17233 23681 17267 23715
rect 17417 23681 17451 23715
rect 17601 23681 17635 23715
rect 18245 23681 18279 23715
rect 18797 23681 18831 23715
rect 19073 23681 19107 23715
rect 25605 23681 25639 23715
rect 25753 23681 25787 23715
rect 26070 23681 26104 23715
rect 27537 23681 27571 23715
rect 1961 23613 1995 23647
rect 5181 23613 5215 23647
rect 5641 23613 5675 23647
rect 7389 23613 7423 23647
rect 11897 23613 11931 23647
rect 12633 23613 12667 23647
rect 17877 23613 17911 23647
rect 19901 23613 19935 23647
rect 21649 23613 21683 23647
rect 23305 23613 23339 23647
rect 23581 23613 23615 23647
rect 23765 23613 23799 23647
rect 24041 23613 24075 23647
rect 25513 23613 25547 23647
rect 6193 23545 6227 23579
rect 7665 23545 7699 23579
rect 13185 23545 13219 23579
rect 16865 23545 16899 23579
rect 10425 23477 10459 23511
rect 15025 23477 15059 23511
rect 16037 23477 16071 23511
rect 17785 23477 17819 23511
rect 17969 23477 18003 23511
rect 18337 23477 18371 23511
rect 18521 23477 18555 23511
rect 21833 23477 21867 23511
rect 27721 23477 27755 23511
rect 8585 23273 8619 23307
rect 9965 23273 9999 23307
rect 12265 23273 12299 23307
rect 12817 23273 12851 23307
rect 19257 23273 19291 23307
rect 22201 23273 22235 23307
rect 22385 23273 22419 23307
rect 22753 23273 22787 23307
rect 24133 23273 24167 23307
rect 26801 23273 26835 23307
rect 26985 23273 27019 23307
rect 9689 23205 9723 23239
rect 11437 23205 11471 23239
rect 16957 23205 16991 23239
rect 22661 23205 22695 23239
rect 22845 23205 22879 23239
rect 27261 23205 27295 23239
rect 4997 23137 5031 23171
rect 5457 23137 5491 23171
rect 12173 23137 12207 23171
rect 13001 23137 13035 23171
rect 14197 23137 14231 23171
rect 22477 23137 22511 23171
rect 24409 23137 24443 23171
rect 24777 23137 24811 23171
rect 24869 23137 24903 23171
rect 27077 23137 27111 23171
rect 1501 23069 1535 23103
rect 1685 23069 1719 23103
rect 2605 23069 2639 23103
rect 2789 23069 2823 23103
rect 2973 23069 3007 23103
rect 3065 23069 3099 23103
rect 3249 23069 3283 23103
rect 4905 23069 4939 23103
rect 5089 23069 5123 23103
rect 6837 23069 6871 23103
rect 7021 23069 7055 23103
rect 9597 23069 9631 23103
rect 10149 23069 10183 23103
rect 10241 23069 10275 23103
rect 10425 23069 10459 23103
rect 10517 23069 10551 23103
rect 10609 23069 10643 23103
rect 10701 23069 10735 23103
rect 10885 23069 10919 23103
rect 11161 23069 11195 23103
rect 11437 23069 11471 23103
rect 12449 23069 12483 23103
rect 12725 23069 12759 23103
rect 14289 23069 14323 23103
rect 16865 23069 16899 23103
rect 17049 23069 17083 23103
rect 19441 23069 19475 23103
rect 19717 23069 19751 23103
rect 21925 23069 21959 23103
rect 22753 23069 22787 23103
rect 23121 23069 23155 23103
rect 23949 23069 23983 23103
rect 24133 23069 24167 23103
rect 25421 23069 25455 23103
rect 25605 23069 25639 23103
rect 27353 23069 27387 23103
rect 27629 23069 27663 23103
rect 2881 23001 2915 23035
rect 6285 23001 6319 23035
rect 8401 23001 8435 23035
rect 11345 23001 11379 23035
rect 22017 23001 22051 23035
rect 22845 23001 22879 23035
rect 25053 23001 25087 23035
rect 26617 23001 26651 23035
rect 2329 22933 2363 22967
rect 3157 22933 3191 22967
rect 8601 22933 8635 22967
rect 8769 22933 8803 22967
rect 11069 22933 11103 22967
rect 12633 22933 12667 22967
rect 13001 22933 13035 22967
rect 14657 22933 14691 22967
rect 19625 22933 19659 22967
rect 21741 22933 21775 22967
rect 22227 22933 22261 22967
rect 23029 22933 23063 22967
rect 25421 22933 25455 22967
rect 26817 22933 26851 22967
rect 27353 22933 27387 22967
rect 27445 22933 27479 22967
rect 2513 22729 2547 22763
rect 3985 22729 4019 22763
rect 4077 22729 4111 22763
rect 6929 22729 6963 22763
rect 7941 22729 7975 22763
rect 9689 22729 9723 22763
rect 10057 22729 10091 22763
rect 18889 22729 18923 22763
rect 25329 22729 25363 22763
rect 26249 22729 26283 22763
rect 3801 22661 3835 22695
rect 7573 22661 7607 22695
rect 8125 22661 8159 22695
rect 8861 22661 8895 22695
rect 9229 22661 9263 22695
rect 18613 22661 18647 22695
rect 19349 22661 19383 22695
rect 20269 22661 20303 22695
rect 22201 22661 22235 22695
rect 22385 22661 22419 22695
rect 25237 22661 25271 22695
rect 25497 22661 25531 22695
rect 25697 22661 25731 22695
rect 1869 22593 1903 22627
rect 4169 22593 4203 22627
rect 6745 22593 6779 22627
rect 6929 22593 6963 22627
rect 7481 22593 7515 22627
rect 7665 22593 7699 22627
rect 7849 22593 7883 22627
rect 9045 22593 9079 22627
rect 9597 22593 9631 22627
rect 9873 22593 9907 22627
rect 12633 22593 12667 22627
rect 12817 22593 12851 22627
rect 18153 22593 18187 22627
rect 18337 22593 18371 22627
rect 18429 22593 18463 22627
rect 18703 22615 18737 22649
rect 18797 22599 18831 22633
rect 19073 22593 19107 22627
rect 20177 22593 20211 22627
rect 20361 22593 20395 22627
rect 26341 22593 26375 22627
rect 27169 22593 27203 22627
rect 27537 22593 27571 22627
rect 1961 22525 1995 22559
rect 2881 22525 2915 22559
rect 3617 22525 3651 22559
rect 12541 22525 12575 22559
rect 24777 22525 24811 22559
rect 26985 22525 27019 22559
rect 4353 22457 4387 22491
rect 8125 22457 8159 22491
rect 19073 22457 19107 22491
rect 19717 22457 19751 22491
rect 24961 22457 24995 22491
rect 27721 22457 27755 22491
rect 13001 22389 13035 22423
rect 18245 22389 18279 22423
rect 18521 22389 18555 22423
rect 19165 22389 19199 22423
rect 19349 22389 19383 22423
rect 25513 22389 25547 22423
rect 27353 22389 27387 22423
rect 12633 22185 12667 22219
rect 14657 22185 14691 22219
rect 17141 22185 17175 22219
rect 21189 22185 21223 22219
rect 24041 22185 24075 22219
rect 25513 22185 25547 22219
rect 25789 22185 25823 22219
rect 25881 22117 25915 22151
rect 26433 22117 26467 22151
rect 3065 22049 3099 22083
rect 9505 22049 9539 22083
rect 9873 22049 9907 22083
rect 10701 22049 10735 22083
rect 20729 22049 20763 22083
rect 21097 22049 21131 22083
rect 1409 21981 1443 22015
rect 2697 21981 2731 22015
rect 2881 21981 2915 22015
rect 3985 21981 4019 22015
rect 4179 21981 4213 22015
rect 4353 21981 4387 22015
rect 4813 21981 4847 22015
rect 5273 21981 5307 22015
rect 9413 21981 9447 22015
rect 9597 21981 9631 22015
rect 10149 21981 10183 22015
rect 11621 21981 11655 22015
rect 11805 21981 11839 22015
rect 11897 21981 11931 22015
rect 12173 21981 12207 22015
rect 12449 21981 12483 22015
rect 12725 21981 12759 22015
rect 14933 21981 14967 22015
rect 15117 21981 15151 22015
rect 20913 21981 20947 22015
rect 21189 21981 21223 22015
rect 21373 21981 21407 22015
rect 24593 21981 24627 22015
rect 24685 21981 24719 22015
rect 24869 21981 24903 22015
rect 25789 21981 25823 22015
rect 26065 21981 26099 22015
rect 26157 21981 26191 22015
rect 26433 21981 26467 22015
rect 27537 21981 27571 22015
rect 1961 21913 1995 21947
rect 12357 21913 12391 21947
rect 14473 21913 14507 21947
rect 14673 21913 14707 21947
rect 17120 21913 17154 21947
rect 17325 21913 17359 21947
rect 23857 21913 23891 21947
rect 25329 21913 25363 21947
rect 1593 21845 1627 21879
rect 3985 21845 4019 21879
rect 4445 21845 4479 21879
rect 11713 21845 11747 21879
rect 11989 21845 12023 21879
rect 13001 21845 13035 21879
rect 14841 21845 14875 21879
rect 15025 21845 15059 21879
rect 16957 21845 16991 21879
rect 24067 21845 24101 21879
rect 24225 21845 24259 21879
rect 25053 21845 25087 21879
rect 25529 21845 25563 21879
rect 25697 21845 25731 21879
rect 26249 21845 26283 21879
rect 27721 21845 27755 21879
rect 14289 21641 14323 21675
rect 14473 21641 14507 21675
rect 16313 21641 16347 21675
rect 24961 21641 24995 21675
rect 26801 21641 26835 21675
rect 2513 21573 2547 21607
rect 2881 21573 2915 21607
rect 14381 21573 14415 21607
rect 16497 21573 16531 21607
rect 17693 21573 17727 21607
rect 25329 21573 25363 21607
rect 27077 21573 27111 21607
rect 1409 21505 1443 21539
rect 2237 21505 2271 21539
rect 3617 21505 3651 21539
rect 3985 21505 4019 21539
rect 4905 21505 4939 21539
rect 5089 21505 5123 21539
rect 7573 21505 7607 21539
rect 7757 21505 7791 21539
rect 15025 21505 15059 21539
rect 15301 21505 15335 21539
rect 15393 21505 15427 21539
rect 15577 21505 15611 21539
rect 16221 21505 16255 21539
rect 16957 21505 16991 21539
rect 17785 21505 17819 21539
rect 18245 21505 18279 21539
rect 18613 21505 18647 21539
rect 18981 21505 19015 21539
rect 19533 21505 19567 21539
rect 24317 21505 24351 21539
rect 24501 21505 24535 21539
rect 24777 21505 24811 21539
rect 27813 21505 27847 21539
rect 4629 21437 4663 21471
rect 4997 21437 5031 21471
rect 5365 21437 5399 21471
rect 5733 21437 5767 21471
rect 5825 21437 5859 21471
rect 14013 21437 14047 21471
rect 14749 21437 14783 21471
rect 16773 21437 16807 21471
rect 16865 21437 16899 21471
rect 17141 21437 17175 21471
rect 19441 21437 19475 21471
rect 25053 21437 25087 21471
rect 27261 21437 27295 21471
rect 8585 21369 8619 21403
rect 14105 21369 14139 21403
rect 15669 21369 15703 21403
rect 17325 21369 17359 21403
rect 19901 21369 19935 21403
rect 6009 21301 6043 21335
rect 13921 21301 13955 21335
rect 14933 21301 14967 21335
rect 15117 21301 15151 21335
rect 16497 21301 16531 21335
rect 27629 21301 27663 21335
rect 12265 21097 12299 21131
rect 14565 21097 14599 21131
rect 17233 21097 17267 21131
rect 14105 21029 14139 21063
rect 16497 21029 16531 21063
rect 17325 21029 17359 21063
rect 19901 21029 19935 21063
rect 20453 21029 20487 21063
rect 2513 20961 2547 20995
rect 11529 20961 11563 20995
rect 12081 20961 12115 20995
rect 14473 20961 14507 20995
rect 14841 20961 14875 20995
rect 15025 20961 15059 20995
rect 15117 20961 15151 20995
rect 16957 20961 16991 20995
rect 17049 20961 17083 20995
rect 17509 20961 17543 20995
rect 17601 20961 17635 20995
rect 17877 20961 17911 20995
rect 19625 20961 19659 20995
rect 22569 20961 22603 20995
rect 24961 20961 24995 20995
rect 4997 20893 5031 20927
rect 5273 20893 5307 20927
rect 5365 20893 5399 20927
rect 5549 20893 5583 20927
rect 6101 20893 6135 20927
rect 7573 20893 7607 20927
rect 11161 20893 11195 20927
rect 11253 20893 11287 20927
rect 11621 20893 11655 20927
rect 12357 20893 12391 20927
rect 13461 20893 13495 20927
rect 13645 20893 13679 20927
rect 14289 20893 14323 20927
rect 14565 20893 14599 20927
rect 14933 20893 14967 20927
rect 15669 20893 15703 20927
rect 15853 20893 15887 20927
rect 16037 20893 16071 20927
rect 16313 20893 16347 20927
rect 17969 20893 18003 20927
rect 18245 20893 18279 20927
rect 18521 20893 18555 20927
rect 18797 20893 18831 20927
rect 19073 20893 19107 20927
rect 19533 20893 19567 20927
rect 19809 20893 19843 20927
rect 19993 20893 20027 20927
rect 20085 20893 20119 20927
rect 20269 20893 20303 20927
rect 21649 20893 21683 20927
rect 21741 20893 21775 20927
rect 21925 20893 21959 20927
rect 22109 20893 22143 20927
rect 22201 20893 22235 20927
rect 22385 20893 22419 20927
rect 22661 20893 22695 20927
rect 24685 20893 24719 20927
rect 1961 20825 1995 20859
rect 8309 20825 8343 20859
rect 11897 20825 11931 20859
rect 16497 20825 16531 20859
rect 18613 20825 18647 20859
rect 18981 20825 19015 20859
rect 13553 20757 13587 20791
rect 14657 20757 14691 20791
rect 15393 20757 15427 20791
rect 16221 20757 16255 20791
rect 17785 20757 17819 20791
rect 18061 20757 18095 20791
rect 18429 20757 18463 20791
rect 19349 20757 19383 20791
rect 22293 20757 22327 20791
rect 26433 20757 26467 20791
rect 10793 20553 10827 20587
rect 13093 20553 13127 20587
rect 14841 20553 14875 20587
rect 15669 20553 15703 20587
rect 18797 20553 18831 20587
rect 20913 20553 20947 20587
rect 23581 20553 23615 20587
rect 11529 20485 11563 20519
rect 13461 20485 13495 20519
rect 17325 20485 17359 20519
rect 17509 20485 17543 20519
rect 20545 20485 20579 20519
rect 20761 20485 20795 20519
rect 22109 20485 22143 20519
rect 25513 20485 25547 20519
rect 25697 20485 25731 20519
rect 2053 20417 2087 20451
rect 2237 20417 2271 20451
rect 3525 20417 3559 20451
rect 3709 20417 3743 20451
rect 6745 20417 6779 20451
rect 6929 20417 6963 20451
rect 7941 20417 7975 20451
rect 8217 20417 8251 20451
rect 10977 20417 11011 20451
rect 11069 20417 11103 20451
rect 11253 20417 11287 20451
rect 11345 20417 11379 20451
rect 11621 20417 11655 20451
rect 11897 20417 11931 20451
rect 12081 20417 12115 20451
rect 12357 20417 12391 20451
rect 12449 20417 12483 20451
rect 13277 20417 13311 20451
rect 13737 20417 13771 20451
rect 13921 20417 13955 20451
rect 14013 20417 14047 20451
rect 14289 20417 14323 20451
rect 14473 20417 14507 20451
rect 15025 20417 15059 20451
rect 15117 20417 15151 20451
rect 15301 20417 15335 20451
rect 15393 20417 15427 20451
rect 15485 20417 15519 20451
rect 16681 20417 16715 20451
rect 16957 20417 16991 20451
rect 17969 20417 18003 20451
rect 18061 20417 18095 20451
rect 18981 20417 19015 20451
rect 19073 20417 19107 20451
rect 19257 20417 19291 20451
rect 19349 20417 19383 20451
rect 19533 20417 19567 20451
rect 21189 20417 21223 20451
rect 21281 20417 21315 20451
rect 21373 20417 21407 20451
rect 21557 20417 21591 20451
rect 21649 20417 21683 20451
rect 2145 20349 2179 20383
rect 2605 20349 2639 20383
rect 3433 20349 3467 20383
rect 6837 20349 6871 20383
rect 7205 20349 7239 20383
rect 14657 20349 14691 20383
rect 17785 20349 17819 20383
rect 21833 20349 21867 20383
rect 7665 20281 7699 20315
rect 17233 20281 17267 20315
rect 18061 20281 18095 20315
rect 3525 20213 3559 20247
rect 13553 20213 13587 20247
rect 13921 20213 13955 20247
rect 16773 20213 16807 20247
rect 17693 20213 17727 20247
rect 19625 20213 19659 20247
rect 20729 20213 20763 20247
rect 21005 20213 21039 20247
rect 12173 20009 12207 20043
rect 13461 20009 13495 20043
rect 19533 20009 19567 20043
rect 22201 20009 22235 20043
rect 22661 20009 22695 20043
rect 27813 20009 27847 20043
rect 12725 19941 12759 19975
rect 14105 19941 14139 19975
rect 2053 19873 2087 19907
rect 2697 19873 2731 19907
rect 3157 19873 3191 19907
rect 3341 19873 3375 19907
rect 3433 19873 3467 19907
rect 3617 19873 3651 19907
rect 7757 19873 7791 19907
rect 10333 19873 10367 19907
rect 12081 19873 12115 19907
rect 14381 19873 14415 19907
rect 21005 19873 21039 19907
rect 21557 19873 21591 19907
rect 22569 19873 22603 19907
rect 26065 19873 26099 19907
rect 1409 19805 1443 19839
rect 2145 19805 2179 19839
rect 3249 19805 3283 19839
rect 4445 19805 4479 19839
rect 4721 19805 4755 19839
rect 5365 19805 5399 19839
rect 5549 19805 5583 19839
rect 7665 19805 7699 19839
rect 12357 19805 12391 19839
rect 12633 19805 12667 19839
rect 12817 19805 12851 19839
rect 13645 19805 13679 19839
rect 13829 19805 13863 19839
rect 14473 19805 14507 19839
rect 19717 19805 19751 19839
rect 19901 19805 19935 19839
rect 21189 19805 21223 19839
rect 21281 19805 21315 19839
rect 21741 19805 21775 19839
rect 21833 19805 21867 19839
rect 22017 19805 22051 19839
rect 22109 19805 22143 19839
rect 22385 19805 22419 19839
rect 10609 19737 10643 19771
rect 12541 19737 12575 19771
rect 22661 19737 22695 19771
rect 26341 19737 26375 19771
rect 1593 19669 1627 19703
rect 5273 19669 5307 19703
rect 5549 19669 5583 19703
rect 8033 19669 8067 19703
rect 21005 19669 21039 19703
rect 8033 19465 8067 19499
rect 20729 19465 20763 19499
rect 21833 19465 21867 19499
rect 2881 19397 2915 19431
rect 4537 19397 4571 19431
rect 18429 19397 18463 19431
rect 18613 19397 18647 19431
rect 19165 19397 19199 19431
rect 21985 19397 22019 19431
rect 22201 19397 22235 19431
rect 22293 19397 22327 19431
rect 2789 19329 2823 19363
rect 2973 19329 3007 19363
rect 3341 19329 3375 19363
rect 4445 19329 4479 19363
rect 4997 19329 5031 19363
rect 5089 19329 5123 19363
rect 5457 19329 5491 19363
rect 6009 19329 6043 19363
rect 6377 19329 6411 19363
rect 6561 19329 6595 19363
rect 7941 19329 7975 19363
rect 8217 19329 8251 19363
rect 8585 19329 8619 19363
rect 8769 19329 8803 19363
rect 12817 19329 12851 19363
rect 18705 19329 18739 19363
rect 18981 19329 19015 19363
rect 19441 19329 19475 19363
rect 19809 19329 19843 19363
rect 20269 19329 20303 19363
rect 20545 19329 20579 19363
rect 20637 19329 20671 19363
rect 20821 19329 20855 19363
rect 22477 19329 22511 19363
rect 22569 19329 22603 19363
rect 3433 19261 3467 19295
rect 4077 19261 4111 19295
rect 12725 19261 12759 19295
rect 12909 19261 12943 19295
rect 13001 19261 13035 19295
rect 19533 19261 19567 19295
rect 19717 19261 19751 19295
rect 9781 19193 9815 19227
rect 18797 19193 18831 19227
rect 19809 19193 19843 19227
rect 20453 19193 20487 19227
rect 22293 19193 22327 19227
rect 6193 19125 6227 19159
rect 6469 19125 6503 19159
rect 8217 19125 8251 19159
rect 12541 19125 12575 19159
rect 18429 19125 18463 19159
rect 22017 19125 22051 19159
rect 8217 18921 8251 18955
rect 13001 18921 13035 18955
rect 14105 18921 14139 18955
rect 24225 18921 24259 18955
rect 8677 18785 8711 18819
rect 9045 18785 9079 18819
rect 12449 18785 12483 18819
rect 13829 18785 13863 18819
rect 21833 18785 21867 18819
rect 22477 18785 22511 18819
rect 4905 18717 4939 18751
rect 5365 18717 5399 18751
rect 6101 18717 6135 18751
rect 6561 18717 6595 18751
rect 8401 18717 8435 18751
rect 8493 18717 8527 18751
rect 8769 18717 8803 18751
rect 9137 18717 9171 18751
rect 9597 18717 9631 18751
rect 9781 18717 9815 18751
rect 12357 18717 12391 18751
rect 12817 18717 12851 18751
rect 12909 18717 12943 18751
rect 13737 18717 13771 18751
rect 14381 18717 14415 18751
rect 14473 18717 14507 18751
rect 14565 18717 14599 18751
rect 14749 18717 14783 18751
rect 17969 18717 18003 18751
rect 18153 18717 18187 18751
rect 18429 18717 18463 18751
rect 18613 18717 18647 18751
rect 18705 18717 18739 18751
rect 18061 18649 18095 18683
rect 18291 18649 18325 18683
rect 20085 18649 20119 18683
rect 22753 18649 22787 18683
rect 5733 18581 5767 18615
rect 9505 18581 9539 18615
rect 9689 18581 9723 18615
rect 12725 18581 12759 18615
rect 13185 18581 13219 18615
rect 17785 18581 17819 18615
rect 18889 18581 18923 18615
rect 4997 18377 5031 18411
rect 7297 18377 7331 18411
rect 12449 18377 12483 18411
rect 12541 18377 12575 18411
rect 15945 18377 15979 18411
rect 18429 18377 18463 18411
rect 20729 18377 20763 18411
rect 21925 18377 21959 18411
rect 1961 18309 1995 18343
rect 2329 18309 2363 18343
rect 6745 18309 6779 18343
rect 10241 18309 10275 18343
rect 17141 18309 17175 18343
rect 22661 18309 22695 18343
rect 1501 18241 1535 18275
rect 3249 18241 3283 18275
rect 4905 18241 4939 18275
rect 5089 18241 5123 18275
rect 6377 18241 6411 18275
rect 7297 18241 7331 18275
rect 9229 18241 9263 18275
rect 9413 18241 9447 18275
rect 9505 18241 9539 18275
rect 9873 18241 9907 18275
rect 10149 18241 10183 18275
rect 12173 18241 12207 18275
rect 12633 18241 12667 18275
rect 12725 18241 12759 18275
rect 14013 18241 14047 18275
rect 14657 18241 14691 18275
rect 15025 18241 15059 18275
rect 15209 18241 15243 18275
rect 16129 18241 16163 18275
rect 16773 18241 16807 18275
rect 18981 18241 19015 18275
rect 21833 18241 21867 18275
rect 22109 18241 22143 18275
rect 2973 18173 3007 18207
rect 3065 18173 3099 18207
rect 3157 18173 3191 18207
rect 7389 18173 7423 18207
rect 10057 18173 10091 18207
rect 12265 18173 12299 18207
rect 12817 18173 12851 18207
rect 14841 18173 14875 18207
rect 14933 18173 14967 18207
rect 16313 18173 16347 18207
rect 19257 18173 19291 18207
rect 9597 18105 9631 18139
rect 1593 18037 1627 18071
rect 3433 18037 3467 18071
rect 6469 18037 6503 18071
rect 9413 18037 9447 18071
rect 11989 18037 12023 18071
rect 14105 18037 14139 18071
rect 14473 18037 14507 18071
rect 22293 18037 22327 18071
rect 22937 18037 22971 18071
rect 3249 17833 3283 17867
rect 9321 17833 9355 17867
rect 12173 17833 12207 17867
rect 12265 17833 12299 17867
rect 14749 17765 14783 17799
rect 15117 17765 15151 17799
rect 15761 17765 15795 17799
rect 16313 17765 16347 17799
rect 16957 17765 16991 17799
rect 17877 17765 17911 17799
rect 1685 17697 1719 17731
rect 1961 17697 1995 17731
rect 2329 17697 2363 17731
rect 8309 17697 8343 17731
rect 10057 17697 10091 17731
rect 12265 17697 12299 17731
rect 14657 17697 14691 17731
rect 17509 17697 17543 17731
rect 21649 17697 21683 17731
rect 22385 17697 22419 17731
rect 22477 17697 22511 17731
rect 1593 17629 1627 17663
rect 3249 17629 3283 17663
rect 3433 17629 3467 17663
rect 7573 17629 7607 17663
rect 7665 17629 7699 17663
rect 9229 17629 9263 17663
rect 9413 17629 9447 17663
rect 9873 17629 9907 17663
rect 14565 17629 14599 17663
rect 14841 17629 14875 17663
rect 15117 17629 15151 17663
rect 15301 17629 15335 17663
rect 15761 17629 15795 17663
rect 16037 17629 16071 17663
rect 16313 17629 16347 17663
rect 16497 17629 16531 17663
rect 16589 17629 16623 17663
rect 16773 17629 16807 17663
rect 16865 17629 16899 17663
rect 17233 17629 17267 17663
rect 17693 17629 17727 17663
rect 18061 17629 18095 17663
rect 18337 17629 18371 17663
rect 18613 17629 18647 17663
rect 18889 17629 18923 17663
rect 20729 17629 20763 17663
rect 20913 17629 20947 17663
rect 21005 17629 21039 17663
rect 21097 17629 21131 17663
rect 21281 17629 21315 17663
rect 21465 17629 21499 17663
rect 21557 17629 21591 17663
rect 21833 17629 21867 17663
rect 22017 17629 22051 17663
rect 2881 17561 2915 17595
rect 11897 17561 11931 17595
rect 22753 17561 22787 17595
rect 10609 17493 10643 17527
rect 11989 17493 12023 17527
rect 15025 17493 15059 17527
rect 15945 17493 15979 17527
rect 18705 17493 18739 17527
rect 19073 17493 19107 17527
rect 24225 17493 24259 17527
rect 2421 17289 2455 17323
rect 7757 17289 7791 17323
rect 9321 17289 9355 17323
rect 19441 17289 19475 17323
rect 22385 17289 22419 17323
rect 11345 17221 11379 17255
rect 15853 17221 15887 17255
rect 22753 17221 22787 17255
rect 23581 17221 23615 17255
rect 1869 17153 1903 17187
rect 2329 17153 2363 17187
rect 2513 17153 2547 17187
rect 3525 17153 3559 17187
rect 3893 17153 3927 17187
rect 4629 17153 4663 17187
rect 4813 17153 4847 17187
rect 7573 17153 7607 17187
rect 7849 17153 7883 17187
rect 9045 17153 9079 17187
rect 9689 17153 9723 17187
rect 9873 17153 9907 17187
rect 11713 17153 11747 17187
rect 13645 17153 13679 17187
rect 13829 17153 13863 17187
rect 14473 17153 14507 17187
rect 14565 17153 14599 17187
rect 15669 17153 15703 17187
rect 15761 17153 15795 17187
rect 15991 17153 16025 17187
rect 16129 17153 16163 17187
rect 16865 17153 16899 17187
rect 17049 17153 17083 17187
rect 19349 17153 19383 17187
rect 19533 17153 19567 17187
rect 20085 17153 20119 17187
rect 21281 17153 21315 17187
rect 21373 17153 21407 17187
rect 22569 17153 22603 17187
rect 23029 17153 23063 17187
rect 23213 17153 23247 17187
rect 23489 17153 23523 17187
rect 23673 17153 23707 17187
rect 25237 17153 25271 17187
rect 1961 17085 1995 17119
rect 4537 17085 4571 17119
rect 8861 17085 8895 17119
rect 8953 17085 8987 17119
rect 9137 17085 9171 17119
rect 11989 17085 12023 17119
rect 14289 17085 14323 17119
rect 16957 17085 16991 17119
rect 19809 17085 19843 17119
rect 19993 17085 20027 17119
rect 23397 17085 23431 17119
rect 24961 17085 24995 17119
rect 2237 17017 2271 17051
rect 7573 17017 7607 17051
rect 15485 17017 15519 17051
rect 19257 17017 19291 17051
rect 4721 16949 4755 16983
rect 13461 16949 13495 16983
rect 13645 16949 13679 16983
rect 14381 16949 14415 16983
rect 19717 16949 19751 16983
rect 20361 16949 20395 16983
rect 12909 16745 12943 16779
rect 15853 16745 15887 16779
rect 16037 16745 16071 16779
rect 22017 16745 22051 16779
rect 23121 16745 23155 16779
rect 8953 16677 8987 16711
rect 20453 16677 20487 16711
rect 24869 16677 24903 16711
rect 2973 16609 3007 16643
rect 3525 16609 3559 16643
rect 8125 16609 8159 16643
rect 9321 16609 9355 16643
rect 12357 16609 12391 16643
rect 12817 16609 12851 16643
rect 14105 16609 14139 16643
rect 20545 16609 20579 16643
rect 20909 16609 20943 16643
rect 21097 16609 21131 16643
rect 21741 16609 21775 16643
rect 23029 16609 23063 16643
rect 2881 16541 2915 16575
rect 4721 16541 4755 16575
rect 5365 16541 5399 16575
rect 7389 16541 7423 16575
rect 7573 16541 7607 16575
rect 9413 16541 9447 16575
rect 9873 16541 9907 16575
rect 10241 16541 10275 16575
rect 10609 16541 10643 16575
rect 12081 16541 12115 16575
rect 12265 16541 12299 16575
rect 12449 16541 12483 16575
rect 12633 16541 12667 16575
rect 13093 16541 13127 16575
rect 13185 16541 13219 16575
rect 16129 16541 16163 16575
rect 19901 16541 19935 16575
rect 20315 16541 20349 16575
rect 20729 16541 20763 16575
rect 20821 16541 20855 16575
rect 21189 16541 21223 16575
rect 21649 16541 21683 16575
rect 21925 16541 21959 16575
rect 22109 16541 22143 16575
rect 22385 16541 22419 16575
rect 22477 16541 22511 16575
rect 22569 16541 22603 16575
rect 22753 16541 22787 16575
rect 22845 16541 22879 16575
rect 23305 16541 23339 16575
rect 23489 16541 23523 16575
rect 23581 16541 23615 16575
rect 23857 16541 23891 16575
rect 24133 16541 24167 16575
rect 12909 16473 12943 16507
rect 14381 16473 14415 16507
rect 20085 16473 20119 16507
rect 20177 16473 20211 16507
rect 23673 16473 23707 16507
rect 24685 16473 24719 16507
rect 13369 16405 13403 16439
rect 20545 16405 20579 16439
rect 20913 16405 20947 16439
rect 21281 16405 21315 16439
rect 22293 16405 22327 16439
rect 24041 16405 24075 16439
rect 2973 16201 3007 16235
rect 7481 16201 7515 16235
rect 10333 16201 10367 16235
rect 11989 16201 12023 16235
rect 14473 16201 14507 16235
rect 14749 16201 14783 16235
rect 17141 16201 17175 16235
rect 19625 16201 19659 16235
rect 23213 16201 23247 16235
rect 12633 16133 12667 16167
rect 23673 16133 23707 16167
rect 1409 16065 1443 16099
rect 2881 16065 2915 16099
rect 3065 16065 3099 16099
rect 3157 16065 3191 16099
rect 3617 16065 3651 16099
rect 3801 16065 3835 16099
rect 3893 16065 3927 16099
rect 4261 16065 4295 16099
rect 4629 16065 4663 16099
rect 5181 16065 5215 16099
rect 5641 16065 5675 16099
rect 5825 16065 5859 16099
rect 6929 16065 6963 16099
rect 7205 16065 7239 16099
rect 7297 16065 7331 16099
rect 7665 16065 7699 16099
rect 8309 16065 8343 16099
rect 9597 16065 9631 16099
rect 9965 16065 9999 16099
rect 10241 16065 10275 16099
rect 10425 16065 10459 16099
rect 12173 16065 12207 16099
rect 12265 16065 12299 16099
rect 12541 16065 12575 16099
rect 14565 16065 14599 16099
rect 14657 16065 14691 16099
rect 14933 16065 14967 16099
rect 15393 16065 15427 16099
rect 16681 16065 16715 16099
rect 16957 16065 16991 16099
rect 17417 16065 17451 16099
rect 17877 16065 17911 16099
rect 18061 16065 18095 16099
rect 18153 16065 18187 16099
rect 18889 16065 18923 16099
rect 19533 16065 19567 16099
rect 19809 16065 19843 16099
rect 23305 16065 23339 16099
rect 23397 16065 23431 16099
rect 1685 15997 1719 16031
rect 3249 15997 3283 16031
rect 4813 15997 4847 16031
rect 10057 15997 10091 16031
rect 14197 15997 14231 16031
rect 16865 15997 16899 16031
rect 18797 15997 18831 16031
rect 25145 15997 25179 16031
rect 15025 15929 15059 15963
rect 17693 15929 17727 15963
rect 3801 15861 3835 15895
rect 5733 15861 5767 15895
rect 7021 15861 7055 15895
rect 9321 15861 9355 15895
rect 9689 15861 9723 15895
rect 13829 15861 13863 15895
rect 14105 15861 14139 15895
rect 14289 15861 14323 15895
rect 15117 15861 15151 15895
rect 16681 15861 16715 15895
rect 17325 15861 17359 15895
rect 19993 15861 20027 15895
rect 12173 15657 12207 15691
rect 16129 15657 16163 15691
rect 16589 15657 16623 15691
rect 23949 15657 23983 15691
rect 24593 15657 24627 15691
rect 23397 15589 23431 15623
rect 23489 15589 23523 15623
rect 24409 15589 24443 15623
rect 4445 15521 4479 15555
rect 16221 15521 16255 15555
rect 17049 15521 17083 15555
rect 19073 15521 19107 15555
rect 20269 15521 20303 15555
rect 4353 15453 4387 15487
rect 7297 15453 7331 15487
rect 8125 15453 8159 15487
rect 9321 15453 9355 15487
rect 9781 15453 9815 15487
rect 11621 15453 11655 15487
rect 11805 15453 11839 15487
rect 11989 15453 12023 15487
rect 16405 15453 16439 15487
rect 16773 15453 16807 15487
rect 16957 15453 16991 15487
rect 19993 15453 20027 15487
rect 20177 15453 20211 15487
rect 20913 15453 20947 15487
rect 21097 15453 21131 15487
rect 23213 15453 23247 15487
rect 23581 15453 23615 15487
rect 23673 15453 23707 15487
rect 8769 15385 8803 15419
rect 11897 15385 11931 15419
rect 16129 15385 16163 15419
rect 16865 15385 16899 15419
rect 17325 15385 17359 15419
rect 24777 15385 24811 15419
rect 4721 15317 4755 15351
rect 19809 15317 19843 15351
rect 21097 15317 21131 15351
rect 24567 15317 24601 15351
rect 8585 15113 8619 15147
rect 12357 15113 12391 15147
rect 14197 15113 14231 15147
rect 16865 15113 16899 15147
rect 17417 15113 17451 15147
rect 20821 15113 20855 15147
rect 23397 15113 23431 15147
rect 8217 15045 8251 15079
rect 8401 15045 8435 15079
rect 9045 15045 9079 15079
rect 20729 15045 20763 15079
rect 23765 15045 23799 15079
rect 2513 14977 2547 15011
rect 2697 14977 2731 15011
rect 3433 14977 3467 15011
rect 3525 14977 3559 15011
rect 4169 14977 4203 15011
rect 4353 14977 4387 15011
rect 5089 14977 5123 15011
rect 5273 14977 5307 15011
rect 6377 14977 6411 15011
rect 7297 14977 7331 15011
rect 7481 14977 7515 15011
rect 8677 14977 8711 15011
rect 8861 14977 8895 15011
rect 9873 14977 9907 15011
rect 10333 14977 10367 15011
rect 11805 14977 11839 15011
rect 11989 14977 12023 15011
rect 12081 14977 12115 15011
rect 12173 14977 12207 15011
rect 12633 14977 12667 15011
rect 12725 14977 12759 15011
rect 12909 14977 12943 15011
rect 13001 14977 13035 15011
rect 14289 14977 14323 15011
rect 14565 14977 14599 15011
rect 17049 14977 17083 15011
rect 17325 14977 17359 15011
rect 17601 14977 17635 15011
rect 17969 14977 18003 15011
rect 18153 14977 18187 15011
rect 19993 14977 20027 15011
rect 20269 14977 20303 15011
rect 21005 14977 21039 15011
rect 21281 14977 21315 15011
rect 21465 14977 21499 15011
rect 21649 14977 21683 15011
rect 23121 14977 23155 15011
rect 23949 14977 23983 15011
rect 24041 14977 24075 15011
rect 4077 14909 4111 14943
rect 6101 14909 6135 14943
rect 14197 14909 14231 14943
rect 14381 14909 14415 14943
rect 14657 14909 14691 14943
rect 17233 14909 17267 14943
rect 17785 14909 17819 14943
rect 17877 14909 17911 14943
rect 20453 14909 20487 14943
rect 6745 14841 6779 14875
rect 21097 14841 21131 14875
rect 21189 14841 21223 14875
rect 23765 14841 23799 14875
rect 2697 14773 2731 14807
rect 4261 14773 4295 14807
rect 12449 14773 12483 14807
rect 17325 14773 17359 14807
rect 18705 14773 18739 14807
rect 20085 14773 20119 14807
rect 20637 14773 20671 14807
rect 21465 14773 21499 14807
rect 3341 14569 3375 14603
rect 15117 14569 15151 14603
rect 17601 14569 17635 14603
rect 18429 14569 18463 14603
rect 18613 14569 18647 14603
rect 22109 14569 22143 14603
rect 2605 14501 2639 14535
rect 4077 14501 4111 14535
rect 5549 14501 5583 14535
rect 6377 14501 6411 14535
rect 17371 14501 17405 14535
rect 19441 14501 19475 14535
rect 20637 14501 20671 14535
rect 23397 14501 23431 14535
rect 2329 14433 2363 14467
rect 2881 14433 2915 14467
rect 3157 14433 3191 14467
rect 4353 14433 4387 14467
rect 5273 14433 5307 14467
rect 5733 14433 5767 14467
rect 6929 14433 6963 14467
rect 11069 14433 11103 14467
rect 14887 14433 14921 14467
rect 15025 14433 15059 14467
rect 16957 14433 16991 14467
rect 17141 14433 17175 14467
rect 18245 14433 18279 14467
rect 19625 14433 19659 14467
rect 20913 14433 20947 14467
rect 23857 14433 23891 14467
rect 2237 14365 2271 14399
rect 2973 14365 3007 14399
rect 3065 14365 3099 14399
rect 3893 14365 3927 14399
rect 3985 14365 4019 14399
rect 4169 14365 4203 14399
rect 6101 14365 6135 14399
rect 6745 14365 6779 14399
rect 13185 14365 13219 14399
rect 13461 14365 13495 14399
rect 14749 14365 14783 14399
rect 15209 14365 15243 14399
rect 16865 14365 16899 14399
rect 17233 14365 17267 14399
rect 17509 14365 17543 14399
rect 17693 14365 17727 14399
rect 18429 14365 18463 14399
rect 19441 14365 19475 14399
rect 19809 14365 19843 14399
rect 21005 14365 21039 14399
rect 22477 14365 22511 14399
rect 22569 14365 22603 14399
rect 22753 14365 22787 14399
rect 22845 14365 22879 14399
rect 23489 14365 23523 14399
rect 23765 14365 23799 14399
rect 23949 14365 23983 14399
rect 24041 14365 24075 14399
rect 11345 14297 11379 14331
rect 18153 14297 18187 14331
rect 22017 14297 22051 14331
rect 24501 14297 24535 14331
rect 12817 14229 12851 14263
rect 13001 14229 13035 14263
rect 13369 14229 13403 14263
rect 17141 14229 17175 14263
rect 23029 14229 23063 14263
rect 23581 14229 23615 14263
rect 24593 14229 24627 14263
rect 11621 14025 11655 14059
rect 11897 14025 11931 14059
rect 15853 14025 15887 14059
rect 22385 14025 22419 14059
rect 22569 14025 22603 14059
rect 25329 14025 25363 14059
rect 27629 14025 27663 14059
rect 3249 13957 3283 13991
rect 3893 13957 3927 13991
rect 15485 13957 15519 13991
rect 15577 13957 15611 13991
rect 18613 13957 18647 13991
rect 23857 13957 23891 13991
rect 25513 13957 25547 13991
rect 1409 13889 1443 13923
rect 2697 13889 2731 13923
rect 3157 13889 3191 13923
rect 3341 13889 3375 13923
rect 3807 13889 3841 13923
rect 3985 13889 4019 13923
rect 4169 13889 4203 13923
rect 4353 13889 4387 13923
rect 6561 13889 6595 13923
rect 10609 13889 10643 13923
rect 11713 13889 11747 13923
rect 12173 13889 12207 13923
rect 12357 13889 12391 13923
rect 12541 13889 12575 13923
rect 14381 13889 14415 13923
rect 14565 13889 14599 13923
rect 14933 13889 14967 13923
rect 15301 13889 15335 13923
rect 15669 13889 15703 13923
rect 18061 13889 18095 13923
rect 18337 13889 18371 13923
rect 18429 13889 18463 13923
rect 22017 13889 22051 13923
rect 22109 13889 22143 13923
rect 22937 13889 22971 13923
rect 23305 13889 23339 13923
rect 23397 13889 23431 13923
rect 27813 13889 27847 13923
rect 2145 13821 2179 13855
rect 2789 13821 2823 13855
rect 5181 13821 5215 13855
rect 6653 13821 6687 13855
rect 8493 13821 8527 13855
rect 10701 13821 10735 13855
rect 12081 13821 12115 13855
rect 12265 13821 12299 13855
rect 14657 13821 14691 13855
rect 14749 13821 14783 13855
rect 18153 13821 18187 13855
rect 21925 13821 21959 13855
rect 22201 13821 22235 13855
rect 22477 13821 22511 13855
rect 23029 13821 23063 13855
rect 23581 13821 23615 13855
rect 25789 13821 25823 13855
rect 3065 13753 3099 13787
rect 8769 13753 8803 13787
rect 15117 13753 15151 13787
rect 6837 13685 6871 13719
rect 8953 13685 8987 13719
rect 12633 13685 12667 13719
rect 14381 13685 14415 13719
rect 2421 13481 2455 13515
rect 7389 13481 7423 13515
rect 8677 13481 8711 13515
rect 12173 13481 12207 13515
rect 12449 13481 12483 13515
rect 22937 13481 22971 13515
rect 23213 13481 23247 13515
rect 7849 13413 7883 13447
rect 15945 13413 15979 13447
rect 17417 13413 17451 13447
rect 24409 13413 24443 13447
rect 1961 13345 1995 13379
rect 2237 13345 2271 13379
rect 14105 13345 14139 13379
rect 17693 13345 17727 13379
rect 23489 13345 23523 13379
rect 24685 13345 24719 13379
rect 1869 13277 1903 13311
rect 2329 13277 2363 13311
rect 2513 13277 2547 13311
rect 6837 13277 6871 13311
rect 7113 13277 7147 13311
rect 7481 13277 7515 13311
rect 7573 13277 7607 13311
rect 8125 13277 8159 13311
rect 8217 13277 8251 13311
rect 8401 13277 8435 13311
rect 8493 13277 8527 13311
rect 9045 13277 9079 13311
rect 9229 13277 9263 13311
rect 12357 13277 12391 13311
rect 12449 13277 12483 13311
rect 13001 13277 13035 13311
rect 16129 13277 16163 13311
rect 16405 13277 16439 13311
rect 17509 13277 17543 13311
rect 17601 13277 17635 13311
rect 17877 13277 17911 13311
rect 20177 13277 20211 13311
rect 20545 13277 20579 13311
rect 21925 13277 21959 13311
rect 22109 13277 22143 13311
rect 22477 13277 22511 13311
rect 22845 13277 22879 13311
rect 22937 13277 22971 13311
rect 23581 13277 23615 13311
rect 24777 13277 24811 13311
rect 7665 13209 7699 13243
rect 7849 13209 7883 13243
rect 10057 13209 10091 13243
rect 12633 13209 12667 13243
rect 14381 13209 14415 13243
rect 17325 13209 17359 13243
rect 12817 13141 12851 13175
rect 15853 13141 15887 13175
rect 16313 13141 16347 13175
rect 20085 13141 20119 13175
rect 20453 13141 20487 13175
rect 22293 13141 22327 13175
rect 23121 13141 23155 13175
rect 6653 12937 6687 12971
rect 8125 12937 8159 12971
rect 8493 12937 8527 12971
rect 12265 12937 12299 12971
rect 12449 12937 12483 12971
rect 14933 12937 14967 12971
rect 21281 12937 21315 12971
rect 23397 12937 23431 12971
rect 11897 12869 11931 12903
rect 12097 12869 12131 12903
rect 15853 12869 15887 12903
rect 19257 12869 19291 12903
rect 22201 12869 22235 12903
rect 1961 12801 1995 12835
rect 6193 12801 6227 12835
rect 6469 12801 6503 12835
rect 6653 12801 6687 12835
rect 8033 12801 8067 12835
rect 8309 12801 8343 12835
rect 8861 12801 8895 12835
rect 12357 12801 12391 12835
rect 12541 12801 12575 12835
rect 15117 12801 15151 12835
rect 15301 12801 15335 12835
rect 15485 12801 15519 12835
rect 15669 12801 15703 12835
rect 15761 12801 15795 12835
rect 18061 12801 18095 12835
rect 18429 12801 18463 12835
rect 21833 12801 21867 12835
rect 22017 12801 22051 12835
rect 23397 12801 23431 12835
rect 23765 12801 23799 12835
rect 2053 12733 2087 12767
rect 5365 12733 5399 12767
rect 8769 12733 8803 12767
rect 9689 12733 9723 12767
rect 15393 12733 15427 12767
rect 17785 12733 17819 12767
rect 18337 12733 18371 12767
rect 19533 12733 19567 12767
rect 19809 12733 19843 12767
rect 23213 12733 23247 12767
rect 18889 12665 18923 12699
rect 2237 12597 2271 12631
rect 12081 12597 12115 12631
rect 17877 12597 17911 12631
rect 17969 12597 18003 12631
rect 19257 12597 19291 12631
rect 19441 12597 19475 12631
rect 19533 12393 19567 12427
rect 21649 12393 21683 12427
rect 4629 12325 4663 12359
rect 5549 12325 5583 12359
rect 16589 12325 16623 12359
rect 21189 12325 21223 12359
rect 3157 12257 3191 12291
rect 8309 12257 8343 12291
rect 12265 12257 12299 12291
rect 12449 12257 12483 12291
rect 12725 12257 12759 12291
rect 16405 12257 16439 12291
rect 20545 12257 20579 12291
rect 21281 12257 21315 12291
rect 3249 12189 3283 12223
rect 3801 12189 3835 12223
rect 3985 12189 4019 12223
rect 4537 12189 4571 12223
rect 4721 12189 4755 12223
rect 4905 12189 4939 12223
rect 5457 12189 5491 12223
rect 5641 12189 5675 12223
rect 6193 12189 6227 12223
rect 6561 12189 6595 12223
rect 7389 12189 7423 12223
rect 11345 12189 11379 12223
rect 11621 12189 11655 12223
rect 11897 12189 11931 12223
rect 12173 12189 12207 12223
rect 12357 12189 12391 12223
rect 12633 12189 12667 12223
rect 12909 12189 12943 12223
rect 16129 12189 16163 12223
rect 16313 12189 16347 12223
rect 16589 12189 16623 12223
rect 16957 12189 16991 12223
rect 17233 12189 17267 12223
rect 18153 12189 18187 12223
rect 18613 12189 18647 12223
rect 18797 12189 18831 12223
rect 18889 12189 18923 12223
rect 19073 12189 19107 12223
rect 19257 12189 19291 12223
rect 19441 12189 19475 12223
rect 19717 12189 19751 12223
rect 19993 12189 20027 12223
rect 20269 12189 20303 12223
rect 20453 12189 20487 12223
rect 20637 12189 20671 12223
rect 20821 12189 20855 12223
rect 21005 12189 21039 12223
rect 21189 12189 21223 12223
rect 21465 12189 21499 12223
rect 3893 12121 3927 12155
rect 4261 12121 4295 12155
rect 7205 12121 7239 12155
rect 19349 12121 19383 12155
rect 19901 12121 19935 12155
rect 3617 12053 3651 12087
rect 11161 12053 11195 12087
rect 11529 12053 11563 12087
rect 13093 12053 13127 12087
rect 16497 12053 16531 12087
rect 16773 12053 16807 12087
rect 17141 12053 17175 12087
rect 18245 12053 18279 12087
rect 18705 12053 18739 12087
rect 18981 12053 19015 12087
rect 20085 12053 20119 12087
rect 3709 11849 3743 11883
rect 7665 11849 7699 11883
rect 11345 11849 11379 11883
rect 11529 11849 11563 11883
rect 16405 11849 16439 11883
rect 19349 11849 19383 11883
rect 21097 11849 21131 11883
rect 23029 11849 23063 11883
rect 10977 11781 11011 11815
rect 12541 11781 12575 11815
rect 23397 11781 23431 11815
rect 1409 11713 1443 11747
rect 2881 11713 2915 11747
rect 3065 11713 3099 11747
rect 4629 11713 4663 11747
rect 5089 11713 5123 11747
rect 5273 11713 5307 11747
rect 7573 11713 7607 11747
rect 7757 11713 7791 11747
rect 10885 11713 10919 11747
rect 11161 11713 11195 11747
rect 11713 11713 11747 11747
rect 11805 11713 11839 11747
rect 11989 11713 12023 11747
rect 12081 11713 12115 11747
rect 12173 11713 12207 11747
rect 12265 11713 12299 11747
rect 12357 11713 12391 11747
rect 12633 11713 12667 11747
rect 15485 11713 15519 11747
rect 15577 11713 15611 11747
rect 15761 11713 15795 11747
rect 15853 11713 15887 11747
rect 16129 11713 16163 11747
rect 16221 11713 16255 11747
rect 16497 11713 16531 11747
rect 16681 11713 16715 11747
rect 18705 11713 18739 11747
rect 18889 11713 18923 11747
rect 19073 11713 19107 11747
rect 19165 11713 19199 11747
rect 19533 11713 19567 11747
rect 19809 11713 19843 11747
rect 23213 11713 23247 11747
rect 23305 11713 23339 11747
rect 23581 11713 23615 11747
rect 23673 11713 23707 11747
rect 1685 11645 1719 11679
rect 2973 11645 3007 11679
rect 3249 11645 3283 11679
rect 3341 11645 3375 11679
rect 3433 11645 3467 11679
rect 3525 11645 3559 11679
rect 4537 11645 4571 11679
rect 5181 11645 5215 11679
rect 16313 11645 16347 11679
rect 18981 11645 19015 11679
rect 4997 11577 5031 11611
rect 16037 11577 16071 11611
rect 2697 11305 2731 11339
rect 10057 11305 10091 11339
rect 10241 11305 10275 11339
rect 11713 11305 11747 11339
rect 12541 11305 12575 11339
rect 13001 11305 13035 11339
rect 15117 11305 15151 11339
rect 18245 11305 18279 11339
rect 19441 11305 19475 11339
rect 19901 11305 19935 11339
rect 20177 11305 20211 11339
rect 23581 11305 23615 11339
rect 11621 11237 11655 11271
rect 15025 11237 15059 11271
rect 22845 11237 22879 11271
rect 23213 11237 23247 11271
rect 23305 11237 23339 11271
rect 2237 11169 2271 11203
rect 7205 11169 7239 11203
rect 10977 11169 11011 11203
rect 11069 11169 11103 11203
rect 11437 11169 11471 11203
rect 16129 11169 16163 11203
rect 19717 11169 19751 11203
rect 20361 11169 20395 11203
rect 24593 11169 24627 11203
rect 2329 11101 2363 11135
rect 7113 11101 7147 11135
rect 10517 11101 10551 11135
rect 10609 11101 10643 11135
rect 10793 11101 10827 11135
rect 10885 11101 10919 11135
rect 11345 11101 11379 11135
rect 11851 11101 11885 11135
rect 12265 11101 12299 11135
rect 12357 11101 12391 11135
rect 12449 11101 12483 11135
rect 12909 11101 12943 11135
rect 13093 11101 13127 11135
rect 14473 11101 14507 11135
rect 14657 11101 14691 11135
rect 14749 11101 14783 11135
rect 14841 11101 14875 11135
rect 15301 11101 15335 11135
rect 15669 11101 15703 11135
rect 15761 11101 15795 11135
rect 16037 11101 16071 11135
rect 18061 11101 18095 11135
rect 19993 11101 20027 11135
rect 20453 11101 20487 11135
rect 20913 11101 20947 11135
rect 21097 11101 21131 11135
rect 21189 11101 21223 11135
rect 22569 11101 22603 11135
rect 22937 11101 22971 11135
rect 23122 11101 23156 11135
rect 23397 11101 23431 11135
rect 6561 11033 6595 11067
rect 9873 11033 9907 11067
rect 10333 11033 10367 11067
rect 11989 11033 12023 11067
rect 12081 11033 12115 11067
rect 15393 11033 15427 11067
rect 15485 11033 15519 11067
rect 16405 11033 16439 11067
rect 22845 11033 22879 11067
rect 23857 11033 23891 11067
rect 24041 11033 24075 11067
rect 24869 11033 24903 11067
rect 7113 10965 7147 10999
rect 10073 10965 10107 10999
rect 12725 10965 12759 10999
rect 15945 10965 15979 10999
rect 17877 10965 17911 10999
rect 20729 10965 20763 10999
rect 22661 10965 22695 10999
rect 23673 10965 23707 10999
rect 2421 10761 2455 10795
rect 6745 10761 6779 10795
rect 8125 10761 8159 10795
rect 11253 10761 11287 10795
rect 12930 10761 12964 10795
rect 14289 10761 14323 10795
rect 15117 10761 15151 10795
rect 15669 10761 15703 10795
rect 18521 10761 18555 10795
rect 7757 10693 7791 10727
rect 7941 10693 7975 10727
rect 9137 10693 9171 10727
rect 12725 10693 12759 10727
rect 14565 10693 14599 10727
rect 14749 10693 14783 10727
rect 15209 10693 15243 10727
rect 16773 10693 16807 10727
rect 18429 10693 18463 10727
rect 20453 10693 20487 10727
rect 20637 10693 20671 10727
rect 21373 10693 21407 10727
rect 22845 10693 22879 10727
rect 23061 10693 23095 10727
rect 23581 10693 23615 10727
rect 1869 10625 1903 10659
rect 2329 10625 2363 10659
rect 2513 10625 2547 10659
rect 3065 10625 3099 10659
rect 3525 10625 3559 10659
rect 3709 10625 3743 10659
rect 5641 10625 5675 10659
rect 6377 10625 6411 10659
rect 6470 10625 6504 10659
rect 7021 10625 7055 10659
rect 7573 10625 7607 10659
rect 8401 10625 8435 10659
rect 8677 10625 8711 10659
rect 8861 10625 8895 10659
rect 8953 10625 8987 10659
rect 9321 10625 9355 10659
rect 11161 10625 11195 10659
rect 11345 10625 11379 10659
rect 11713 10625 11747 10659
rect 11897 10625 11931 10659
rect 12081 10625 12115 10659
rect 12265 10625 12299 10659
rect 14197 10625 14231 10659
rect 14473 10625 14507 10659
rect 14657 10625 14691 10659
rect 14933 10625 14967 10659
rect 15485 10625 15519 10659
rect 15761 10625 15795 10659
rect 15945 10625 15979 10659
rect 16129 10625 16163 10659
rect 16313 10625 16347 10659
rect 18981 10625 19015 10659
rect 19809 10625 19843 10659
rect 20085 10625 20119 10659
rect 20269 10625 20303 10659
rect 20545 10625 20579 10659
rect 20821 10625 20855 10659
rect 20913 10625 20947 10659
rect 21097 10625 21131 10659
rect 21189 10625 21223 10659
rect 21465 10625 21499 10659
rect 23305 10625 23339 10659
rect 25145 10625 25179 10659
rect 25329 10625 25363 10659
rect 1961 10557 1995 10591
rect 2973 10557 3007 10591
rect 3617 10557 3651 10591
rect 5549 10557 5583 10591
rect 6929 10557 6963 10591
rect 8033 10557 8067 10591
rect 8585 10557 8619 10591
rect 11989 10557 12023 10591
rect 15393 10557 15427 10591
rect 16037 10557 16071 10591
rect 18705 10557 18739 10591
rect 18797 10557 18831 10591
rect 18889 10557 18923 10591
rect 25237 10557 25271 10591
rect 3433 10489 3467 10523
rect 6009 10489 6043 10523
rect 7389 10489 7423 10523
rect 8769 10489 8803 10523
rect 13093 10489 13127 10523
rect 25053 10489 25087 10523
rect 2237 10421 2271 10455
rect 12449 10421 12483 10455
rect 12909 10421 12943 10455
rect 15485 10421 15519 10455
rect 16497 10421 16531 10455
rect 19901 10421 19935 10455
rect 23029 10421 23063 10455
rect 23213 10421 23247 10455
rect 7665 10217 7699 10251
rect 9137 10217 9171 10251
rect 9321 10217 9355 10251
rect 9965 10217 9999 10251
rect 10149 10217 10183 10251
rect 13921 10217 13955 10251
rect 14841 10217 14875 10251
rect 15292 10217 15326 10251
rect 16037 10217 16071 10251
rect 17141 10217 17175 10251
rect 18337 10217 18371 10251
rect 21925 10217 21959 10251
rect 23305 10217 23339 10251
rect 23765 10217 23799 10251
rect 8217 10149 8251 10183
rect 12725 10149 12759 10183
rect 15485 10149 15519 10183
rect 2145 10081 2179 10115
rect 18521 10081 18555 10115
rect 20177 10081 20211 10115
rect 20453 10081 20487 10115
rect 23397 10081 23431 10115
rect 24409 10081 24443 10115
rect 24685 10081 24719 10115
rect 2237 10013 2271 10047
rect 7573 10013 7607 10047
rect 7757 10013 7791 10047
rect 7849 10013 7883 10047
rect 8033 10013 8067 10047
rect 8493 10013 8527 10047
rect 8769 10013 8803 10047
rect 9781 10013 9815 10047
rect 10057 10013 10091 10047
rect 11161 10013 11195 10047
rect 12449 10013 12483 10047
rect 12909 10013 12943 10047
rect 13093 10013 13127 10047
rect 13277 10013 13311 10047
rect 13461 10013 13495 10047
rect 13737 10013 13771 10047
rect 14105 10013 14139 10047
rect 14289 10013 14323 10047
rect 14381 10013 14415 10047
rect 14473 10013 14507 10047
rect 14841 10013 14875 10047
rect 15025 10013 15059 10047
rect 16129 10013 16163 10047
rect 16497 10013 16531 10047
rect 16645 10013 16679 10047
rect 16962 10013 16996 10047
rect 17233 10013 17267 10047
rect 17969 10013 18003 10047
rect 18153 10013 18187 10047
rect 18429 10013 18463 10047
rect 23305 10013 23339 10047
rect 23581 10013 23615 10047
rect 23949 10013 23983 10047
rect 24041 10013 24075 10047
rect 8953 9945 8987 9979
rect 9153 9945 9187 9979
rect 9413 9945 9447 9979
rect 12541 9945 12575 9979
rect 12725 9945 12759 9979
rect 15117 9945 15151 9979
rect 16773 9945 16807 9979
rect 16865 9945 16899 9979
rect 17601 9945 17635 9979
rect 2605 9877 2639 9911
rect 7941 9877 7975 9911
rect 8401 9877 8435 9911
rect 8585 9877 8619 9911
rect 9597 9877 9631 9911
rect 9689 9877 9723 9911
rect 11069 9877 11103 9911
rect 13001 9877 13035 9911
rect 14657 9877 14691 9911
rect 15317 9877 15351 9911
rect 26157 9877 26191 9911
rect 5549 9673 5583 9707
rect 8769 9673 8803 9707
rect 15761 9673 15795 9707
rect 18337 9673 18371 9707
rect 18981 9673 19015 9707
rect 7481 9605 7515 9639
rect 8585 9605 8619 9639
rect 16221 9605 16255 9639
rect 20361 9605 20395 9639
rect 20821 9605 20855 9639
rect 20591 9571 20625 9605
rect 4077 9537 4111 9571
rect 4537 9537 4571 9571
rect 4721 9537 4755 9571
rect 5089 9537 5123 9571
rect 5365 9537 5399 9571
rect 7389 9537 7423 9571
rect 7573 9537 7607 9571
rect 8125 9537 8159 9571
rect 8309 9537 8343 9571
rect 8401 9537 8435 9571
rect 12817 9537 12851 9571
rect 12909 9537 12943 9571
rect 13001 9537 13035 9571
rect 13277 9537 13311 9571
rect 15117 9537 15151 9571
rect 15301 9537 15335 9571
rect 15393 9537 15427 9571
rect 15577 9537 15611 9571
rect 16129 9537 16163 9571
rect 16313 9537 16347 9571
rect 18153 9537 18187 9571
rect 18889 9537 18923 9571
rect 19073 9537 19107 9571
rect 21097 9537 21131 9571
rect 21557 9537 21591 9571
rect 24225 9537 24259 9571
rect 3985 9469 4019 9503
rect 4629 9469 4663 9503
rect 7941 9469 7975 9503
rect 17877 9469 17911 9503
rect 18245 9469 18279 9503
rect 18337 9469 18371 9503
rect 21373 9469 21407 9503
rect 4445 9401 4479 9435
rect 5181 9401 5215 9435
rect 5273 9401 5307 9435
rect 17969 9401 18003 9435
rect 20729 9401 20763 9435
rect 21281 9401 21315 9435
rect 12541 9333 12575 9367
rect 13093 9333 13127 9367
rect 14933 9333 14967 9367
rect 15393 9333 15427 9367
rect 20545 9333 20579 9367
rect 21189 9333 21223 9367
rect 24317 9333 24351 9367
rect 4445 9129 4479 9163
rect 8125 9129 8159 9163
rect 12449 9129 12483 9163
rect 13001 9129 13035 9163
rect 18521 9129 18555 9163
rect 21005 9129 21039 9163
rect 11989 9061 12023 9095
rect 3341 8993 3375 9027
rect 3617 8993 3651 9027
rect 4077 8993 4111 9027
rect 5181 8993 5215 9027
rect 10517 8993 10551 9027
rect 19257 8993 19291 9027
rect 3249 8925 3283 8959
rect 3985 8925 4019 8959
rect 4169 8925 4203 8959
rect 4261 8925 4295 8959
rect 5273 8925 5307 8959
rect 7941 8925 7975 8959
rect 8125 8925 8159 8959
rect 10241 8925 10275 8959
rect 12725 8925 12759 8959
rect 12817 8925 12851 8959
rect 18429 8925 18463 8959
rect 18521 8925 18555 8959
rect 19441 8925 19475 8959
rect 20729 8925 20763 8959
rect 20821 8925 20855 8959
rect 21005 8925 21039 8959
rect 23489 8925 23523 8959
rect 23673 8925 23707 8959
rect 23949 8925 23983 8959
rect 12357 8857 12391 8891
rect 18245 8857 18279 8891
rect 19625 8857 19659 8891
rect 5641 8789 5675 8823
rect 23765 8789 23799 8823
rect 3617 8585 3651 8619
rect 5457 8585 5491 8619
rect 7757 8585 7791 8619
rect 8033 8585 8067 8619
rect 10149 8585 10183 8619
rect 11897 8585 11931 8619
rect 17233 8585 17267 8619
rect 18245 8585 18279 8619
rect 23029 8585 23063 8619
rect 7205 8517 7239 8551
rect 10333 8517 10367 8551
rect 16681 8517 16715 8551
rect 16897 8517 16931 8551
rect 23305 8517 23339 8551
rect 24225 8517 24259 8551
rect 24945 8517 24979 8551
rect 25145 8517 25179 8551
rect 3065 8449 3099 8483
rect 3525 8449 3559 8483
rect 3709 8449 3743 8483
rect 3801 8449 3835 8483
rect 3985 8449 4019 8483
rect 5365 8449 5399 8483
rect 5549 8449 5583 8483
rect 7021 8449 7055 8483
rect 7113 8449 7147 8483
rect 7389 8449 7423 8483
rect 7481 8449 7515 8483
rect 7573 8449 7607 8483
rect 7757 8449 7791 8483
rect 7849 8449 7883 8483
rect 8033 8449 8067 8483
rect 9137 8449 9171 8483
rect 9321 8449 9355 8483
rect 10057 8449 10091 8483
rect 10701 8449 10735 8483
rect 10793 8449 10827 8483
rect 11805 8449 11839 8483
rect 11989 8449 12023 8483
rect 17141 8449 17175 8483
rect 17417 8449 17451 8483
rect 17877 8449 17911 8483
rect 23213 8449 23247 8483
rect 23397 8449 23431 8483
rect 23581 8449 23615 8483
rect 23949 8449 23983 8483
rect 24317 8449 24351 8483
rect 24501 8449 24535 8483
rect 25237 8449 25271 8483
rect 2973 8381 3007 8415
rect 7205 8381 7239 8415
rect 10425 8381 10459 8415
rect 17785 8381 17819 8415
rect 24133 8381 24167 8415
rect 3433 8313 3467 8347
rect 3893 8313 3927 8347
rect 6745 8313 6779 8347
rect 9229 8313 9263 8347
rect 10977 8313 11011 8347
rect 23765 8313 23799 8347
rect 24777 8313 24811 8347
rect 25421 8313 25455 8347
rect 7113 8245 7147 8279
rect 16865 8245 16899 8279
rect 17049 8245 17083 8279
rect 17417 8245 17451 8279
rect 24133 8245 24167 8279
rect 24685 8245 24719 8279
rect 24961 8245 24995 8279
rect 8493 8041 8527 8075
rect 9321 8041 9355 8075
rect 11989 8041 12023 8075
rect 12725 8041 12759 8075
rect 15393 8041 15427 8075
rect 15853 8041 15887 8075
rect 17233 8041 17267 8075
rect 24133 8041 24167 8075
rect 26157 8041 26191 8075
rect 4353 7973 4387 8007
rect 21281 7973 21315 8007
rect 3893 7905 3927 7939
rect 4721 7905 4755 7939
rect 6929 7905 6963 7939
rect 7389 7905 7423 7939
rect 11529 7905 11563 7939
rect 17049 7905 17083 7939
rect 19625 7905 19659 7939
rect 24409 7905 24443 7939
rect 24685 7905 24719 7939
rect 3985 7837 4019 7871
rect 4629 7837 4663 7871
rect 7021 7837 7055 7871
rect 8401 7837 8435 7871
rect 8585 7837 8619 7871
rect 8953 7837 8987 7871
rect 9137 7837 9171 7871
rect 11437 7837 11471 7871
rect 11713 7837 11747 7871
rect 11805 7837 11839 7871
rect 12909 7837 12943 7871
rect 13001 7837 13035 7871
rect 13185 7837 13219 7871
rect 13277 7837 13311 7871
rect 15393 7837 15427 7871
rect 15577 7837 15611 7871
rect 15669 7837 15703 7871
rect 16957 7837 16991 7871
rect 17233 7837 17267 7871
rect 18061 7837 18095 7871
rect 18153 7837 18187 7871
rect 18337 7837 18371 7871
rect 18429 7837 18463 7871
rect 18705 7837 18739 7871
rect 18883 7837 18917 7871
rect 19257 7837 19291 7871
rect 19441 7837 19475 7871
rect 19717 7837 19751 7871
rect 19809 7837 19843 7871
rect 20545 7837 20579 7871
rect 20637 7837 20671 7871
rect 20821 7837 20855 7871
rect 20913 7837 20947 7871
rect 21189 7837 21223 7871
rect 21373 7837 21407 7871
rect 21465 7837 21499 7871
rect 22845 7837 22879 7871
rect 23673 7837 23707 7871
rect 23857 7837 23891 7871
rect 23949 7837 23983 7871
rect 24133 7837 24167 7871
rect 18797 7769 18831 7803
rect 21741 7769 21775 7803
rect 22661 7769 22695 7803
rect 23305 7769 23339 7803
rect 4997 7701 5031 7735
rect 16773 7701 16807 7735
rect 18613 7701 18647 7735
rect 20361 7701 20395 7735
rect 21005 7701 21039 7735
rect 21833 7701 21867 7735
rect 23029 7701 23063 7735
rect 23489 7701 23523 7735
rect 4353 7497 4387 7531
rect 6469 7497 6503 7531
rect 11253 7497 11287 7531
rect 15669 7497 15703 7531
rect 17969 7497 18003 7531
rect 21005 7497 21039 7531
rect 21649 7497 21683 7531
rect 23029 7497 23063 7531
rect 23121 7497 23155 7531
rect 6653 7429 6687 7463
rect 6837 7429 6871 7463
rect 8677 7429 8711 7463
rect 9321 7429 9355 7463
rect 9781 7429 9815 7463
rect 11621 7429 11655 7463
rect 12173 7429 12207 7463
rect 12389 7429 12423 7463
rect 15231 7429 15265 7463
rect 16221 7429 16255 7463
rect 21833 7429 21867 7463
rect 22201 7429 22235 7463
rect 22753 7429 22787 7463
rect 22937 7429 22971 7463
rect 4169 7361 4203 7395
rect 4353 7361 4387 7395
rect 6377 7361 6411 7395
rect 6745 7361 6779 7395
rect 6929 7361 6963 7395
rect 8493 7361 8527 7395
rect 8861 7361 8895 7395
rect 8953 7361 8987 7395
rect 9137 7361 9171 7395
rect 9413 7361 9447 7395
rect 9597 7361 9631 7395
rect 10701 7361 10735 7395
rect 10793 7361 10827 7395
rect 10977 7361 11011 7395
rect 11069 7361 11103 7395
rect 11529 7361 11563 7395
rect 11713 7361 11747 7395
rect 11989 7361 12023 7395
rect 13001 7361 13035 7395
rect 14473 7361 14507 7395
rect 14749 7361 14783 7395
rect 14841 7361 14875 7395
rect 14933 7361 14967 7395
rect 15945 7361 15979 7395
rect 17417 7361 17451 7395
rect 17877 7361 17911 7395
rect 18613 7361 18647 7395
rect 18981 7361 19015 7395
rect 19901 7361 19935 7395
rect 20361 7361 20395 7395
rect 20453 7361 20487 7395
rect 20545 7361 20579 7395
rect 20729 7361 20763 7395
rect 20821 7361 20855 7395
rect 21281 7361 21315 7395
rect 22017 7361 22051 7395
rect 22293 7361 22327 7395
rect 22661 7361 22695 7395
rect 23765 7361 23799 7395
rect 24225 7361 24259 7395
rect 24317 7361 24351 7395
rect 14657 7293 14691 7327
rect 15117 7293 15151 7327
rect 15853 7293 15887 7327
rect 16313 7293 16347 7327
rect 18705 7293 18739 7327
rect 18889 7293 18923 7327
rect 21189 7293 21223 7327
rect 23397 7293 23431 7327
rect 23857 7293 23891 7327
rect 11897 7225 11931 7259
rect 15301 7225 15335 7259
rect 19625 7225 19659 7259
rect 19993 7225 20027 7259
rect 20085 7225 20119 7259
rect 22477 7225 22511 7259
rect 23305 7225 23339 7259
rect 6653 7157 6687 7191
rect 12357 7157 12391 7191
rect 12541 7157 12575 7191
rect 12909 7157 12943 7191
rect 14473 7157 14507 7191
rect 15025 7157 15059 7191
rect 17509 7157 17543 7191
rect 20177 7157 20211 7191
rect 24041 7157 24075 7191
rect 8677 6953 8711 6987
rect 9321 6953 9355 6987
rect 10425 6953 10459 6987
rect 10793 6953 10827 6987
rect 14289 6953 14323 6987
rect 18797 6953 18831 6987
rect 19441 6953 19475 6987
rect 20066 6953 20100 6987
rect 21557 6953 21591 6987
rect 21833 6953 21867 6987
rect 22740 6953 22774 6987
rect 24225 6953 24259 6987
rect 5457 6885 5491 6919
rect 7389 6885 7423 6919
rect 7849 6885 7883 6919
rect 15209 6885 15243 6919
rect 6009 6817 6043 6851
rect 6285 6817 6319 6851
rect 6377 6817 6411 6851
rect 6929 6817 6963 6851
rect 8953 6817 8987 6851
rect 11989 6817 12023 6851
rect 12541 6817 12575 6851
rect 12725 6817 12759 6851
rect 15945 6817 15979 6851
rect 16773 6817 16807 6851
rect 17233 6817 17267 6851
rect 17509 6817 17543 6851
rect 19809 6817 19843 6851
rect 22477 6817 22511 6851
rect 5181 6749 5215 6783
rect 5917 6749 5951 6783
rect 6561 6749 6595 6783
rect 6745 6749 6779 6783
rect 7021 6749 7055 6783
rect 8217 6749 8251 6783
rect 8401 6749 8435 6783
rect 8493 6749 8527 6783
rect 8677 6749 8711 6783
rect 9137 6749 9171 6783
rect 9413 6749 9447 6783
rect 9597 6749 9631 6783
rect 10425 6749 10459 6783
rect 10701 6749 10735 6783
rect 10977 6749 11011 6783
rect 11253 6749 11287 6783
rect 11529 6749 11563 6783
rect 11621 6749 11655 6783
rect 11805 6749 11839 6783
rect 11897 6749 11931 6783
rect 12081 6749 12115 6783
rect 12449 6749 12483 6783
rect 12817 6749 12851 6783
rect 13083 6743 13117 6777
rect 13185 6749 13219 6783
rect 13369 6749 13403 6783
rect 13461 6749 13495 6783
rect 14197 6749 14231 6783
rect 14473 6749 14507 6783
rect 14565 6749 14599 6783
rect 14933 6749 14967 6783
rect 15393 6749 15427 6783
rect 15485 6749 15519 6783
rect 15669 6749 15703 6783
rect 15761 6749 15795 6783
rect 15853 6749 15887 6783
rect 16681 6749 16715 6783
rect 17049 6749 17083 6783
rect 17325 6749 17359 6783
rect 17693 6749 17727 6783
rect 17785 6749 17819 6783
rect 17969 6749 18003 6783
rect 18061 6749 18095 6783
rect 18337 6749 18371 6783
rect 18613 6749 18647 6783
rect 18889 6749 18923 6783
rect 19441 6749 19475 6783
rect 19625 6749 19659 6783
rect 19717 6749 19751 6783
rect 22017 6749 22051 6783
rect 7573 6681 7607 6715
rect 8309 6681 8343 6715
rect 11161 6681 11195 6715
rect 13645 6681 13679 6715
rect 14749 6681 14783 6715
rect 14841 6681 14875 6715
rect 18521 6681 18555 6715
rect 5641 6613 5675 6647
rect 9505 6613 9539 6647
rect 10609 6613 10643 6647
rect 11345 6613 11379 6647
rect 15117 6613 15151 6647
rect 18153 6613 18187 6647
rect 6193 6409 6227 6443
rect 6561 6409 6595 6443
rect 11805 6409 11839 6443
rect 14841 6409 14875 6443
rect 15301 6409 15335 6443
rect 19165 6409 19199 6443
rect 21005 6409 21039 6443
rect 23029 6409 23063 6443
rect 27629 6409 27663 6443
rect 6929 6341 6963 6375
rect 12633 6341 12667 6375
rect 12817 6341 12851 6375
rect 14933 6341 14967 6375
rect 17693 6341 17727 6375
rect 5825 6273 5859 6307
rect 6469 6273 6503 6307
rect 6745 6273 6779 6307
rect 7297 6273 7331 6307
rect 12081 6273 12115 6307
rect 12265 6273 12299 6307
rect 12541 6273 12575 6307
rect 12909 6273 12943 6307
rect 13829 6273 13863 6307
rect 14461 6273 14495 6307
rect 15117 6273 15151 6307
rect 15393 6273 15427 6307
rect 21097 6273 21131 6307
rect 22937 6273 22971 6307
rect 27813 6273 27847 6307
rect 5917 6205 5951 6239
rect 7205 6205 7239 6239
rect 7665 6205 7699 6239
rect 13737 6205 13771 6239
rect 14565 6205 14599 6239
rect 17417 6205 17451 6239
rect 12173 6137 12207 6171
rect 12633 6137 12667 6171
rect 14197 6137 14231 6171
rect 12357 6069 12391 6103
rect 14657 6069 14691 6103
rect 11989 5865 12023 5899
rect 15853 5865 15887 5899
rect 17969 5865 18003 5899
rect 27629 5865 27663 5899
rect 10241 5729 10275 5763
rect 14105 5729 14139 5763
rect 16221 5729 16255 5763
rect 27813 5661 27847 5695
rect 10517 5593 10551 5627
rect 14381 5593 14415 5627
rect 16497 5593 16531 5627
rect 13277 5321 13311 5355
rect 11805 5253 11839 5287
rect 11529 5185 11563 5219
rect 6101 2601 6135 2635
rect 8677 2601 8711 2635
rect 5917 2397 5951 2431
rect 8493 2397 8527 2431
<< metal1 >>
rect 16758 28908 16764 28960
rect 16816 28948 16822 28960
rect 17494 28948 17500 28960
rect 16816 28920 17500 28948
rect 16816 28908 16822 28920
rect 17494 28908 17500 28920
rect 17552 28908 17558 28960
rect 1104 28858 28152 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 28152 28858
rect 1104 28784 28152 28806
rect 12894 28704 12900 28756
rect 12952 28744 12958 28756
rect 12989 28747 13047 28753
rect 12989 28744 13001 28747
rect 12952 28716 13001 28744
rect 12952 28704 12958 28716
rect 12989 28713 13001 28716
rect 13035 28713 13047 28747
rect 12989 28707 13047 28713
rect 13538 28704 13544 28756
rect 13596 28704 13602 28756
rect 14366 28704 14372 28756
rect 14424 28704 14430 28756
rect 14826 28704 14832 28756
rect 14884 28744 14890 28756
rect 15013 28747 15071 28753
rect 15013 28744 15025 28747
rect 14884 28716 15025 28744
rect 14884 28704 14890 28716
rect 15013 28713 15025 28716
rect 15059 28713 15071 28747
rect 15013 28707 15071 28713
rect 15654 28704 15660 28756
rect 15712 28704 15718 28756
rect 16114 28704 16120 28756
rect 16172 28744 16178 28756
rect 16761 28747 16819 28753
rect 16761 28744 16773 28747
rect 16172 28716 16773 28744
rect 16172 28704 16178 28716
rect 16761 28713 16773 28716
rect 16807 28713 16819 28747
rect 16761 28707 16819 28713
rect 17402 28704 17408 28756
rect 17460 28744 17466 28756
rect 17865 28747 17923 28753
rect 17865 28744 17877 28747
rect 17460 28716 17877 28744
rect 17460 28704 17466 28716
rect 17865 28713 17877 28716
rect 17911 28713 17923 28747
rect 17865 28707 17923 28713
rect 18046 28704 18052 28756
rect 18104 28744 18110 28756
rect 18509 28747 18567 28753
rect 18509 28744 18521 28747
rect 18104 28716 18521 28744
rect 18104 28704 18110 28716
rect 18509 28713 18521 28716
rect 18555 28713 18567 28747
rect 18509 28707 18567 28713
rect 19334 28704 19340 28756
rect 19392 28744 19398 28756
rect 19889 28747 19947 28753
rect 19889 28744 19901 28747
rect 19392 28716 19901 28744
rect 19392 28704 19398 28716
rect 19889 28713 19901 28716
rect 19935 28713 19947 28747
rect 19889 28707 19947 28713
rect 20622 28704 20628 28756
rect 20680 28744 20686 28756
rect 21085 28747 21143 28753
rect 21085 28744 21097 28747
rect 20680 28716 21097 28744
rect 20680 28704 20686 28716
rect 21085 28713 21097 28716
rect 21131 28713 21143 28747
rect 21085 28707 21143 28713
rect 21910 28704 21916 28756
rect 21968 28744 21974 28756
rect 21968 28716 22324 28744
rect 21968 28704 21974 28716
rect 17218 28636 17224 28688
rect 17276 28676 17282 28688
rect 17276 28648 17356 28676
rect 17276 28636 17282 28648
rect 15289 28543 15347 28549
rect 15289 28509 15301 28543
rect 15335 28540 15347 28543
rect 17126 28540 17132 28552
rect 15335 28512 17132 28540
rect 15335 28509 15347 28512
rect 15289 28503 15347 28509
rect 17126 28500 17132 28512
rect 17184 28500 17190 28552
rect 17328 28549 17356 28648
rect 17494 28636 17500 28688
rect 17552 28636 17558 28688
rect 18690 28636 18696 28688
rect 18748 28676 18754 28688
rect 19521 28679 19579 28685
rect 19521 28676 19533 28679
rect 18748 28648 19533 28676
rect 18748 28636 18754 28648
rect 19521 28645 19533 28648
rect 19567 28645 19579 28679
rect 19521 28639 19579 28645
rect 19978 28636 19984 28688
rect 20036 28676 20042 28688
rect 20717 28679 20775 28685
rect 20717 28676 20729 28679
rect 20036 28648 20729 28676
rect 20036 28636 20042 28648
rect 20717 28645 20729 28648
rect 20763 28645 20775 28679
rect 20717 28639 20775 28645
rect 21266 28636 21272 28688
rect 21324 28676 21330 28688
rect 22097 28679 22155 28685
rect 22097 28676 22109 28679
rect 21324 28648 22109 28676
rect 21324 28636 21330 28648
rect 22097 28645 22109 28648
rect 22143 28645 22155 28679
rect 22296 28676 22324 28716
rect 22554 28704 22560 28756
rect 22612 28744 22618 28756
rect 23109 28747 23167 28753
rect 23109 28744 23121 28747
rect 22612 28716 23121 28744
rect 22612 28704 22618 28716
rect 23109 28713 23121 28716
rect 23155 28713 23167 28747
rect 23109 28707 23167 28713
rect 23198 28704 23204 28756
rect 23256 28744 23262 28756
rect 23661 28747 23719 28753
rect 23661 28744 23673 28747
rect 23256 28716 23673 28744
rect 23256 28704 23262 28716
rect 23661 28713 23673 28716
rect 23707 28713 23719 28747
rect 23661 28707 23719 28713
rect 23842 28704 23848 28756
rect 23900 28744 23906 28756
rect 24581 28747 24639 28753
rect 24581 28744 24593 28747
rect 23900 28716 24593 28744
rect 23900 28704 23906 28716
rect 24581 28713 24593 28716
rect 24627 28713 24639 28747
rect 24581 28707 24639 28713
rect 25130 28704 25136 28756
rect 25188 28744 25194 28756
rect 25685 28747 25743 28753
rect 25685 28744 25697 28747
rect 25188 28716 25697 28744
rect 25188 28704 25194 28716
rect 25685 28713 25697 28716
rect 25731 28713 25743 28747
rect 25685 28707 25743 28713
rect 25774 28704 25780 28756
rect 25832 28744 25838 28756
rect 26145 28747 26203 28753
rect 26145 28744 26157 28747
rect 25832 28716 26157 28744
rect 25832 28704 25838 28716
rect 26145 28713 26157 28716
rect 26191 28713 26203 28747
rect 26145 28707 26203 28713
rect 26418 28704 26424 28756
rect 26476 28744 26482 28756
rect 27157 28747 27215 28753
rect 27157 28744 27169 28747
rect 26476 28716 27169 28744
rect 26476 28704 26482 28716
rect 27157 28713 27169 28716
rect 27203 28713 27215 28747
rect 27157 28707 27215 28713
rect 22649 28679 22707 28685
rect 22649 28676 22661 28679
rect 22296 28648 22661 28676
rect 22097 28639 22155 28645
rect 22649 28645 22661 28648
rect 22695 28645 22707 28679
rect 22649 28639 22707 28645
rect 24486 28636 24492 28688
rect 24544 28676 24550 28688
rect 25225 28679 25283 28685
rect 25225 28676 25237 28679
rect 24544 28648 25237 28676
rect 24544 28636 24550 28648
rect 25225 28645 25237 28648
rect 25271 28645 25283 28679
rect 25225 28639 25283 28645
rect 17313 28543 17371 28549
rect 17313 28509 17325 28543
rect 17359 28509 17371 28543
rect 17313 28503 17371 28509
rect 26050 28500 26056 28552
rect 26108 28540 26114 28552
rect 27065 28543 27123 28549
rect 27065 28540 27077 28543
rect 26108 28512 27077 28540
rect 26108 28500 26114 28512
rect 27065 28509 27077 28512
rect 27111 28509 27123 28543
rect 27065 28503 27123 28509
rect 13262 28432 13268 28484
rect 13320 28432 13326 28484
rect 13817 28475 13875 28481
rect 13817 28441 13829 28475
rect 13863 28441 13875 28475
rect 13817 28435 13875 28441
rect 13832 28404 13860 28435
rect 14642 28432 14648 28484
rect 14700 28432 14706 28484
rect 15933 28475 15991 28481
rect 15933 28441 15945 28475
rect 15979 28472 15991 28475
rect 16850 28472 16856 28484
rect 15979 28444 16856 28472
rect 15979 28441 15991 28444
rect 15933 28435 15991 28441
rect 16850 28432 16856 28444
rect 16908 28432 16914 28484
rect 17037 28475 17095 28481
rect 17037 28441 17049 28475
rect 17083 28472 17095 28475
rect 17083 28444 18092 28472
rect 17083 28441 17095 28444
rect 17037 28435 17095 28441
rect 17770 28404 17776 28416
rect 13832 28376 17776 28404
rect 17770 28364 17776 28376
rect 17828 28364 17834 28416
rect 18064 28404 18092 28444
rect 18138 28432 18144 28484
rect 18196 28432 18202 28484
rect 18414 28432 18420 28484
rect 18472 28432 18478 28484
rect 19334 28432 19340 28484
rect 19392 28432 19398 28484
rect 20070 28432 20076 28484
rect 20128 28472 20134 28484
rect 20165 28475 20223 28481
rect 20165 28472 20177 28475
rect 20128 28444 20177 28472
rect 20128 28432 20134 28444
rect 20165 28441 20177 28444
rect 20211 28441 20223 28475
rect 20165 28435 20223 28441
rect 20438 28432 20444 28484
rect 20496 28432 20502 28484
rect 20990 28432 20996 28484
rect 21048 28432 21054 28484
rect 21450 28432 21456 28484
rect 21508 28472 21514 28484
rect 21913 28475 21971 28481
rect 21913 28472 21925 28475
rect 21508 28444 21925 28472
rect 21508 28432 21514 28444
rect 21913 28441 21925 28444
rect 21959 28441 21971 28475
rect 21913 28435 21971 28441
rect 22462 28432 22468 28484
rect 22520 28432 22526 28484
rect 23014 28432 23020 28484
rect 23072 28432 23078 28484
rect 23106 28432 23112 28484
rect 23164 28472 23170 28484
rect 23569 28475 23627 28481
rect 23569 28472 23581 28475
rect 23164 28444 23581 28472
rect 23164 28432 23170 28444
rect 23569 28441 23581 28444
rect 23615 28441 23627 28475
rect 23569 28435 23627 28441
rect 24486 28432 24492 28484
rect 24544 28432 24550 28484
rect 25038 28432 25044 28484
rect 25096 28432 25102 28484
rect 25590 28432 25596 28484
rect 25648 28432 25654 28484
rect 26418 28432 26424 28484
rect 26476 28432 26482 28484
rect 22002 28404 22008 28416
rect 18064 28376 22008 28404
rect 22002 28364 22008 28376
rect 22060 28364 22066 28416
rect 1104 28314 28152 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 28152 28314
rect 1104 28240 28152 28262
rect 18049 28203 18107 28209
rect 18049 28169 18061 28203
rect 18095 28200 18107 28203
rect 18414 28200 18420 28212
rect 18095 28172 18420 28200
rect 18095 28169 18107 28172
rect 18049 28163 18107 28169
rect 18414 28160 18420 28172
rect 18472 28160 18478 28212
rect 19061 28203 19119 28209
rect 19061 28200 19073 28203
rect 18524 28172 19073 28200
rect 10134 28092 10140 28144
rect 10192 28132 10198 28144
rect 10192 28104 11928 28132
rect 10192 28092 10198 28104
rect 6362 28024 6368 28076
rect 6420 28064 6426 28076
rect 6825 28067 6883 28073
rect 6825 28064 6837 28067
rect 6420 28036 6837 28064
rect 6420 28024 6426 28036
rect 6825 28033 6837 28036
rect 6871 28033 6883 28067
rect 6825 28027 6883 28033
rect 6914 28024 6920 28076
rect 6972 28064 6978 28076
rect 7009 28067 7067 28073
rect 7009 28064 7021 28067
rect 6972 28036 7021 28064
rect 6972 28024 6978 28036
rect 7009 28033 7021 28036
rect 7055 28033 7067 28067
rect 7009 28027 7067 28033
rect 10962 28024 10968 28076
rect 11020 28024 11026 28076
rect 11790 28064 11796 28076
rect 11072 28036 11796 28064
rect 9398 27956 9404 28008
rect 9456 27996 9462 28008
rect 11072 27996 11100 28036
rect 11790 28024 11796 28036
rect 11848 28024 11854 28076
rect 11900 28073 11928 28104
rect 13262 28092 13268 28144
rect 13320 28132 13326 28144
rect 18524 28132 18552 28172
rect 19061 28169 19073 28172
rect 19107 28169 19119 28203
rect 19978 28200 19984 28212
rect 19061 28163 19119 28169
rect 19168 28172 19984 28200
rect 19168 28132 19196 28172
rect 19978 28160 19984 28172
rect 20036 28160 20042 28212
rect 20070 28160 20076 28212
rect 20128 28160 20134 28212
rect 20165 28203 20223 28209
rect 20165 28169 20177 28203
rect 20211 28200 20223 28203
rect 20438 28200 20444 28212
rect 20211 28172 20444 28200
rect 20211 28169 20223 28172
rect 20165 28163 20223 28169
rect 20438 28160 20444 28172
rect 20496 28160 20502 28212
rect 22373 28203 22431 28209
rect 22373 28169 22385 28203
rect 22419 28200 22431 28203
rect 23014 28200 23020 28212
rect 22419 28172 23020 28200
rect 22419 28169 22431 28172
rect 22373 28163 22431 28169
rect 23014 28160 23020 28172
rect 23072 28160 23078 28212
rect 27062 28160 27068 28212
rect 27120 28200 27126 28212
rect 27341 28203 27399 28209
rect 27341 28200 27353 28203
rect 27120 28172 27353 28200
rect 27120 28160 27126 28172
rect 27341 28169 27353 28172
rect 27387 28169 27399 28203
rect 27341 28163 27399 28169
rect 13320 28104 18552 28132
rect 19076 28104 19196 28132
rect 19229 28135 19287 28141
rect 13320 28092 13326 28104
rect 11885 28067 11943 28073
rect 11885 28033 11897 28067
rect 11931 28064 11943 28067
rect 12250 28064 12256 28076
rect 11931 28036 12256 28064
rect 11931 28033 11943 28036
rect 11885 28027 11943 28033
rect 12250 28024 12256 28036
rect 12308 28024 12314 28076
rect 17954 28024 17960 28076
rect 18012 28024 18018 28076
rect 18141 28067 18199 28073
rect 18141 28033 18153 28067
rect 18187 28064 18199 28067
rect 19076 28064 19104 28104
rect 19229 28101 19241 28135
rect 19275 28101 19287 28135
rect 19229 28095 19287 28101
rect 18187 28036 19104 28064
rect 18187 28033 18199 28036
rect 18141 28027 18199 28033
rect 9456 27968 11100 27996
rect 11241 27999 11299 28005
rect 9456 27956 9462 27968
rect 11241 27965 11253 27999
rect 11287 27996 11299 27999
rect 12066 27996 12072 28008
rect 11287 27968 12072 27996
rect 11287 27965 11299 27968
rect 11241 27959 11299 27965
rect 12066 27956 12072 27968
rect 12124 27956 12130 28008
rect 17586 27956 17592 28008
rect 17644 27996 17650 28008
rect 18156 27996 18184 28027
rect 17644 27968 18184 27996
rect 17644 27956 17650 27968
rect 19150 27956 19156 28008
rect 19208 27996 19214 28008
rect 19244 27996 19272 28095
rect 19426 28092 19432 28144
rect 19484 28092 19490 28144
rect 19521 28135 19579 28141
rect 19521 28101 19533 28135
rect 19567 28132 19579 28135
rect 19610 28132 19616 28144
rect 19567 28104 19616 28132
rect 19567 28101 19579 28104
rect 19521 28095 19579 28101
rect 19610 28092 19616 28104
rect 19668 28092 19674 28144
rect 20317 28135 20375 28141
rect 20317 28101 20329 28135
rect 20363 28132 20375 28135
rect 20533 28135 20591 28141
rect 20363 28101 20392 28132
rect 20317 28095 20392 28101
rect 20533 28101 20545 28135
rect 20579 28132 20591 28135
rect 20898 28132 20904 28144
rect 20579 28104 20904 28132
rect 20579 28101 20591 28104
rect 20533 28095 20591 28101
rect 19702 28024 19708 28076
rect 19760 28024 19766 28076
rect 19794 28024 19800 28076
rect 19852 28024 19858 28076
rect 19889 28067 19947 28073
rect 19889 28033 19901 28067
rect 19935 28064 19947 28067
rect 20364 28064 20392 28095
rect 20898 28092 20904 28104
rect 20956 28092 20962 28144
rect 21910 28132 21916 28144
rect 21100 28104 21916 28132
rect 21100 28073 21128 28104
rect 21910 28092 21916 28104
rect 21968 28132 21974 28144
rect 22189 28135 22247 28141
rect 22189 28132 22201 28135
rect 21968 28104 22201 28132
rect 21968 28092 21974 28104
rect 22189 28101 22201 28104
rect 22235 28101 22247 28135
rect 22189 28095 22247 28101
rect 25961 28135 26019 28141
rect 25961 28101 25973 28135
rect 26007 28132 26019 28135
rect 27249 28135 27307 28141
rect 27249 28132 27261 28135
rect 26007 28104 27261 28132
rect 26007 28101 26019 28104
rect 25961 28095 26019 28101
rect 27249 28101 27261 28104
rect 27295 28101 27307 28135
rect 27249 28095 27307 28101
rect 21085 28067 21143 28073
rect 21085 28064 21097 28067
rect 19935 28036 21097 28064
rect 19935 28033 19947 28036
rect 19889 28027 19947 28033
rect 21085 28033 21097 28036
rect 21131 28033 21143 28067
rect 21085 28027 21143 28033
rect 21174 28024 21180 28076
rect 21232 28024 21238 28076
rect 22005 28067 22063 28073
rect 22005 28033 22017 28067
rect 22051 28033 22063 28067
rect 22005 28027 22063 28033
rect 22097 28067 22155 28073
rect 22097 28033 22109 28067
rect 22143 28064 22155 28067
rect 22370 28064 22376 28076
rect 22143 28036 22376 28064
rect 22143 28033 22155 28036
rect 22097 28027 22155 28033
rect 19208 27968 19748 27996
rect 19208 27956 19214 27968
rect 19058 27888 19064 27940
rect 19116 27928 19122 27940
rect 19426 27928 19432 27940
rect 19116 27900 19432 27928
rect 19116 27888 19122 27900
rect 19426 27888 19432 27900
rect 19484 27888 19490 27940
rect 6454 27820 6460 27872
rect 6512 27860 6518 27872
rect 7006 27860 7012 27872
rect 6512 27832 7012 27860
rect 6512 27820 6518 27832
rect 7006 27820 7012 27832
rect 7064 27820 7070 27872
rect 10226 27820 10232 27872
rect 10284 27860 10290 27872
rect 10781 27863 10839 27869
rect 10781 27860 10793 27863
rect 10284 27832 10793 27860
rect 10284 27820 10290 27832
rect 10781 27829 10793 27832
rect 10827 27829 10839 27863
rect 10781 27823 10839 27829
rect 10870 27820 10876 27872
rect 10928 27860 10934 27872
rect 11149 27863 11207 27869
rect 11149 27860 11161 27863
rect 10928 27832 11161 27860
rect 10928 27820 10934 27832
rect 11149 27829 11161 27832
rect 11195 27829 11207 27863
rect 11149 27823 11207 27829
rect 11698 27820 11704 27872
rect 11756 27820 11762 27872
rect 19245 27863 19303 27869
rect 19245 27829 19257 27863
rect 19291 27860 19303 27863
rect 19610 27860 19616 27872
rect 19291 27832 19616 27860
rect 19291 27829 19303 27832
rect 19245 27823 19303 27829
rect 19610 27820 19616 27832
rect 19668 27820 19674 27872
rect 19720 27860 19748 27968
rect 19978 27956 19984 28008
rect 20036 27996 20042 28008
rect 21192 27996 21220 28024
rect 20036 27968 21220 27996
rect 22020 27996 22048 28027
rect 22370 28024 22376 28036
rect 22428 28024 22434 28076
rect 24578 28024 24584 28076
rect 24636 28064 24642 28076
rect 24673 28067 24731 28073
rect 24673 28064 24685 28067
rect 24636 28036 24685 28064
rect 24636 28024 24642 28036
rect 24673 28033 24685 28036
rect 24719 28033 24731 28067
rect 24673 28027 24731 28033
rect 24762 28024 24768 28076
rect 24820 28064 24826 28076
rect 25133 28067 25191 28073
rect 25133 28064 25145 28067
rect 24820 28036 25145 28064
rect 24820 28024 24826 28036
rect 25133 28033 25145 28036
rect 25179 28033 25191 28067
rect 25133 28027 25191 28033
rect 25774 28024 25780 28076
rect 25832 28064 25838 28076
rect 25869 28067 25927 28073
rect 25869 28064 25881 28067
rect 25832 28036 25881 28064
rect 25832 28024 25838 28036
rect 25869 28033 25881 28036
rect 25915 28033 25927 28067
rect 25869 28027 25927 28033
rect 26053 28067 26111 28073
rect 26053 28033 26065 28067
rect 26099 28033 26111 28067
rect 26053 28027 26111 28033
rect 24394 27996 24400 28008
rect 22020 27968 24400 27996
rect 20036 27956 20042 27968
rect 24394 27956 24400 27968
rect 24452 27956 24458 28008
rect 25041 27999 25099 28005
rect 25041 27965 25053 27999
rect 25087 27996 25099 27999
rect 25222 27996 25228 28008
rect 25087 27968 25228 27996
rect 25087 27965 25099 27968
rect 25041 27959 25099 27965
rect 25222 27956 25228 27968
rect 25280 27956 25286 28008
rect 19886 27888 19892 27940
rect 19944 27928 19950 27940
rect 20622 27928 20628 27940
rect 19944 27900 20628 27928
rect 19944 27888 19950 27900
rect 20622 27888 20628 27900
rect 20680 27928 20686 27940
rect 21821 27931 21879 27937
rect 21821 27928 21833 27931
rect 20680 27900 21833 27928
rect 20680 27888 20686 27900
rect 21821 27897 21833 27900
rect 21867 27897 21879 27931
rect 21821 27891 21879 27897
rect 25130 27888 25136 27940
rect 25188 27928 25194 27940
rect 26068 27928 26096 28027
rect 26326 28024 26332 28076
rect 26384 28064 26390 28076
rect 26421 28067 26479 28073
rect 26421 28064 26433 28067
rect 26384 28036 26433 28064
rect 26384 28024 26390 28036
rect 26421 28033 26433 28036
rect 26467 28033 26479 28067
rect 26421 28027 26479 28033
rect 26789 28067 26847 28073
rect 26789 28033 26801 28067
rect 26835 28064 26847 28067
rect 28994 28064 29000 28076
rect 26835 28036 29000 28064
rect 26835 28033 26847 28036
rect 26789 28027 26847 28033
rect 28994 28024 29000 28036
rect 29052 28024 29058 28076
rect 26142 27928 26148 27940
rect 25188 27900 26148 27928
rect 25188 27888 25194 27900
rect 26142 27888 26148 27900
rect 26200 27888 26206 27940
rect 20349 27863 20407 27869
rect 20349 27860 20361 27863
rect 19720 27832 20361 27860
rect 20349 27829 20361 27832
rect 20395 27829 20407 27863
rect 20349 27823 20407 27829
rect 24854 27820 24860 27872
rect 24912 27820 24918 27872
rect 25314 27820 25320 27872
rect 25372 27820 25378 27872
rect 1104 27770 28152 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 28152 27770
rect 1104 27696 28152 27718
rect 5629 27659 5687 27665
rect 5629 27625 5641 27659
rect 5675 27625 5687 27659
rect 5629 27619 5687 27625
rect 2746 27560 5396 27588
rect 2222 27480 2228 27532
rect 2280 27520 2286 27532
rect 2746 27520 2774 27560
rect 2280 27492 2774 27520
rect 5077 27523 5135 27529
rect 2280 27480 2286 27492
rect 5077 27489 5089 27523
rect 5123 27520 5135 27523
rect 5258 27520 5264 27532
rect 5123 27492 5264 27520
rect 5123 27489 5135 27492
rect 5077 27483 5135 27489
rect 5258 27480 5264 27492
rect 5316 27480 5322 27532
rect 5368 27520 5396 27560
rect 5442 27548 5448 27600
rect 5500 27588 5506 27600
rect 5644 27588 5672 27619
rect 6362 27616 6368 27668
rect 6420 27656 6426 27668
rect 10413 27659 10471 27665
rect 6420 27628 7696 27656
rect 6420 27616 6426 27628
rect 6914 27588 6920 27600
rect 5500 27560 5672 27588
rect 5736 27560 6920 27588
rect 5500 27548 5506 27560
rect 5736 27520 5764 27560
rect 6914 27548 6920 27560
rect 6972 27588 6978 27600
rect 7668 27588 7696 27628
rect 10413 27625 10425 27659
rect 10459 27656 10471 27659
rect 10870 27656 10876 27668
rect 10459 27628 10876 27656
rect 10459 27625 10471 27628
rect 10413 27619 10471 27625
rect 10870 27616 10876 27628
rect 10928 27616 10934 27668
rect 11057 27659 11115 27665
rect 11057 27625 11069 27659
rect 11103 27656 11115 27659
rect 11238 27656 11244 27668
rect 11103 27628 11244 27656
rect 11103 27625 11115 27628
rect 11057 27619 11115 27625
rect 11238 27616 11244 27628
rect 11296 27616 11302 27668
rect 11790 27616 11796 27668
rect 11848 27656 11854 27668
rect 11848 27628 12434 27656
rect 11848 27616 11854 27628
rect 10134 27588 10140 27600
rect 6972 27560 7604 27588
rect 6972 27548 6978 27560
rect 7009 27523 7067 27529
rect 5368 27492 5764 27520
rect 5828 27492 6960 27520
rect 3789 27455 3847 27461
rect 3789 27421 3801 27455
rect 3835 27452 3847 27455
rect 3878 27452 3884 27464
rect 3835 27424 3884 27452
rect 3835 27421 3847 27424
rect 3789 27415 3847 27421
rect 3878 27412 3884 27424
rect 3936 27412 3942 27464
rect 3970 27412 3976 27464
rect 4028 27412 4034 27464
rect 4798 27412 4804 27464
rect 4856 27452 4862 27464
rect 4985 27455 5043 27461
rect 4985 27452 4997 27455
rect 4856 27424 4997 27452
rect 4856 27412 4862 27424
rect 4985 27421 4997 27424
rect 5031 27421 5043 27455
rect 5828 27452 5856 27492
rect 4985 27415 5043 27421
rect 5092 27424 5856 27452
rect 6089 27455 6147 27461
rect 3694 27344 3700 27396
rect 3752 27384 3758 27396
rect 5092 27384 5120 27424
rect 6089 27421 6101 27455
rect 6135 27452 6147 27455
rect 6178 27452 6184 27464
rect 6135 27424 6184 27452
rect 6135 27421 6147 27424
rect 6089 27415 6147 27421
rect 6178 27412 6184 27424
rect 6236 27412 6242 27464
rect 6273 27455 6331 27461
rect 6273 27421 6285 27455
rect 6319 27452 6331 27455
rect 6454 27452 6460 27464
rect 6319 27424 6460 27452
rect 6319 27421 6331 27424
rect 6273 27415 6331 27421
rect 6454 27412 6460 27424
rect 6512 27412 6518 27464
rect 6546 27412 6552 27464
rect 6604 27452 6610 27464
rect 6932 27461 6960 27492
rect 7009 27489 7021 27523
rect 7055 27520 7067 27523
rect 7377 27523 7435 27529
rect 7377 27520 7389 27523
rect 7055 27492 7389 27520
rect 7055 27489 7067 27492
rect 7009 27483 7067 27489
rect 7377 27489 7389 27492
rect 7423 27489 7435 27523
rect 7377 27483 7435 27489
rect 7576 27461 7604 27560
rect 7668 27560 10140 27588
rect 6641 27455 6699 27461
rect 6641 27452 6653 27455
rect 6604 27424 6653 27452
rect 6604 27412 6610 27424
rect 6641 27421 6653 27424
rect 6687 27421 6699 27455
rect 6641 27415 6699 27421
rect 6917 27455 6975 27461
rect 6917 27421 6929 27455
rect 6963 27452 6975 27455
rect 7561 27455 7619 27461
rect 6963 27424 7512 27452
rect 6963 27421 6975 27424
rect 6917 27415 6975 27421
rect 5445 27387 5503 27393
rect 5445 27384 5457 27387
rect 3752 27356 5120 27384
rect 5184 27356 5457 27384
rect 3752 27344 3758 27356
rect 3881 27319 3939 27325
rect 3881 27285 3893 27319
rect 3927 27316 3939 27319
rect 4062 27316 4068 27328
rect 3927 27288 4068 27316
rect 3927 27285 3939 27288
rect 3881 27279 3939 27285
rect 4062 27276 4068 27288
rect 4120 27276 4126 27328
rect 4706 27276 4712 27328
rect 4764 27316 4770 27328
rect 5184 27316 5212 27356
rect 5445 27353 5457 27356
rect 5491 27384 5503 27387
rect 5994 27384 6000 27396
rect 5491 27356 6000 27384
rect 5491 27353 5503 27356
rect 5445 27347 5503 27353
rect 5994 27344 6000 27356
rect 6052 27344 6058 27396
rect 4764 27288 5212 27316
rect 5353 27319 5411 27325
rect 4764 27276 4770 27288
rect 5353 27285 5365 27319
rect 5399 27316 5411 27319
rect 5534 27316 5540 27328
rect 5399 27288 5540 27316
rect 5399 27285 5411 27288
rect 5353 27279 5411 27285
rect 5534 27276 5540 27288
rect 5592 27316 5598 27328
rect 5645 27319 5703 27325
rect 5645 27316 5657 27319
rect 5592 27288 5657 27316
rect 5592 27276 5598 27288
rect 5645 27285 5657 27288
rect 5691 27285 5703 27319
rect 5645 27279 5703 27285
rect 5810 27276 5816 27328
rect 5868 27276 5874 27328
rect 6086 27276 6092 27328
rect 6144 27276 6150 27328
rect 6454 27276 6460 27328
rect 6512 27316 6518 27328
rect 6549 27319 6607 27325
rect 6549 27316 6561 27319
rect 6512 27288 6561 27316
rect 6512 27276 6518 27288
rect 6549 27285 6561 27288
rect 6595 27285 6607 27319
rect 6549 27279 6607 27285
rect 7285 27319 7343 27325
rect 7285 27285 7297 27319
rect 7331 27316 7343 27319
rect 7374 27316 7380 27328
rect 7331 27288 7380 27316
rect 7331 27285 7343 27288
rect 7285 27279 7343 27285
rect 7374 27276 7380 27288
rect 7432 27276 7438 27328
rect 7484 27316 7512 27424
rect 7561 27421 7573 27455
rect 7607 27421 7619 27455
rect 7668 27452 7696 27560
rect 9968 27529 9996 27560
rect 10134 27548 10140 27560
rect 10192 27548 10198 27600
rect 10318 27548 10324 27600
rect 10376 27548 10382 27600
rect 12406 27588 12434 27628
rect 17218 27616 17224 27668
rect 17276 27616 17282 27668
rect 18138 27616 18144 27668
rect 18196 27656 18202 27668
rect 18233 27659 18291 27665
rect 18233 27656 18245 27659
rect 18196 27628 18245 27656
rect 18196 27616 18202 27628
rect 18233 27625 18245 27628
rect 18279 27625 18291 27659
rect 18233 27619 18291 27625
rect 18969 27659 19027 27665
rect 18969 27625 18981 27659
rect 19015 27656 19027 27659
rect 19058 27656 19064 27668
rect 19015 27628 19064 27656
rect 19015 27625 19027 27628
rect 18969 27619 19027 27625
rect 19058 27616 19064 27628
rect 19116 27616 19122 27668
rect 19168 27628 19380 27656
rect 10888 27560 11836 27588
rect 12406 27560 12480 27588
rect 9677 27523 9735 27529
rect 9677 27489 9689 27523
rect 9723 27489 9735 27523
rect 9677 27483 9735 27489
rect 9953 27523 10011 27529
rect 9953 27489 9965 27523
rect 9999 27489 10011 27523
rect 9953 27483 10011 27489
rect 7837 27455 7895 27461
rect 7837 27452 7849 27455
rect 7668 27424 7849 27452
rect 7561 27415 7619 27421
rect 7837 27421 7849 27424
rect 7883 27421 7895 27455
rect 7837 27415 7895 27421
rect 7576 27384 7604 27415
rect 7926 27412 7932 27464
rect 7984 27452 7990 27464
rect 8021 27455 8079 27461
rect 8021 27452 8033 27455
rect 7984 27424 8033 27452
rect 7984 27412 7990 27424
rect 8021 27421 8033 27424
rect 8067 27452 8079 27455
rect 9398 27452 9404 27464
rect 8067 27424 9404 27452
rect 8067 27421 8079 27424
rect 8021 27415 8079 27421
rect 9398 27412 9404 27424
rect 9456 27412 9462 27464
rect 9585 27455 9643 27461
rect 9585 27421 9597 27455
rect 9631 27421 9643 27455
rect 9692 27452 9720 27483
rect 10778 27480 10784 27532
rect 10836 27480 10842 27532
rect 10226 27452 10232 27464
rect 9692 27424 10232 27452
rect 9585 27415 9643 27421
rect 7576 27356 9444 27384
rect 8294 27316 8300 27328
rect 7484 27288 8300 27316
rect 8294 27276 8300 27288
rect 8352 27276 8358 27328
rect 9217 27319 9275 27325
rect 9217 27285 9229 27319
rect 9263 27316 9275 27319
rect 9306 27316 9312 27328
rect 9263 27288 9312 27316
rect 9263 27285 9275 27288
rect 9217 27279 9275 27285
rect 9306 27276 9312 27288
rect 9364 27276 9370 27328
rect 9416 27316 9444 27356
rect 9490 27344 9496 27396
rect 9548 27384 9554 27396
rect 9600 27384 9628 27415
rect 10226 27412 10232 27424
rect 10284 27412 10290 27464
rect 10888 27461 10916 27560
rect 11808 27520 11836 27560
rect 11072 27492 11560 27520
rect 11808 27492 11928 27520
rect 10597 27455 10655 27461
rect 10597 27421 10609 27455
rect 10643 27421 10655 27455
rect 10597 27415 10655 27421
rect 10689 27455 10747 27461
rect 10689 27421 10701 27455
rect 10735 27421 10747 27455
rect 10689 27415 10747 27421
rect 10873 27455 10931 27461
rect 10873 27421 10885 27455
rect 10919 27421 10931 27455
rect 10873 27415 10931 27421
rect 9548 27356 9628 27384
rect 9548 27344 9554 27356
rect 10612 27316 10640 27415
rect 10704 27384 10732 27415
rect 11072 27384 11100 27492
rect 11149 27455 11207 27461
rect 11149 27421 11161 27455
rect 11195 27421 11207 27455
rect 11149 27415 11207 27421
rect 10704 27356 11100 27384
rect 11164 27316 11192 27415
rect 11330 27412 11336 27464
rect 11388 27412 11394 27464
rect 11532 27461 11560 27492
rect 11517 27455 11575 27461
rect 11517 27421 11529 27455
rect 11563 27452 11575 27455
rect 11698 27452 11704 27464
rect 11563 27424 11704 27452
rect 11563 27421 11575 27424
rect 11517 27415 11575 27421
rect 11698 27412 11704 27424
rect 11756 27412 11762 27464
rect 11790 27412 11796 27464
rect 11848 27412 11854 27464
rect 11900 27461 11928 27492
rect 11885 27455 11943 27461
rect 11885 27421 11897 27455
rect 11931 27452 11943 27455
rect 12069 27455 12127 27461
rect 12069 27452 12081 27455
rect 11931 27424 12081 27452
rect 11931 27421 11943 27424
rect 11885 27415 11943 27421
rect 12069 27421 12081 27424
rect 12115 27452 12127 27455
rect 12158 27452 12164 27464
rect 12115 27424 12164 27452
rect 12115 27421 12127 27424
rect 12069 27415 12127 27421
rect 12158 27412 12164 27424
rect 12216 27412 12222 27464
rect 12250 27412 12256 27464
rect 12308 27461 12314 27464
rect 12452 27461 12480 27560
rect 17126 27548 17132 27600
rect 17184 27588 17190 27600
rect 17497 27591 17555 27597
rect 17497 27588 17509 27591
rect 17184 27560 17509 27588
rect 17184 27548 17190 27560
rect 17497 27557 17509 27560
rect 17543 27557 17555 27591
rect 17497 27551 17555 27557
rect 17770 27548 17776 27600
rect 17828 27548 17834 27600
rect 19168 27588 19196 27628
rect 18616 27560 19196 27588
rect 19245 27591 19303 27597
rect 17236 27492 17540 27520
rect 17236 27461 17264 27492
rect 17512 27461 17540 27492
rect 17696 27492 18276 27520
rect 12308 27455 12341 27461
rect 12329 27421 12341 27455
rect 12308 27415 12341 27421
rect 12437 27455 12495 27461
rect 12437 27421 12449 27455
rect 12483 27452 12495 27455
rect 17221 27455 17279 27461
rect 12483 27424 12848 27452
rect 12483 27421 12495 27424
rect 12437 27415 12495 27421
rect 12308 27412 12314 27415
rect 11808 27384 11836 27412
rect 12820 27396 12848 27424
rect 17221 27421 17233 27455
rect 17267 27421 17279 27455
rect 17221 27415 17279 27421
rect 17405 27455 17463 27461
rect 17405 27421 17417 27455
rect 17451 27421 17463 27455
rect 17405 27415 17463 27421
rect 17497 27455 17555 27461
rect 17497 27421 17509 27455
rect 17543 27452 17555 27455
rect 17586 27452 17592 27464
rect 17543 27424 17592 27452
rect 17543 27421 17555 27424
rect 17497 27415 17555 27421
rect 12529 27387 12587 27393
rect 12529 27384 12541 27387
rect 11808 27356 12541 27384
rect 12529 27353 12541 27356
rect 12575 27353 12587 27387
rect 12529 27347 12587 27353
rect 12713 27387 12771 27393
rect 12713 27353 12725 27387
rect 12759 27353 12771 27387
rect 12713 27347 12771 27353
rect 11882 27316 11888 27328
rect 9416 27288 11888 27316
rect 11882 27276 11888 27288
rect 11940 27276 11946 27328
rect 11974 27276 11980 27328
rect 12032 27316 12038 27328
rect 12728 27316 12756 27347
rect 12802 27344 12808 27396
rect 12860 27384 12866 27396
rect 12897 27387 12955 27393
rect 12897 27384 12909 27387
rect 12860 27356 12909 27384
rect 12860 27344 12866 27356
rect 12897 27353 12909 27356
rect 12943 27353 12955 27387
rect 17420 27384 17448 27415
rect 17586 27412 17592 27424
rect 17644 27412 17650 27464
rect 17696 27461 17724 27492
rect 17681 27455 17739 27461
rect 17681 27421 17693 27455
rect 17727 27421 17739 27455
rect 17681 27415 17739 27421
rect 17773 27455 17831 27461
rect 17773 27421 17785 27455
rect 17819 27452 17831 27455
rect 17862 27452 17868 27464
rect 17819 27424 17868 27452
rect 17819 27421 17831 27424
rect 17773 27415 17831 27421
rect 17862 27412 17868 27424
rect 17920 27412 17926 27464
rect 17957 27455 18015 27461
rect 17957 27421 17969 27455
rect 18003 27452 18015 27455
rect 18046 27452 18052 27464
rect 18003 27424 18052 27452
rect 18003 27421 18015 27424
rect 17957 27415 18015 27421
rect 18046 27412 18052 27424
rect 18104 27412 18110 27464
rect 18248 27461 18276 27492
rect 18616 27461 18644 27560
rect 19245 27557 19257 27591
rect 19291 27557 19303 27591
rect 19245 27551 19303 27557
rect 19260 27520 19288 27551
rect 18708 27492 19288 27520
rect 18233 27455 18291 27461
rect 18233 27421 18245 27455
rect 18279 27452 18291 27455
rect 18601 27455 18659 27461
rect 18279 27424 18552 27452
rect 18279 27421 18291 27424
rect 18233 27415 18291 27421
rect 18524 27384 18552 27424
rect 18601 27421 18613 27455
rect 18647 27421 18659 27455
rect 18601 27415 18659 27421
rect 18708 27384 18736 27492
rect 18785 27455 18843 27461
rect 18785 27421 18797 27455
rect 18831 27452 18843 27455
rect 19061 27455 19119 27461
rect 18831 27424 18920 27452
rect 18831 27421 18843 27424
rect 18785 27415 18843 27421
rect 17420 27356 18460 27384
rect 18524 27356 18736 27384
rect 12897 27347 12955 27353
rect 12986 27316 12992 27328
rect 12032 27288 12992 27316
rect 12032 27276 12038 27288
rect 12986 27276 12992 27288
rect 13044 27276 13050 27328
rect 18230 27276 18236 27328
rect 18288 27316 18294 27328
rect 18432 27325 18460 27356
rect 18417 27319 18475 27325
rect 18417 27316 18429 27319
rect 18288 27288 18429 27316
rect 18288 27276 18294 27288
rect 18417 27285 18429 27288
rect 18463 27285 18475 27319
rect 18892 27316 18920 27424
rect 19061 27421 19073 27455
rect 19107 27421 19119 27455
rect 19352 27452 19380 27628
rect 19426 27616 19432 27668
rect 19484 27616 19490 27668
rect 20809 27659 20867 27665
rect 20809 27625 20821 27659
rect 20855 27656 20867 27659
rect 20990 27656 20996 27668
rect 20855 27628 20996 27656
rect 20855 27625 20867 27628
rect 20809 27619 20867 27625
rect 20990 27616 20996 27628
rect 21048 27616 21054 27668
rect 21269 27659 21327 27665
rect 21269 27625 21281 27659
rect 21315 27656 21327 27659
rect 21913 27659 21971 27665
rect 21913 27656 21925 27659
rect 21315 27628 21925 27656
rect 21315 27625 21327 27628
rect 21269 27619 21327 27625
rect 21913 27625 21925 27628
rect 21959 27656 21971 27659
rect 22097 27659 22155 27665
rect 21959 27628 22048 27656
rect 21959 27625 21971 27628
rect 21913 27619 21971 27625
rect 19886 27588 19892 27600
rect 19720 27560 19892 27588
rect 19518 27480 19524 27532
rect 19576 27480 19582 27532
rect 19429 27455 19487 27461
rect 19429 27452 19441 27455
rect 19352 27424 19441 27452
rect 19061 27415 19119 27421
rect 19429 27421 19441 27424
rect 19475 27452 19487 27455
rect 19720 27452 19748 27560
rect 19886 27548 19892 27560
rect 19944 27548 19950 27600
rect 19978 27548 19984 27600
rect 20036 27548 20042 27600
rect 20070 27548 20076 27600
rect 20128 27588 20134 27600
rect 20128 27560 20944 27588
rect 20128 27548 20134 27560
rect 19794 27480 19800 27532
rect 19852 27520 19858 27532
rect 19852 27492 20116 27520
rect 19852 27480 19858 27492
rect 19475 27424 19748 27452
rect 20088 27452 20116 27492
rect 20162 27480 20168 27532
rect 20220 27520 20226 27532
rect 20220 27492 20668 27520
rect 20220 27480 20226 27492
rect 20257 27455 20315 27461
rect 20257 27452 20269 27455
rect 20088 27424 20269 27452
rect 19475 27421 19487 27424
rect 19429 27415 19487 27421
rect 20257 27421 20269 27424
rect 20303 27452 20315 27455
rect 20346 27452 20352 27464
rect 20303 27424 20352 27452
rect 20303 27421 20315 27424
rect 20257 27415 20315 27421
rect 19076 27384 19104 27415
rect 20346 27412 20352 27424
rect 20404 27412 20410 27464
rect 20640 27461 20668 27492
rect 20916 27461 20944 27560
rect 21450 27548 21456 27600
rect 21508 27548 21514 27600
rect 22020 27588 22048 27628
rect 22097 27625 22109 27659
rect 22143 27656 22155 27659
rect 22462 27656 22468 27668
rect 22143 27628 22468 27656
rect 22143 27625 22155 27628
rect 22097 27619 22155 27625
rect 22462 27616 22468 27628
rect 22520 27616 22526 27668
rect 23477 27659 23535 27665
rect 23477 27625 23489 27659
rect 23523 27656 23535 27659
rect 24486 27656 24492 27668
rect 23523 27628 24492 27656
rect 23523 27625 23535 27628
rect 23477 27619 23535 27625
rect 24486 27616 24492 27628
rect 24544 27616 24550 27668
rect 24578 27616 24584 27668
rect 24636 27656 24642 27668
rect 24857 27659 24915 27665
rect 24857 27656 24869 27659
rect 24636 27628 24869 27656
rect 24636 27616 24642 27628
rect 24857 27625 24869 27628
rect 24903 27656 24915 27659
rect 24946 27656 24952 27668
rect 24903 27628 24952 27656
rect 24903 27625 24915 27628
rect 24857 27619 24915 27625
rect 24946 27616 24952 27628
rect 25004 27616 25010 27668
rect 25130 27616 25136 27668
rect 25188 27616 25194 27668
rect 25498 27616 25504 27668
rect 25556 27656 25562 27668
rect 25685 27659 25743 27665
rect 25685 27656 25697 27659
rect 25556 27628 25697 27656
rect 25556 27616 25562 27628
rect 25685 27625 25697 27628
rect 25731 27625 25743 27659
rect 25685 27619 25743 27625
rect 26329 27659 26387 27665
rect 26329 27625 26341 27659
rect 26375 27656 26387 27659
rect 26418 27656 26424 27668
rect 26375 27628 26424 27656
rect 26375 27625 26387 27628
rect 26329 27619 26387 27625
rect 26418 27616 26424 27628
rect 26476 27616 26482 27668
rect 23017 27591 23075 27597
rect 22020 27560 22692 27588
rect 20625 27455 20683 27461
rect 20625 27421 20637 27455
rect 20671 27421 20683 27455
rect 20625 27415 20683 27421
rect 20809 27455 20867 27461
rect 20809 27421 20821 27455
rect 20855 27421 20867 27455
rect 20809 27415 20867 27421
rect 20901 27455 20959 27461
rect 20901 27421 20913 27455
rect 20947 27452 20959 27455
rect 21545 27455 21603 27461
rect 21545 27452 21557 27455
rect 20947 27424 21557 27452
rect 20947 27421 20959 27424
rect 20901 27415 20959 27421
rect 21545 27421 21557 27424
rect 21591 27452 21603 27455
rect 21634 27452 21640 27464
rect 21591 27424 21640 27452
rect 21591 27421 21603 27424
rect 21545 27415 21603 27421
rect 19518 27384 19524 27396
rect 19076 27356 19524 27384
rect 19518 27344 19524 27356
rect 19576 27344 19582 27396
rect 19794 27344 19800 27396
rect 19852 27384 19858 27396
rect 19889 27387 19947 27393
rect 19889 27384 19901 27387
rect 19852 27356 19901 27384
rect 19852 27344 19858 27356
rect 19889 27353 19901 27356
rect 19935 27384 19947 27387
rect 20070 27384 20076 27396
rect 19935 27356 20076 27384
rect 19935 27353 19947 27356
rect 19889 27347 19947 27353
rect 20070 27344 20076 27356
rect 20128 27344 20134 27396
rect 20180 27356 20484 27384
rect 20180 27328 20208 27356
rect 19426 27316 19432 27328
rect 18892 27288 19432 27316
rect 18417 27279 18475 27285
rect 19426 27276 19432 27288
rect 19484 27276 19490 27328
rect 20162 27276 20168 27328
rect 20220 27276 20226 27328
rect 20254 27276 20260 27328
rect 20312 27316 20318 27328
rect 20349 27319 20407 27325
rect 20349 27316 20361 27319
rect 20312 27288 20361 27316
rect 20312 27276 20318 27288
rect 20349 27285 20361 27288
rect 20395 27285 20407 27319
rect 20456 27316 20484 27356
rect 20530 27344 20536 27396
rect 20588 27344 20594 27396
rect 20824 27384 20852 27415
rect 21634 27412 21640 27424
rect 21692 27412 21698 27464
rect 22373 27455 22431 27461
rect 22373 27421 22385 27455
rect 22419 27452 22431 27455
rect 22554 27452 22560 27464
rect 22419 27424 22560 27452
rect 22419 27421 22431 27424
rect 22373 27415 22431 27421
rect 22554 27412 22560 27424
rect 22612 27412 22618 27464
rect 22664 27452 22692 27560
rect 23017 27557 23029 27591
rect 23063 27588 23075 27591
rect 23106 27588 23112 27600
rect 23063 27560 23112 27588
rect 23063 27557 23075 27560
rect 23017 27551 23075 27557
rect 23106 27548 23112 27560
rect 23164 27548 23170 27600
rect 24213 27591 24271 27597
rect 24213 27557 24225 27591
rect 24259 27588 24271 27591
rect 25038 27588 25044 27600
rect 24259 27560 25044 27588
rect 24259 27557 24271 27560
rect 24213 27551 24271 27557
rect 25038 27548 25044 27560
rect 25096 27548 25102 27600
rect 27706 27548 27712 27600
rect 27764 27548 27770 27600
rect 22741 27523 22799 27529
rect 22741 27489 22753 27523
rect 22787 27520 22799 27523
rect 24854 27520 24860 27532
rect 22787 27492 23336 27520
rect 22787 27489 22799 27492
rect 22741 27483 22799 27489
rect 23308 27464 23336 27492
rect 24228 27492 24860 27520
rect 23201 27455 23259 27461
rect 23201 27452 23213 27455
rect 22664 27424 23213 27452
rect 23201 27421 23213 27424
rect 23247 27421 23259 27455
rect 23201 27415 23259 27421
rect 21174 27384 21180 27396
rect 20824 27356 21180 27384
rect 21174 27344 21180 27356
rect 21232 27384 21238 27396
rect 21232 27356 21404 27384
rect 21232 27344 21238 27356
rect 21269 27319 21327 27325
rect 21269 27316 21281 27319
rect 20456 27288 21281 27316
rect 20349 27279 20407 27285
rect 21269 27285 21281 27288
rect 21315 27285 21327 27319
rect 21376 27316 21404 27356
rect 21910 27344 21916 27396
rect 21968 27344 21974 27396
rect 22858 27387 22916 27393
rect 22066 27356 22784 27384
rect 22066 27316 22094 27356
rect 21376 27288 22094 27316
rect 21269 27279 21327 27285
rect 22646 27276 22652 27328
rect 22704 27276 22710 27328
rect 22756 27316 22784 27356
rect 22858 27353 22870 27387
rect 22904 27384 22916 27387
rect 23014 27384 23020 27396
rect 22904 27356 23020 27384
rect 22904 27353 22916 27356
rect 22858 27347 22916 27353
rect 23014 27344 23020 27356
rect 23072 27344 23078 27396
rect 23216 27384 23244 27415
rect 23290 27412 23296 27464
rect 23348 27412 23354 27464
rect 24026 27412 24032 27464
rect 24084 27412 24090 27464
rect 24228 27461 24256 27492
rect 24854 27480 24860 27492
rect 24912 27520 24918 27532
rect 24912 27492 26096 27520
rect 24912 27480 24918 27492
rect 24213 27455 24271 27461
rect 24213 27421 24225 27455
rect 24259 27421 24271 27455
rect 24213 27415 24271 27421
rect 24486 27412 24492 27464
rect 24544 27412 24550 27464
rect 24581 27455 24639 27461
rect 24581 27421 24593 27455
rect 24627 27452 24639 27455
rect 24762 27452 24768 27464
rect 24627 27424 24768 27452
rect 24627 27421 24639 27424
rect 24581 27415 24639 27421
rect 23382 27384 23388 27396
rect 23216 27356 23388 27384
rect 23382 27344 23388 27356
rect 23440 27344 23446 27396
rect 24302 27344 24308 27396
rect 24360 27384 24366 27396
rect 24596 27384 24624 27415
rect 24762 27412 24768 27424
rect 24820 27412 24826 27464
rect 24949 27455 25007 27461
rect 24949 27421 24961 27455
rect 24995 27421 25007 27455
rect 24949 27415 25007 27421
rect 24360 27356 24624 27384
rect 24964 27384 24992 27415
rect 25038 27412 25044 27464
rect 25096 27452 25102 27464
rect 25317 27455 25375 27461
rect 25317 27452 25329 27455
rect 25096 27424 25329 27452
rect 25096 27412 25102 27424
rect 25317 27421 25329 27424
rect 25363 27421 25375 27455
rect 25317 27415 25375 27421
rect 25406 27412 25412 27464
rect 25464 27412 25470 27464
rect 26068 27461 26096 27492
rect 26142 27480 26148 27532
rect 26200 27520 26206 27532
rect 26200 27492 26556 27520
rect 26200 27480 26206 27492
rect 25777 27455 25835 27461
rect 25777 27421 25789 27455
rect 25823 27421 25835 27455
rect 25777 27415 25835 27421
rect 26053 27455 26111 27461
rect 26053 27421 26065 27455
rect 26099 27421 26111 27455
rect 26053 27415 26111 27421
rect 25792 27384 25820 27415
rect 26234 27412 26240 27464
rect 26292 27452 26298 27464
rect 26528 27461 26556 27492
rect 26329 27455 26387 27461
rect 26329 27452 26341 27455
rect 26292 27424 26341 27452
rect 26292 27412 26298 27424
rect 26329 27421 26341 27424
rect 26375 27421 26387 27455
rect 26329 27415 26387 27421
rect 26513 27455 26571 27461
rect 26513 27421 26525 27455
rect 26559 27421 26571 27455
rect 27433 27455 27491 27461
rect 27433 27452 27445 27455
rect 26513 27415 26571 27421
rect 26988 27424 27445 27452
rect 24964 27356 25820 27384
rect 24360 27344 24366 27356
rect 25148 27328 25176 27356
rect 25866 27344 25872 27396
rect 25924 27384 25930 27396
rect 26881 27387 26939 27393
rect 26881 27384 26893 27387
rect 25924 27356 26893 27384
rect 25924 27344 25930 27356
rect 26881 27353 26893 27356
rect 26927 27353 26939 27387
rect 26881 27347 26939 27353
rect 24946 27316 24952 27328
rect 22756 27288 24952 27316
rect 24946 27276 24952 27288
rect 25004 27276 25010 27328
rect 25130 27276 25136 27328
rect 25188 27276 25194 27328
rect 25958 27276 25964 27328
rect 26016 27276 26022 27328
rect 26145 27319 26203 27325
rect 26145 27285 26157 27319
rect 26191 27316 26203 27319
rect 26988 27316 27016 27424
rect 27433 27421 27445 27424
rect 27479 27421 27491 27455
rect 27433 27415 27491 27421
rect 27249 27387 27307 27393
rect 27249 27353 27261 27387
rect 27295 27384 27307 27387
rect 28350 27384 28356 27396
rect 27295 27356 28356 27384
rect 27295 27353 27307 27356
rect 27249 27347 27307 27353
rect 28350 27344 28356 27356
rect 28408 27344 28414 27396
rect 26191 27288 27016 27316
rect 26191 27285 26203 27288
rect 26145 27279 26203 27285
rect 1104 27226 28152 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 28152 27226
rect 1104 27152 28152 27174
rect 3513 27115 3571 27121
rect 3513 27081 3525 27115
rect 3559 27112 3571 27115
rect 3970 27112 3976 27124
rect 3559 27084 3976 27112
rect 3559 27081 3571 27084
rect 3513 27075 3571 27081
rect 3970 27072 3976 27084
rect 4028 27072 4034 27124
rect 5258 27072 5264 27124
rect 5316 27072 5322 27124
rect 5718 27112 5724 27124
rect 5368 27084 5724 27112
rect 3142 27004 3148 27056
rect 3200 27004 3206 27056
rect 3345 27047 3403 27053
rect 3345 27044 3357 27047
rect 3252 27016 3357 27044
rect 2222 26936 2228 26988
rect 2280 26976 2286 26988
rect 2409 26979 2467 26985
rect 2409 26976 2421 26979
rect 2280 26948 2421 26976
rect 2280 26936 2286 26948
rect 2409 26945 2421 26948
rect 2455 26945 2467 26979
rect 3252 26976 3280 27016
rect 3345 27013 3357 27016
rect 3391 27044 3403 27047
rect 3881 27047 3939 27053
rect 3881 27044 3893 27047
rect 3391 27016 3893 27044
rect 3391 27013 3403 27016
rect 3345 27007 3403 27013
rect 3881 27013 3893 27016
rect 3927 27013 3939 27047
rect 5368 27044 5396 27084
rect 5718 27072 5724 27084
rect 5776 27112 5782 27124
rect 6365 27115 6423 27121
rect 6365 27112 6377 27115
rect 5776 27084 6377 27112
rect 5776 27072 5782 27084
rect 6365 27081 6377 27084
rect 6411 27081 6423 27115
rect 6914 27112 6920 27124
rect 6365 27075 6423 27081
rect 6656 27084 6920 27112
rect 5626 27044 5632 27056
rect 3881 27007 3939 27013
rect 5184 27016 5396 27044
rect 5460 27016 5632 27044
rect 3605 26979 3663 26985
rect 3605 26976 3617 26979
rect 2409 26939 2467 26945
rect 2792 26948 3280 26976
rect 3344 26948 3617 26976
rect 1854 26868 1860 26920
rect 1912 26908 1918 26920
rect 2314 26908 2320 26920
rect 1912 26880 2320 26908
rect 1912 26868 1918 26880
rect 2314 26868 2320 26880
rect 2372 26868 2378 26920
rect 2792 26917 2820 26948
rect 2777 26911 2835 26917
rect 2777 26877 2789 26911
rect 2823 26877 2835 26911
rect 2777 26871 2835 26877
rect 2866 26732 2872 26784
rect 2924 26772 2930 26784
rect 3344 26781 3372 26948
rect 3605 26945 3617 26948
rect 3651 26945 3663 26979
rect 3605 26939 3663 26945
rect 3694 26936 3700 26988
rect 3752 26936 3758 26988
rect 4062 26936 4068 26988
rect 4120 26936 4126 26988
rect 4433 26979 4491 26985
rect 4433 26945 4445 26979
rect 4479 26976 4491 26979
rect 4614 26976 4620 26988
rect 4479 26948 4620 26976
rect 4479 26945 4491 26948
rect 4433 26939 4491 26945
rect 4614 26936 4620 26948
rect 4672 26936 4678 26988
rect 5184 26985 5212 27016
rect 5169 26979 5227 26985
rect 5169 26945 5181 26979
rect 5215 26945 5227 26979
rect 5169 26939 5227 26945
rect 5353 26979 5411 26985
rect 5353 26945 5365 26979
rect 5399 26976 5411 26979
rect 5460 26976 5488 27016
rect 5626 27004 5632 27016
rect 5684 27004 5690 27056
rect 5810 27004 5816 27056
rect 5868 27004 5874 27056
rect 5399 26948 5488 26976
rect 5536 26979 5594 26985
rect 5399 26945 5411 26948
rect 5353 26939 5411 26945
rect 5536 26945 5548 26979
rect 5582 26974 5594 26979
rect 5828 26976 5856 27004
rect 5644 26974 5856 26976
rect 5582 26948 5856 26974
rect 5582 26946 5672 26948
rect 5582 26945 5594 26946
rect 5536 26939 5594 26945
rect 5994 26936 6000 26988
rect 6052 26976 6058 26988
rect 6546 26976 6552 26988
rect 6052 26948 6552 26976
rect 6052 26936 6058 26948
rect 6546 26936 6552 26948
rect 6604 26936 6610 26988
rect 6656 26985 6684 27084
rect 6914 27072 6920 27084
rect 6972 27072 6978 27124
rect 7929 27115 7987 27121
rect 7208 27084 7788 27112
rect 6641 26979 6699 26985
rect 6641 26945 6653 26979
rect 6687 26945 6699 26979
rect 6641 26939 6699 26945
rect 6730 26936 6736 26988
rect 6788 26976 6794 26988
rect 6917 26979 6975 26985
rect 6917 26976 6929 26979
rect 6788 26948 6929 26976
rect 6788 26936 6794 26948
rect 6917 26945 6929 26948
rect 6963 26976 6975 26979
rect 7208 26976 7236 27084
rect 7285 27047 7343 27053
rect 7285 27013 7297 27047
rect 7331 27044 7343 27047
rect 7331 27016 7696 27044
rect 7331 27013 7343 27016
rect 7285 27007 7343 27013
rect 6963 26948 7236 26976
rect 6963 26945 6975 26948
rect 6917 26939 6975 26945
rect 7374 26936 7380 26988
rect 7432 26976 7438 26988
rect 7469 26979 7527 26985
rect 7469 26976 7481 26979
rect 7432 26948 7481 26976
rect 7432 26936 7438 26948
rect 7469 26945 7481 26948
rect 7515 26945 7527 26979
rect 7469 26939 7527 26945
rect 5077 26911 5135 26917
rect 5077 26877 5089 26911
rect 5123 26908 5135 26911
rect 5258 26908 5264 26920
rect 5123 26880 5264 26908
rect 5123 26877 5135 26880
rect 5077 26871 5135 26877
rect 5258 26868 5264 26880
rect 5316 26868 5322 26920
rect 5629 26911 5687 26917
rect 5629 26908 5641 26911
rect 5552 26880 5641 26908
rect 4798 26800 4804 26852
rect 4856 26840 4862 26852
rect 5552 26840 5580 26880
rect 5629 26877 5641 26880
rect 5675 26877 5687 26911
rect 5629 26871 5687 26877
rect 5718 26868 5724 26920
rect 5776 26868 5782 26920
rect 5813 26911 5871 26917
rect 5813 26877 5825 26911
rect 5859 26908 5871 26911
rect 6086 26908 6092 26920
rect 5859 26880 6092 26908
rect 5859 26877 5871 26880
rect 5813 26871 5871 26877
rect 4856 26812 5580 26840
rect 4856 26800 4862 26812
rect 3329 26775 3387 26781
rect 3329 26772 3341 26775
rect 2924 26744 3341 26772
rect 2924 26732 2930 26744
rect 3329 26741 3341 26744
rect 3375 26741 3387 26775
rect 3329 26735 3387 26741
rect 3878 26732 3884 26784
rect 3936 26732 3942 26784
rect 5718 26732 5724 26784
rect 5776 26772 5782 26784
rect 5828 26772 5856 26871
rect 6086 26868 6092 26880
rect 6144 26868 6150 26920
rect 6362 26868 6368 26920
rect 6420 26868 6426 26920
rect 7006 26868 7012 26920
rect 7064 26908 7070 26920
rect 7193 26911 7251 26917
rect 7193 26908 7205 26911
rect 7064 26880 7205 26908
rect 7064 26868 7070 26880
rect 7193 26877 7205 26880
rect 7239 26908 7251 26911
rect 7561 26911 7619 26917
rect 7561 26908 7573 26911
rect 7239 26880 7573 26908
rect 7239 26877 7251 26880
rect 7193 26871 7251 26877
rect 7561 26877 7573 26880
rect 7607 26877 7619 26911
rect 7668 26908 7696 27016
rect 7760 26985 7788 27084
rect 7929 27081 7941 27115
rect 7975 27112 7987 27115
rect 10689 27115 10747 27121
rect 7975 27084 8248 27112
rect 7975 27081 7987 27084
rect 7929 27075 7987 27081
rect 7745 26979 7803 26985
rect 7745 26945 7757 26979
rect 7791 26976 7803 26979
rect 7926 26976 7932 26988
rect 7791 26948 7932 26976
rect 7791 26945 7803 26948
rect 7745 26939 7803 26945
rect 7926 26936 7932 26948
rect 7984 26936 7990 26988
rect 8220 26985 8248 27084
rect 10689 27081 10701 27115
rect 10735 27112 10747 27115
rect 10962 27112 10968 27124
rect 10735 27084 10968 27112
rect 10735 27081 10747 27084
rect 10689 27075 10747 27081
rect 10962 27072 10968 27084
rect 11020 27112 11026 27124
rect 11517 27115 11575 27121
rect 11517 27112 11529 27115
rect 11020 27084 11529 27112
rect 11020 27072 11026 27084
rect 11517 27081 11529 27084
rect 11563 27081 11575 27115
rect 11517 27075 11575 27081
rect 12066 27072 12072 27124
rect 12124 27112 12130 27124
rect 12161 27115 12219 27121
rect 12161 27112 12173 27115
rect 12124 27084 12173 27112
rect 12124 27072 12130 27084
rect 12161 27081 12173 27084
rect 12207 27081 12219 27115
rect 12161 27075 12219 27081
rect 16850 27072 16856 27124
rect 16908 27112 16914 27124
rect 17865 27115 17923 27121
rect 17865 27112 17877 27115
rect 16908 27084 17877 27112
rect 16908 27072 16914 27084
rect 17865 27081 17877 27084
rect 17911 27081 17923 27115
rect 17865 27075 17923 27081
rect 18325 27115 18383 27121
rect 18325 27081 18337 27115
rect 18371 27112 18383 27115
rect 19334 27112 19340 27124
rect 18371 27084 19340 27112
rect 18371 27081 18383 27084
rect 18325 27075 18383 27081
rect 19334 27072 19340 27084
rect 19392 27072 19398 27124
rect 19610 27072 19616 27124
rect 19668 27112 19674 27124
rect 20162 27112 20168 27124
rect 19668 27084 20168 27112
rect 19668 27072 19674 27084
rect 20162 27072 20168 27084
rect 20220 27112 20226 27124
rect 20257 27115 20315 27121
rect 20257 27112 20269 27115
rect 20220 27084 20269 27112
rect 20220 27072 20226 27084
rect 20257 27081 20269 27084
rect 20303 27081 20315 27115
rect 20257 27075 20315 27081
rect 8294 27004 8300 27056
rect 8352 27044 8358 27056
rect 11149 27047 11207 27053
rect 8352 27016 11100 27044
rect 8352 27004 8358 27016
rect 8021 26979 8079 26985
rect 8021 26945 8033 26979
rect 8067 26945 8079 26979
rect 8021 26939 8079 26945
rect 8205 26979 8263 26985
rect 8205 26945 8217 26979
rect 8251 26976 8263 26979
rect 9122 26976 9128 26988
rect 8251 26948 9128 26976
rect 8251 26945 8263 26948
rect 8205 26939 8263 26945
rect 8036 26908 8064 26939
rect 9122 26936 9128 26948
rect 9180 26936 9186 26988
rect 10045 26979 10103 26985
rect 10045 26945 10057 26979
rect 10091 26976 10103 26979
rect 10594 26976 10600 26988
rect 10091 26948 10600 26976
rect 10091 26945 10103 26948
rect 10045 26939 10103 26945
rect 10594 26936 10600 26948
rect 10652 26976 10658 26988
rect 10965 26979 11023 26985
rect 10965 26976 10977 26979
rect 10652 26948 10977 26976
rect 10652 26936 10658 26948
rect 10965 26945 10977 26948
rect 11011 26945 11023 26979
rect 10965 26939 11023 26945
rect 7668 26880 8064 26908
rect 7561 26871 7619 26877
rect 10226 26868 10232 26920
rect 10284 26868 10290 26920
rect 10321 26911 10379 26917
rect 10321 26877 10333 26911
rect 10367 26877 10379 26911
rect 10321 26871 10379 26877
rect 6546 26800 6552 26852
rect 6604 26840 6610 26852
rect 10336 26840 10364 26871
rect 6604 26812 10364 26840
rect 6604 26800 6610 26812
rect 5776 26744 5856 26772
rect 5776 26732 5782 26744
rect 5994 26732 6000 26784
rect 6052 26732 6058 26784
rect 6914 26732 6920 26784
rect 6972 26772 6978 26784
rect 7055 26775 7113 26781
rect 7055 26772 7067 26775
rect 6972 26744 7067 26772
rect 6972 26732 6978 26744
rect 7055 26741 7067 26744
rect 7101 26772 7113 26775
rect 7469 26775 7527 26781
rect 7469 26772 7481 26775
rect 7101 26744 7481 26772
rect 7101 26741 7113 26744
rect 7055 26735 7113 26741
rect 7469 26741 7481 26744
rect 7515 26741 7527 26775
rect 7469 26735 7527 26741
rect 8113 26775 8171 26781
rect 8113 26741 8125 26775
rect 8159 26772 8171 26775
rect 8202 26772 8208 26784
rect 8159 26744 8208 26772
rect 8159 26741 8171 26744
rect 8113 26735 8171 26741
rect 8202 26732 8208 26744
rect 8260 26732 8266 26784
rect 10686 26732 10692 26784
rect 10744 26772 10750 26784
rect 10781 26775 10839 26781
rect 10781 26772 10793 26775
rect 10744 26744 10793 26772
rect 10744 26732 10750 26744
rect 10781 26741 10793 26744
rect 10827 26741 10839 26775
rect 11072 26772 11100 27016
rect 11149 27013 11161 27047
rect 11195 27044 11207 27047
rect 11330 27044 11336 27056
rect 11195 27016 11336 27044
rect 11195 27013 11207 27016
rect 11149 27007 11207 27013
rect 11330 27004 11336 27016
rect 11388 27004 11394 27056
rect 12313 27047 12371 27053
rect 12313 27044 12325 27047
rect 12084 27016 12325 27044
rect 11238 26936 11244 26988
rect 11296 26936 11302 26988
rect 11698 26936 11704 26988
rect 11756 26936 11762 26988
rect 11882 26936 11888 26988
rect 11940 26976 11946 26988
rect 12084 26985 12112 27016
rect 12313 27013 12325 27016
rect 12359 27013 12371 27047
rect 12313 27007 12371 27013
rect 12526 27004 12532 27056
rect 12584 27044 12590 27056
rect 12805 27047 12863 27053
rect 12805 27044 12817 27047
rect 12584 27016 12817 27044
rect 12584 27004 12590 27016
rect 12805 27013 12817 27016
rect 12851 27013 12863 27047
rect 18877 27047 18935 27053
rect 18877 27044 18889 27047
rect 12805 27007 12863 27013
rect 17788 27016 18889 27044
rect 12069 26979 12127 26985
rect 12069 26976 12081 26979
rect 11940 26948 12081 26976
rect 11940 26936 11946 26948
rect 12069 26945 12081 26948
rect 12115 26945 12127 26979
rect 12069 26939 12127 26945
rect 12158 26936 12164 26988
rect 12216 26976 12222 26988
rect 17788 26985 17816 27016
rect 18877 27013 18889 27016
rect 18923 27044 18935 27047
rect 18966 27044 18972 27056
rect 18923 27016 18972 27044
rect 18923 27013 18935 27016
rect 18877 27007 18935 27013
rect 18966 27004 18972 27016
rect 19024 27004 19030 27056
rect 19794 27044 19800 27056
rect 19306 27016 19800 27044
rect 19306 26988 19334 27016
rect 19794 27004 19800 27016
rect 19852 27004 19858 27056
rect 19889 27047 19947 27053
rect 19889 27013 19901 27047
rect 19935 27044 19947 27047
rect 20272 27044 20300 27075
rect 22002 27072 22008 27124
rect 22060 27072 22066 27124
rect 22189 27115 22247 27121
rect 22189 27081 22201 27115
rect 22235 27112 22247 27115
rect 23290 27112 23296 27124
rect 22235 27084 23296 27112
rect 22235 27081 22247 27084
rect 22189 27075 22247 27081
rect 21177 27047 21235 27053
rect 19935 27016 20208 27044
rect 20272 27016 20760 27044
rect 19935 27013 19947 27016
rect 19889 27007 19947 27013
rect 20180 26988 20208 27016
rect 12621 26979 12679 26985
rect 12621 26976 12633 26979
rect 12216 26948 12633 26976
rect 12216 26936 12222 26948
rect 12621 26945 12633 26948
rect 12667 26945 12679 26979
rect 12621 26939 12679 26945
rect 17773 26979 17831 26985
rect 17773 26945 17785 26979
rect 17819 26945 17831 26979
rect 17773 26939 17831 26945
rect 17957 26979 18015 26985
rect 17957 26945 17969 26979
rect 18003 26976 18015 26979
rect 18046 26976 18052 26988
rect 18003 26948 18052 26976
rect 18003 26945 18015 26948
rect 17957 26939 18015 26945
rect 17972 26908 18000 26939
rect 18046 26936 18052 26948
rect 18104 26936 18110 26988
rect 18230 26936 18236 26988
rect 18288 26936 18294 26988
rect 18417 26979 18475 26985
rect 18417 26945 18429 26979
rect 18463 26945 18475 26979
rect 19150 26976 19156 26988
rect 19111 26948 19156 26976
rect 18417 26939 18475 26945
rect 18432 26908 18460 26939
rect 19150 26936 19156 26948
rect 19208 26936 19214 26988
rect 19242 26936 19248 26988
rect 19300 26948 19334 26988
rect 19300 26936 19306 26948
rect 19518 26936 19524 26988
rect 19576 26936 19582 26988
rect 20162 26936 20168 26988
rect 20220 26936 20226 26988
rect 20349 26979 20407 26985
rect 20349 26976 20361 26979
rect 20272 26948 20361 26976
rect 17972 26880 18460 26908
rect 19168 26908 19196 26936
rect 19334 26908 19340 26920
rect 19168 26880 19340 26908
rect 11330 26800 11336 26852
rect 11388 26840 11394 26852
rect 12434 26840 12440 26852
rect 11388 26812 12440 26840
rect 11388 26800 11394 26812
rect 12434 26800 12440 26812
rect 12492 26800 12498 26852
rect 18432 26840 18460 26880
rect 19334 26868 19340 26880
rect 19392 26868 19398 26920
rect 18432 26812 20024 26840
rect 11974 26772 11980 26784
rect 11072 26744 11980 26772
rect 10781 26735 10839 26741
rect 11974 26732 11980 26744
rect 12032 26732 12038 26784
rect 12250 26732 12256 26784
rect 12308 26772 12314 26784
rect 12345 26775 12403 26781
rect 12345 26772 12357 26775
rect 12308 26744 12357 26772
rect 12308 26732 12314 26744
rect 12345 26741 12357 26744
rect 12391 26741 12403 26775
rect 12345 26735 12403 26741
rect 12989 26775 13047 26781
rect 12989 26741 13001 26775
rect 13035 26772 13047 26775
rect 13078 26772 13084 26784
rect 13035 26744 13084 26772
rect 13035 26741 13047 26744
rect 12989 26735 13047 26741
rect 13078 26732 13084 26744
rect 13136 26732 13142 26784
rect 19426 26732 19432 26784
rect 19484 26772 19490 26784
rect 19794 26772 19800 26784
rect 19484 26744 19800 26772
rect 19484 26732 19490 26744
rect 19794 26732 19800 26744
rect 19852 26772 19858 26784
rect 19889 26775 19947 26781
rect 19889 26772 19901 26775
rect 19852 26744 19901 26772
rect 19852 26732 19858 26744
rect 19889 26741 19901 26744
rect 19935 26741 19947 26775
rect 19996 26772 20024 26812
rect 20070 26800 20076 26852
rect 20128 26800 20134 26852
rect 20272 26772 20300 26948
rect 20349 26945 20361 26948
rect 20395 26945 20407 26979
rect 20349 26939 20407 26945
rect 20438 26936 20444 26988
rect 20496 26976 20502 26988
rect 20732 26985 20760 27016
rect 21177 27013 21189 27047
rect 21223 27044 21235 27047
rect 22204 27044 22232 27075
rect 23290 27072 23296 27084
rect 23348 27072 23354 27124
rect 24854 27072 24860 27124
rect 24912 27072 24918 27124
rect 25041 27115 25099 27121
rect 25041 27081 25053 27115
rect 25087 27112 25099 27115
rect 25590 27112 25596 27124
rect 25087 27084 25596 27112
rect 25087 27081 25099 27084
rect 25041 27075 25099 27081
rect 25590 27072 25596 27084
rect 25648 27072 25654 27124
rect 25777 27115 25835 27121
rect 25777 27081 25789 27115
rect 25823 27112 25835 27115
rect 25866 27112 25872 27124
rect 25823 27084 25872 27112
rect 25823 27081 25835 27084
rect 25777 27075 25835 27081
rect 25866 27072 25872 27084
rect 25924 27072 25930 27124
rect 26050 27072 26056 27124
rect 26108 27072 26114 27124
rect 26234 27112 26240 27124
rect 26160 27084 26240 27112
rect 21223 27016 22232 27044
rect 22741 27047 22799 27053
rect 21223 27013 21235 27016
rect 21177 27007 21235 27013
rect 22741 27013 22753 27047
rect 22787 27044 22799 27047
rect 22830 27044 22836 27056
rect 22787 27016 22836 27044
rect 22787 27013 22799 27016
rect 22741 27007 22799 27013
rect 22830 27004 22836 27016
rect 22888 27004 22894 27056
rect 22925 27047 22983 27053
rect 22925 27013 22937 27047
rect 22971 27044 22983 27047
rect 23014 27044 23020 27056
rect 22971 27016 23020 27044
rect 22971 27013 22983 27016
rect 22925 27007 22983 27013
rect 23014 27004 23020 27016
rect 23072 27004 23078 27056
rect 23106 27004 23112 27056
rect 23164 27053 23170 27056
rect 23164 27047 23199 27053
rect 23187 27044 23199 27047
rect 23385 27047 23443 27053
rect 23385 27044 23397 27047
rect 23187 27016 23397 27044
rect 23187 27013 23199 27016
rect 23164 27007 23199 27013
rect 23385 27013 23397 27016
rect 23431 27013 23443 27047
rect 23385 27007 23443 27013
rect 23569 27047 23627 27053
rect 23569 27013 23581 27047
rect 23615 27044 23627 27047
rect 24486 27044 24492 27056
rect 23615 27016 24492 27044
rect 23615 27013 23627 27016
rect 23569 27007 23627 27013
rect 23164 27004 23170 27007
rect 24486 27004 24492 27016
rect 24544 27044 24550 27056
rect 26160 27044 26188 27084
rect 26234 27072 26240 27084
rect 26292 27072 26298 27124
rect 26326 27072 26332 27124
rect 26384 27072 26390 27124
rect 24544 27016 24900 27044
rect 24544 27004 24550 27016
rect 20533 26979 20591 26985
rect 20533 26976 20545 26979
rect 20496 26948 20545 26976
rect 20496 26936 20502 26948
rect 20533 26945 20545 26948
rect 20579 26945 20591 26979
rect 20533 26939 20591 26945
rect 20717 26979 20775 26985
rect 20717 26945 20729 26979
rect 20763 26945 20775 26979
rect 20717 26939 20775 26945
rect 20548 26908 20576 26939
rect 20990 26936 20996 26988
rect 21048 26976 21054 26988
rect 21544 26979 21602 26985
rect 21544 26976 21556 26979
rect 21048 26948 21556 26976
rect 21048 26936 21054 26948
rect 21544 26945 21556 26948
rect 21590 26945 21602 26979
rect 21544 26939 21602 26945
rect 21269 26911 21327 26917
rect 21269 26908 21281 26911
rect 20548 26880 21281 26908
rect 21269 26877 21281 26880
rect 21315 26877 21327 26911
rect 21559 26908 21587 26939
rect 21634 26936 21640 26988
rect 21692 26976 21698 26988
rect 22186 26976 22192 26988
rect 21692 26948 22192 26976
rect 21692 26936 21698 26948
rect 22186 26936 22192 26948
rect 22244 26936 22250 26988
rect 21559 26880 22232 26908
rect 21269 26871 21327 26877
rect 20346 26800 20352 26852
rect 20404 26840 20410 26852
rect 20809 26843 20867 26849
rect 20809 26840 20821 26843
rect 20404 26812 20821 26840
rect 20404 26800 20410 26812
rect 20809 26809 20821 26812
rect 20855 26809 20867 26843
rect 20809 26803 20867 26809
rect 20901 26843 20959 26849
rect 20901 26809 20913 26843
rect 20947 26840 20959 26843
rect 20990 26840 20996 26852
rect 20947 26812 20996 26840
rect 20947 26809 20959 26812
rect 20901 26803 20959 26809
rect 20990 26800 20996 26812
rect 21048 26800 21054 26852
rect 22204 26840 22232 26880
rect 22278 26868 22284 26920
rect 22336 26868 22342 26920
rect 23032 26908 23060 27004
rect 24210 26936 24216 26988
rect 24268 26936 24274 26988
rect 24394 26936 24400 26988
rect 24452 26976 24458 26988
rect 24670 26976 24676 26988
rect 24452 26948 24676 26976
rect 24452 26936 24458 26948
rect 24670 26936 24676 26948
rect 24728 26936 24734 26988
rect 24412 26908 24440 26936
rect 22756 26880 24440 26908
rect 22646 26840 22652 26852
rect 22020 26812 22140 26840
rect 22204 26812 22652 26840
rect 22020 26772 22048 26812
rect 19996 26744 22048 26772
rect 22112 26772 22140 26812
rect 22646 26800 22652 26812
rect 22704 26800 22710 26852
rect 22756 26849 22784 26880
rect 24486 26868 24492 26920
rect 24544 26868 24550 26920
rect 24872 26908 24900 27016
rect 24964 27016 26188 27044
rect 24964 26988 24992 27016
rect 24946 26936 24952 26988
rect 25004 26936 25010 26988
rect 25133 26979 25191 26985
rect 25133 26945 25145 26979
rect 25179 26976 25191 26979
rect 25314 26976 25320 26988
rect 25179 26948 25320 26976
rect 25179 26945 25191 26948
rect 25133 26939 25191 26945
rect 25314 26936 25320 26948
rect 25372 26976 25378 26988
rect 25685 26979 25743 26985
rect 25685 26976 25697 26979
rect 25372 26948 25697 26976
rect 25372 26936 25378 26948
rect 25685 26945 25697 26948
rect 25731 26945 25743 26979
rect 25685 26939 25743 26945
rect 25774 26936 25780 26988
rect 25832 26976 25838 26988
rect 25869 26979 25927 26985
rect 25869 26976 25881 26979
rect 25832 26948 25881 26976
rect 25832 26936 25838 26948
rect 25869 26945 25881 26948
rect 25915 26945 25927 26979
rect 25869 26939 25927 26945
rect 25498 26908 25504 26920
rect 24872 26880 25504 26908
rect 25498 26868 25504 26880
rect 25556 26868 25562 26920
rect 22741 26843 22799 26849
rect 22741 26809 22753 26843
rect 22787 26809 22799 26843
rect 24026 26840 24032 26852
rect 22741 26803 22799 26809
rect 23032 26812 24032 26840
rect 23032 26772 23060 26812
rect 24026 26800 24032 26812
rect 24084 26840 24090 26852
rect 25884 26840 25912 26939
rect 25958 26936 25964 26988
rect 26016 26936 26022 26988
rect 26160 26985 26188 27016
rect 26145 26979 26203 26985
rect 26145 26945 26157 26979
rect 26191 26945 26203 26979
rect 26145 26939 26203 26945
rect 26237 26979 26295 26985
rect 26237 26945 26249 26979
rect 26283 26945 26295 26979
rect 26237 26939 26295 26945
rect 26421 26979 26479 26985
rect 26421 26945 26433 26979
rect 26467 26945 26479 26979
rect 26421 26939 26479 26945
rect 25976 26908 26004 26936
rect 26252 26908 26280 26939
rect 25976 26880 26280 26908
rect 26436 26840 26464 26939
rect 26510 26936 26516 26988
rect 26568 26976 26574 26988
rect 27525 26979 27583 26985
rect 27525 26976 27537 26979
rect 26568 26948 27537 26976
rect 26568 26936 26574 26948
rect 27525 26945 27537 26948
rect 27571 26945 27583 26979
rect 27525 26939 27583 26945
rect 26786 26840 26792 26852
rect 24084 26812 26792 26840
rect 24084 26800 24090 26812
rect 26786 26800 26792 26812
rect 26844 26800 26850 26852
rect 22112 26744 23060 26772
rect 19889 26735 19947 26741
rect 23106 26732 23112 26784
rect 23164 26732 23170 26784
rect 23293 26775 23351 26781
rect 23293 26741 23305 26775
rect 23339 26772 23351 26775
rect 23382 26772 23388 26784
rect 23339 26744 23388 26772
rect 23339 26741 23351 26744
rect 23293 26735 23351 26741
rect 23382 26732 23388 26744
rect 23440 26732 23446 26784
rect 24302 26732 24308 26784
rect 24360 26772 24366 26784
rect 24578 26772 24584 26784
rect 24360 26744 24584 26772
rect 24360 26732 24366 26744
rect 24578 26732 24584 26744
rect 24636 26732 24642 26784
rect 24670 26732 24676 26784
rect 24728 26772 24734 26784
rect 27062 26772 27068 26784
rect 24728 26744 27068 26772
rect 24728 26732 24734 26744
rect 27062 26732 27068 26744
rect 27120 26732 27126 26784
rect 27706 26732 27712 26784
rect 27764 26732 27770 26784
rect 1104 26682 28152 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 28152 26682
rect 1104 26608 28152 26630
rect 2314 26528 2320 26580
rect 2372 26568 2378 26580
rect 2372 26540 3096 26568
rect 2372 26528 2378 26540
rect 3068 26500 3096 26540
rect 3142 26528 3148 26580
rect 3200 26568 3206 26580
rect 3237 26571 3295 26577
rect 3237 26568 3249 26571
rect 3200 26540 3249 26568
rect 3200 26528 3206 26540
rect 3237 26537 3249 26540
rect 3283 26568 3295 26571
rect 3694 26568 3700 26580
rect 3283 26540 3700 26568
rect 3283 26537 3295 26540
rect 3237 26531 3295 26537
rect 3694 26528 3700 26540
rect 3752 26528 3758 26580
rect 3970 26528 3976 26580
rect 4028 26528 4034 26580
rect 4249 26571 4307 26577
rect 4249 26537 4261 26571
rect 4295 26568 4307 26571
rect 4798 26568 4804 26580
rect 4295 26540 4804 26568
rect 4295 26537 4307 26540
rect 4249 26531 4307 26537
rect 4798 26528 4804 26540
rect 4856 26528 4862 26580
rect 5166 26528 5172 26580
rect 5224 26568 5230 26580
rect 6178 26568 6184 26580
rect 5224 26540 6184 26568
rect 5224 26528 5230 26540
rect 6178 26528 6184 26540
rect 6236 26568 6242 26580
rect 6914 26568 6920 26580
rect 6236 26540 6920 26568
rect 6236 26528 6242 26540
rect 6914 26528 6920 26540
rect 6972 26528 6978 26580
rect 9493 26571 9551 26577
rect 9493 26537 9505 26571
rect 9539 26568 9551 26571
rect 9858 26568 9864 26580
rect 9539 26540 9864 26568
rect 9539 26537 9551 26540
rect 9493 26531 9551 26537
rect 9858 26528 9864 26540
rect 9916 26528 9922 26580
rect 12069 26571 12127 26577
rect 12069 26537 12081 26571
rect 12115 26568 12127 26571
rect 12526 26568 12532 26580
rect 12115 26540 12532 26568
rect 12115 26537 12127 26540
rect 12069 26531 12127 26537
rect 12526 26528 12532 26540
rect 12584 26528 12590 26580
rect 17954 26528 17960 26580
rect 18012 26568 18018 26580
rect 19705 26571 19763 26577
rect 19705 26568 19717 26571
rect 18012 26540 19717 26568
rect 18012 26528 18018 26540
rect 19705 26537 19717 26540
rect 19751 26537 19763 26571
rect 19705 26531 19763 26537
rect 20162 26528 20168 26580
rect 20220 26528 20226 26580
rect 20346 26528 20352 26580
rect 20404 26528 20410 26580
rect 20990 26528 20996 26580
rect 21048 26568 21054 26580
rect 22370 26568 22376 26580
rect 21048 26540 22376 26568
rect 21048 26528 21054 26540
rect 22370 26528 22376 26540
rect 22428 26528 22434 26580
rect 22922 26528 22928 26580
rect 22980 26568 22986 26580
rect 24670 26568 24676 26580
rect 22980 26540 24676 26568
rect 22980 26528 22986 26540
rect 24670 26528 24676 26540
rect 24728 26528 24734 26580
rect 26786 26528 26792 26580
rect 26844 26528 26850 26580
rect 4706 26500 4712 26512
rect 1964 26472 2774 26500
rect 3068 26472 4712 26500
rect 1964 26382 1992 26472
rect 2746 26432 2774 26472
rect 4706 26460 4712 26472
rect 4764 26500 4770 26512
rect 5537 26503 5595 26509
rect 4764 26472 5396 26500
rect 4764 26460 4770 26472
rect 5074 26432 5080 26444
rect 2746 26404 5080 26432
rect 1952 26376 2004 26382
rect 1854 26324 1860 26376
rect 1912 26324 1918 26376
rect 3050 26324 3056 26376
rect 3108 26364 3114 26376
rect 3329 26367 3387 26373
rect 3329 26364 3341 26367
rect 3108 26336 3341 26364
rect 3108 26324 3114 26336
rect 3329 26333 3341 26336
rect 3375 26333 3387 26367
rect 3329 26327 3387 26333
rect 3878 26324 3884 26376
rect 3936 26364 3942 26376
rect 5000 26373 5028 26404
rect 5074 26392 5080 26404
rect 5132 26432 5138 26444
rect 5132 26404 5304 26432
rect 5132 26392 5138 26404
rect 4249 26367 4307 26373
rect 4249 26364 4261 26367
rect 3936 26336 4261 26364
rect 3936 26324 3942 26336
rect 4249 26333 4261 26336
rect 4295 26333 4307 26367
rect 4249 26327 4307 26333
rect 4433 26367 4491 26373
rect 4433 26333 4445 26367
rect 4479 26333 4491 26367
rect 4433 26327 4491 26333
rect 4985 26367 5043 26373
rect 4985 26333 4997 26367
rect 5031 26333 5043 26367
rect 4985 26327 5043 26333
rect 1952 26318 2004 26324
rect 2774 26256 2780 26308
rect 2832 26296 2838 26308
rect 2869 26299 2927 26305
rect 2869 26296 2881 26299
rect 2832 26268 2881 26296
rect 2832 26256 2838 26268
rect 2869 26265 2881 26268
rect 2915 26265 2927 26299
rect 2869 26259 2927 26265
rect 3418 26256 3424 26308
rect 3476 26296 3482 26308
rect 4448 26296 4476 26327
rect 5166 26324 5172 26376
rect 5224 26324 5230 26376
rect 5276 26373 5304 26404
rect 5368 26373 5396 26472
rect 5537 26469 5549 26503
rect 5583 26469 5595 26503
rect 5537 26463 5595 26469
rect 5552 26432 5580 26463
rect 12618 26460 12624 26512
rect 12676 26500 12682 26512
rect 12805 26503 12863 26509
rect 12805 26500 12817 26503
rect 12676 26472 12817 26500
rect 12676 26460 12682 26472
rect 12805 26469 12817 26472
rect 12851 26469 12863 26503
rect 12805 26463 12863 26469
rect 22833 26503 22891 26509
rect 22833 26469 22845 26503
rect 22879 26500 22891 26503
rect 23014 26500 23020 26512
rect 22879 26472 23020 26500
rect 22879 26469 22891 26472
rect 22833 26463 22891 26469
rect 23014 26460 23020 26472
rect 23072 26500 23078 26512
rect 23072 26472 23244 26500
rect 23072 26460 23078 26472
rect 5552 26404 5948 26432
rect 5261 26367 5319 26373
rect 5261 26333 5273 26367
rect 5307 26333 5319 26367
rect 5261 26327 5319 26333
rect 5353 26367 5411 26373
rect 5353 26333 5365 26367
rect 5399 26333 5411 26367
rect 5353 26327 5411 26333
rect 5534 26324 5540 26376
rect 5592 26324 5598 26376
rect 5810 26324 5816 26376
rect 5868 26324 5874 26376
rect 5920 26373 5948 26404
rect 6454 26392 6460 26444
rect 6512 26392 6518 26444
rect 6546 26392 6552 26444
rect 6604 26432 6610 26444
rect 11238 26432 11244 26444
rect 6604 26404 6868 26432
rect 6604 26392 6610 26404
rect 5905 26367 5963 26373
rect 5905 26333 5917 26367
rect 5951 26333 5963 26367
rect 6365 26367 6423 26373
rect 6365 26364 6377 26367
rect 5905 26327 5963 26333
rect 6196 26336 6377 26364
rect 4614 26296 4620 26308
rect 3476 26268 4384 26296
rect 4448 26268 4620 26296
rect 3476 26256 3482 26268
rect 4356 26228 4384 26268
rect 4614 26256 4620 26268
rect 4672 26296 4678 26308
rect 5077 26299 5135 26305
rect 5077 26296 5089 26299
rect 4672 26268 5089 26296
rect 4672 26256 4678 26268
rect 5077 26265 5089 26268
rect 5123 26265 5135 26299
rect 5077 26259 5135 26265
rect 6086 26256 6092 26308
rect 6144 26256 6150 26308
rect 6196 26228 6224 26336
rect 6365 26333 6377 26336
rect 6411 26364 6423 26367
rect 6730 26364 6736 26376
rect 6411 26336 6736 26364
rect 6411 26333 6423 26336
rect 6365 26327 6423 26333
rect 6730 26324 6736 26336
rect 6788 26324 6794 26376
rect 6840 26373 6868 26404
rect 9324 26404 9904 26432
rect 9324 26376 9352 26404
rect 6825 26367 6883 26373
rect 6825 26333 6837 26367
rect 6871 26333 6883 26367
rect 6825 26327 6883 26333
rect 9033 26367 9091 26373
rect 9033 26333 9045 26367
rect 9079 26333 9091 26367
rect 9033 26327 9091 26333
rect 4356 26200 6224 26228
rect 6733 26231 6791 26237
rect 6733 26197 6745 26231
rect 6779 26228 6791 26231
rect 6822 26228 6828 26240
rect 6779 26200 6828 26228
rect 6779 26197 6791 26200
rect 6733 26191 6791 26197
rect 6822 26188 6828 26200
rect 6880 26188 6886 26240
rect 8846 26188 8852 26240
rect 8904 26228 8910 26240
rect 9048 26228 9076 26327
rect 9122 26324 9128 26376
rect 9180 26324 9186 26376
rect 9306 26324 9312 26376
rect 9364 26324 9370 26376
rect 9876 26373 9904 26404
rect 10796 26404 11244 26432
rect 9585 26367 9643 26373
rect 9585 26333 9597 26367
rect 9631 26333 9643 26367
rect 9585 26327 9643 26333
rect 9677 26367 9735 26373
rect 9677 26333 9689 26367
rect 9723 26333 9735 26367
rect 9677 26327 9735 26333
rect 9861 26367 9919 26373
rect 9861 26333 9873 26367
rect 9907 26333 9919 26367
rect 9861 26327 9919 26333
rect 9140 26296 9168 26324
rect 9600 26296 9628 26327
rect 9140 26268 9628 26296
rect 9692 26228 9720 26327
rect 10594 26324 10600 26376
rect 10652 26324 10658 26376
rect 10796 26373 10824 26404
rect 11238 26392 11244 26404
rect 11296 26392 11302 26444
rect 12713 26435 12771 26441
rect 12713 26401 12725 26435
rect 12759 26432 12771 26435
rect 19981 26435 20039 26441
rect 12759 26404 13400 26432
rect 12759 26401 12771 26404
rect 12713 26395 12771 26401
rect 10781 26367 10839 26373
rect 10781 26333 10793 26367
rect 10827 26333 10839 26367
rect 10781 26327 10839 26333
rect 10873 26367 10931 26373
rect 10873 26333 10885 26367
rect 10919 26364 10931 26367
rect 11330 26364 11336 26376
rect 10919 26336 11336 26364
rect 10919 26333 10931 26336
rect 10873 26327 10931 26333
rect 11330 26324 11336 26336
rect 11388 26324 11394 26376
rect 11974 26324 11980 26376
rect 12032 26324 12038 26376
rect 12253 26367 12311 26373
rect 12253 26333 12265 26367
rect 12299 26364 12311 26367
rect 12299 26336 12434 26364
rect 12299 26333 12311 26336
rect 12253 26327 12311 26333
rect 11992 26296 12020 26324
rect 12406 26296 12434 26336
rect 12526 26324 12532 26376
rect 12584 26324 12590 26376
rect 12986 26364 12992 26376
rect 12636 26336 12992 26364
rect 12636 26296 12664 26336
rect 12986 26324 12992 26336
rect 13044 26324 13050 26376
rect 13078 26324 13084 26376
rect 13136 26324 13142 26376
rect 13170 26324 13176 26376
rect 13228 26324 13234 26376
rect 13372 26373 13400 26404
rect 19981 26401 19993 26435
rect 20027 26432 20039 26435
rect 20438 26432 20444 26444
rect 20027 26404 20444 26432
rect 20027 26401 20039 26404
rect 19981 26395 20039 26401
rect 20438 26392 20444 26404
rect 20496 26392 20502 26444
rect 20717 26435 20775 26441
rect 20717 26401 20729 26435
rect 20763 26432 20775 26435
rect 21634 26432 21640 26444
rect 20763 26404 21640 26432
rect 20763 26401 20775 26404
rect 20717 26395 20775 26401
rect 21634 26392 21640 26404
rect 21692 26392 21698 26444
rect 23216 26441 23244 26472
rect 23566 26460 23572 26512
rect 23624 26460 23630 26512
rect 27522 26460 27528 26512
rect 27580 26500 27586 26512
rect 27709 26503 27767 26509
rect 27709 26500 27721 26503
rect 27580 26472 27721 26500
rect 27580 26460 27586 26472
rect 27709 26469 27721 26472
rect 27755 26469 27767 26503
rect 27709 26463 27767 26469
rect 23201 26435 23259 26441
rect 23201 26401 23213 26435
rect 23247 26401 23259 26435
rect 23201 26395 23259 26401
rect 23290 26392 23296 26444
rect 23348 26392 23354 26444
rect 25038 26392 25044 26444
rect 25096 26432 25102 26444
rect 25250 26435 25308 26441
rect 25250 26432 25262 26435
rect 25096 26404 25262 26432
rect 25096 26392 25102 26404
rect 25250 26401 25262 26404
rect 25296 26432 25308 26435
rect 25406 26432 25412 26444
rect 25296 26404 25412 26432
rect 25296 26401 25308 26404
rect 25250 26395 25308 26401
rect 25406 26392 25412 26404
rect 25464 26392 25470 26444
rect 26053 26435 26111 26441
rect 26053 26401 26065 26435
rect 26099 26432 26111 26435
rect 26234 26432 26240 26444
rect 26099 26404 26240 26432
rect 26099 26401 26111 26404
rect 26053 26395 26111 26401
rect 26234 26392 26240 26404
rect 26292 26392 26298 26444
rect 13357 26367 13415 26373
rect 13357 26333 13369 26367
rect 13403 26333 13415 26367
rect 13357 26327 13415 26333
rect 19794 26324 19800 26376
rect 19852 26364 19858 26376
rect 20257 26367 20315 26373
rect 20257 26364 20269 26367
rect 19852 26336 20269 26364
rect 19852 26324 19858 26336
rect 20257 26333 20269 26336
rect 20303 26364 20315 26367
rect 20533 26367 20591 26373
rect 20533 26364 20545 26367
rect 20303 26336 20545 26364
rect 20303 26333 20315 26336
rect 20257 26327 20315 26333
rect 20533 26333 20545 26336
rect 20579 26333 20591 26367
rect 20533 26327 20591 26333
rect 11992 26268 12296 26296
rect 12406 26268 12664 26296
rect 8904 26200 9720 26228
rect 8904 26188 8910 26200
rect 9766 26188 9772 26240
rect 9824 26188 9830 26240
rect 10870 26188 10876 26240
rect 10928 26188 10934 26240
rect 12268 26228 12296 26268
rect 12710 26256 12716 26308
rect 12768 26296 12774 26308
rect 12805 26299 12863 26305
rect 12805 26296 12817 26299
rect 12768 26268 12817 26296
rect 12768 26256 12774 26268
rect 12805 26265 12817 26268
rect 12851 26296 12863 26299
rect 13265 26299 13323 26305
rect 13265 26296 13277 26299
rect 12851 26268 13277 26296
rect 12851 26265 12863 26268
rect 12805 26259 12863 26265
rect 13265 26265 13277 26268
rect 13311 26265 13323 26299
rect 20548 26296 20576 26327
rect 22462 26324 22468 26376
rect 22520 26324 22526 26376
rect 22646 26324 22652 26376
rect 22704 26324 22710 26376
rect 22738 26324 22744 26376
rect 22796 26364 22802 26376
rect 22833 26367 22891 26373
rect 22833 26364 22845 26367
rect 22796 26336 22845 26364
rect 22796 26324 22802 26336
rect 22833 26333 22845 26336
rect 22879 26333 22891 26367
rect 22833 26327 22891 26333
rect 22922 26324 22928 26376
rect 22980 26324 22986 26376
rect 24302 26324 24308 26376
rect 24360 26364 24366 26376
rect 24765 26367 24823 26373
rect 24765 26364 24777 26367
rect 24360 26336 24777 26364
rect 24360 26324 24366 26336
rect 24765 26333 24777 26336
rect 24811 26333 24823 26367
rect 24765 26327 24823 26333
rect 25130 26324 25136 26376
rect 25188 26364 25194 26376
rect 25188 26336 25560 26364
rect 25188 26324 25194 26336
rect 22278 26296 22284 26308
rect 20548 26268 22284 26296
rect 13265 26259 13323 26265
rect 22278 26256 22284 26268
rect 22336 26296 22342 26308
rect 23106 26296 23112 26308
rect 22336 26268 23112 26296
rect 22336 26256 22342 26268
rect 23106 26256 23112 26268
rect 23164 26256 23170 26308
rect 23410 26299 23468 26305
rect 23410 26265 23422 26299
rect 23456 26296 23468 26299
rect 24394 26296 24400 26308
rect 23456 26268 24400 26296
rect 23456 26265 23468 26268
rect 23410 26259 23468 26265
rect 12345 26231 12403 26237
rect 12345 26228 12357 26231
rect 12268 26200 12357 26228
rect 12345 26197 12357 26200
rect 12391 26197 12403 26231
rect 12345 26191 12403 26197
rect 12434 26188 12440 26240
rect 12492 26228 12498 26240
rect 12989 26231 13047 26237
rect 12989 26228 13001 26231
rect 12492 26200 13001 26228
rect 12492 26188 12498 26200
rect 12989 26197 13001 26200
rect 13035 26197 13047 26231
rect 12989 26191 13047 26197
rect 20162 26188 20168 26240
rect 20220 26228 20226 26240
rect 20438 26228 20444 26240
rect 20220 26200 20444 26228
rect 20220 26188 20226 26200
rect 20438 26188 20444 26200
rect 20496 26228 20502 26240
rect 23425 26228 23453 26259
rect 24394 26256 24400 26268
rect 24452 26256 24458 26308
rect 24486 26256 24492 26308
rect 24544 26296 24550 26308
rect 25041 26299 25099 26305
rect 25041 26296 25053 26299
rect 24544 26268 25053 26296
rect 24544 26256 24550 26268
rect 25041 26265 25053 26268
rect 25087 26296 25099 26299
rect 25222 26296 25228 26308
rect 25087 26268 25228 26296
rect 25087 26265 25099 26268
rect 25041 26259 25099 26265
rect 25222 26256 25228 26268
rect 25280 26256 25286 26308
rect 25532 26296 25560 26336
rect 25590 26324 25596 26376
rect 25648 26364 25654 26376
rect 25685 26367 25743 26373
rect 25685 26364 25697 26367
rect 25648 26336 25697 26364
rect 25648 26324 25654 26336
rect 25685 26333 25697 26336
rect 25731 26333 25743 26367
rect 25685 26327 25743 26333
rect 26326 26324 26332 26376
rect 26384 26364 26390 26376
rect 26697 26367 26755 26373
rect 26697 26364 26709 26367
rect 26384 26336 26709 26364
rect 26384 26324 26390 26336
rect 26697 26333 26709 26336
rect 26743 26333 26755 26367
rect 26697 26327 26755 26333
rect 26786 26324 26792 26376
rect 26844 26364 26850 26376
rect 27525 26367 27583 26373
rect 27525 26364 27537 26367
rect 26844 26336 27537 26364
rect 26844 26324 26850 26336
rect 27525 26333 27537 26336
rect 27571 26333 27583 26367
rect 27525 26327 27583 26333
rect 25532 26268 25728 26296
rect 25700 26240 25728 26268
rect 26418 26256 26424 26308
rect 26476 26296 26482 26308
rect 26513 26299 26571 26305
rect 26513 26296 26525 26299
rect 26476 26268 26525 26296
rect 26476 26256 26482 26268
rect 26513 26265 26525 26268
rect 26559 26265 26571 26299
rect 26513 26259 26571 26265
rect 20496 26200 23453 26228
rect 20496 26188 20502 26200
rect 25406 26188 25412 26240
rect 25464 26188 25470 26240
rect 25682 26188 25688 26240
rect 25740 26188 25746 26240
rect 1104 26138 28152 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 28152 26138
rect 1104 26064 28152 26086
rect 7944 25996 8432 26024
rect 5442 25916 5448 25968
rect 5500 25956 5506 25968
rect 7944 25956 7972 25996
rect 5500 25928 7972 25956
rect 5500 25916 5506 25928
rect 2774 25848 2780 25900
rect 2832 25848 2838 25900
rect 3142 25848 3148 25900
rect 3200 25848 3206 25900
rect 5994 25848 6000 25900
rect 6052 25888 6058 25900
rect 7944 25897 7972 25928
rect 8202 25916 8208 25968
rect 8260 25916 8266 25968
rect 8404 25965 8432 25996
rect 12250 25984 12256 26036
rect 12308 25984 12314 26036
rect 12434 25984 12440 26036
rect 12492 25984 12498 26036
rect 12897 26027 12955 26033
rect 12897 25993 12909 26027
rect 12943 26024 12955 26027
rect 13170 26024 13176 26036
rect 12943 25996 13176 26024
rect 12943 25993 12955 25996
rect 12897 25987 12955 25993
rect 13170 25984 13176 25996
rect 13228 25984 13234 26036
rect 25406 25984 25412 26036
rect 25464 26024 25470 26036
rect 26161 26027 26219 26033
rect 26161 26024 26173 26027
rect 25464 25996 26173 26024
rect 25464 25984 25470 25996
rect 26161 25993 26173 25996
rect 26207 25993 26219 26027
rect 26161 25987 26219 25993
rect 26329 26027 26387 26033
rect 26329 25993 26341 26027
rect 26375 26024 26387 26027
rect 26510 26024 26516 26036
rect 26375 25996 26516 26024
rect 26375 25993 26387 25996
rect 26329 25987 26387 25993
rect 26510 25984 26516 25996
rect 26568 25984 26574 26036
rect 8389 25959 8447 25965
rect 8389 25925 8401 25959
rect 8435 25925 8447 25959
rect 8389 25919 8447 25925
rect 8573 25959 8631 25965
rect 8573 25925 8585 25959
rect 8619 25956 8631 25959
rect 12268 25956 12296 25984
rect 12621 25959 12679 25965
rect 12621 25956 12633 25959
rect 8619 25928 8892 25956
rect 12268 25928 12633 25956
rect 8619 25925 8631 25928
rect 8573 25919 8631 25925
rect 6733 25891 6791 25897
rect 6733 25888 6745 25891
rect 6052 25860 6745 25888
rect 6052 25848 6058 25860
rect 6733 25857 6745 25860
rect 6779 25857 6791 25891
rect 6733 25851 6791 25857
rect 7929 25891 7987 25897
rect 7929 25857 7941 25891
rect 7975 25857 7987 25891
rect 7929 25851 7987 25857
rect 8123 25891 8181 25897
rect 8123 25857 8135 25891
rect 8169 25888 8181 25891
rect 8220 25888 8248 25916
rect 8864 25900 8892 25928
rect 12621 25925 12633 25928
rect 12667 25925 12679 25959
rect 12621 25919 12679 25925
rect 12802 25916 12808 25968
rect 12860 25916 12866 25968
rect 22462 25916 22468 25968
rect 22520 25956 22526 25968
rect 23014 25956 23020 25968
rect 22520 25928 23020 25956
rect 22520 25916 22526 25928
rect 23014 25916 23020 25928
rect 23072 25916 23078 25968
rect 23382 25916 23388 25968
rect 23440 25956 23446 25968
rect 25130 25956 25136 25968
rect 23440 25928 25136 25956
rect 23440 25916 23446 25928
rect 25130 25916 25136 25928
rect 25188 25956 25194 25968
rect 25501 25959 25559 25965
rect 25501 25956 25513 25959
rect 25188 25928 25513 25956
rect 25188 25916 25194 25928
rect 25501 25925 25513 25928
rect 25547 25925 25559 25959
rect 25501 25919 25559 25925
rect 25590 25916 25596 25968
rect 25648 25916 25654 25968
rect 25961 25959 26019 25965
rect 25961 25925 25973 25959
rect 26007 25925 26019 25959
rect 25961 25919 26019 25925
rect 8169 25860 8248 25888
rect 8665 25891 8723 25897
rect 8169 25857 8181 25860
rect 8123 25851 8181 25857
rect 8665 25857 8677 25891
rect 8711 25857 8723 25891
rect 8665 25851 8723 25857
rect 2501 25823 2559 25829
rect 2501 25789 2513 25823
rect 2547 25820 2559 25823
rect 2866 25820 2872 25832
rect 2547 25792 2872 25820
rect 2547 25789 2559 25792
rect 2501 25783 2559 25789
rect 2866 25780 2872 25792
rect 2924 25780 2930 25832
rect 6748 25752 6776 25851
rect 6822 25780 6828 25832
rect 6880 25820 6886 25832
rect 7193 25823 7251 25829
rect 7193 25820 7205 25823
rect 6880 25792 7205 25820
rect 6880 25780 6886 25792
rect 7193 25789 7205 25792
rect 7239 25789 7251 25823
rect 7193 25783 7251 25789
rect 8021 25823 8079 25829
rect 8021 25789 8033 25823
rect 8067 25820 8079 25823
rect 8680 25820 8708 25851
rect 8846 25848 8852 25900
rect 8904 25848 8910 25900
rect 12253 25891 12311 25897
rect 12253 25857 12265 25891
rect 12299 25857 12311 25891
rect 12253 25851 12311 25857
rect 12529 25891 12587 25897
rect 12529 25857 12541 25891
rect 12575 25888 12587 25891
rect 12710 25888 12716 25900
rect 12575 25860 12716 25888
rect 12575 25857 12587 25860
rect 12529 25851 12587 25857
rect 8067 25792 8708 25820
rect 12268 25820 12296 25851
rect 12710 25848 12716 25860
rect 12768 25848 12774 25900
rect 12897 25891 12955 25897
rect 12897 25857 12909 25891
rect 12943 25857 12955 25891
rect 12897 25851 12955 25857
rect 12618 25820 12624 25832
rect 12268 25792 12624 25820
rect 8067 25789 8079 25792
rect 8021 25783 8079 25789
rect 12618 25780 12624 25792
rect 12676 25780 12682 25832
rect 12802 25780 12808 25832
rect 12860 25820 12866 25832
rect 12912 25820 12940 25851
rect 20438 25848 20444 25900
rect 20496 25848 20502 25900
rect 20898 25848 20904 25900
rect 20956 25888 20962 25900
rect 22002 25888 22008 25900
rect 20956 25860 22008 25888
rect 20956 25848 20962 25860
rect 22002 25848 22008 25860
rect 22060 25888 22066 25900
rect 22060 25848 22094 25888
rect 22646 25848 22652 25900
rect 22704 25848 22710 25900
rect 22833 25891 22891 25897
rect 22833 25857 22845 25891
rect 22879 25888 22891 25891
rect 24210 25888 24216 25900
rect 22879 25860 24216 25888
rect 22879 25857 22891 25860
rect 22833 25851 22891 25857
rect 12860 25792 12940 25820
rect 22066 25820 22094 25848
rect 22848 25820 22876 25851
rect 24210 25848 24216 25860
rect 24268 25888 24274 25900
rect 24854 25888 24860 25900
rect 24268 25860 24860 25888
rect 24268 25848 24274 25860
rect 24854 25848 24860 25860
rect 24912 25888 24918 25900
rect 25038 25888 25044 25900
rect 24912 25860 25044 25888
rect 24912 25848 24918 25860
rect 25038 25848 25044 25860
rect 25096 25888 25102 25900
rect 25409 25891 25467 25897
rect 25409 25888 25421 25891
rect 25096 25860 25421 25888
rect 25096 25848 25102 25860
rect 25409 25857 25421 25860
rect 25455 25857 25467 25891
rect 25976 25888 26004 25919
rect 26326 25888 26332 25900
rect 25976 25860 26332 25888
rect 25409 25851 25467 25857
rect 26326 25848 26332 25860
rect 26384 25848 26390 25900
rect 26418 25848 26424 25900
rect 26476 25848 26482 25900
rect 22066 25792 22876 25820
rect 25777 25823 25835 25829
rect 12860 25780 12866 25792
rect 25777 25789 25789 25823
rect 25823 25820 25835 25823
rect 26786 25820 26792 25832
rect 25823 25792 26792 25820
rect 25823 25789 25835 25792
rect 25777 25783 25835 25789
rect 26786 25780 26792 25792
rect 26844 25780 26850 25832
rect 7469 25755 7527 25761
rect 7469 25752 7481 25755
rect 6748 25724 7481 25752
rect 7469 25721 7481 25724
rect 7515 25721 7527 25755
rect 7469 25715 7527 25721
rect 25225 25755 25283 25761
rect 25225 25721 25237 25755
rect 25271 25752 25283 25755
rect 25498 25752 25504 25764
rect 25271 25724 25504 25752
rect 25271 25721 25283 25724
rect 25225 25715 25283 25721
rect 25498 25712 25504 25724
rect 25556 25712 25562 25764
rect 25590 25712 25596 25764
rect 25648 25752 25654 25764
rect 26513 25755 26571 25761
rect 26513 25752 26525 25755
rect 25648 25724 26525 25752
rect 25648 25712 25654 25724
rect 7009 25687 7067 25693
rect 7009 25653 7021 25687
rect 7055 25684 7067 25687
rect 7558 25684 7564 25696
rect 7055 25656 7564 25684
rect 7055 25653 7067 25656
rect 7009 25647 7067 25653
rect 7558 25644 7564 25656
rect 7616 25644 7622 25696
rect 7650 25644 7656 25696
rect 7708 25644 7714 25696
rect 8662 25644 8668 25696
rect 8720 25684 8726 25696
rect 8757 25687 8815 25693
rect 8757 25684 8769 25687
rect 8720 25656 8769 25684
rect 8720 25644 8726 25656
rect 8757 25653 8769 25656
rect 8803 25653 8815 25687
rect 8757 25647 8815 25653
rect 12066 25644 12072 25696
rect 12124 25644 12130 25696
rect 20530 25644 20536 25696
rect 20588 25644 20594 25696
rect 26160 25693 26188 25724
rect 26513 25721 26525 25724
rect 26559 25721 26571 25755
rect 26513 25715 26571 25721
rect 26145 25687 26203 25693
rect 26145 25653 26157 25687
rect 26191 25653 26203 25687
rect 26145 25647 26203 25653
rect 1104 25594 28152 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 28152 25594
rect 1104 25520 28152 25542
rect 12434 25440 12440 25492
rect 12492 25480 12498 25492
rect 12986 25480 12992 25492
rect 12492 25452 12992 25480
rect 12492 25440 12498 25452
rect 12986 25440 12992 25452
rect 13044 25440 13050 25492
rect 15933 25483 15991 25489
rect 15933 25449 15945 25483
rect 15979 25480 15991 25483
rect 16945 25483 17003 25489
rect 16945 25480 16957 25483
rect 15979 25452 16957 25480
rect 15979 25449 15991 25452
rect 15933 25443 15991 25449
rect 16945 25449 16957 25452
rect 16991 25480 17003 25483
rect 17402 25480 17408 25492
rect 16991 25452 17408 25480
rect 16991 25449 17003 25452
rect 16945 25443 17003 25449
rect 17402 25440 17408 25452
rect 17460 25440 17466 25492
rect 23014 25440 23020 25492
rect 23072 25480 23078 25492
rect 25685 25483 25743 25489
rect 25685 25480 25697 25483
rect 23072 25452 25697 25480
rect 23072 25440 23078 25452
rect 25685 25449 25697 25452
rect 25731 25480 25743 25483
rect 25866 25480 25872 25492
rect 25731 25452 25872 25480
rect 25731 25449 25743 25452
rect 25685 25443 25743 25449
rect 25866 25440 25872 25452
rect 25924 25440 25930 25492
rect 26326 25440 26332 25492
rect 26384 25480 26390 25492
rect 26513 25483 26571 25489
rect 26513 25480 26525 25483
rect 26384 25452 26525 25480
rect 26384 25440 26390 25452
rect 26513 25449 26525 25452
rect 26559 25449 26571 25483
rect 26513 25443 26571 25449
rect 20530 25372 20536 25424
rect 20588 25412 20594 25424
rect 26234 25412 26240 25424
rect 20588 25384 26240 25412
rect 20588 25372 20594 25384
rect 26234 25372 26240 25384
rect 26292 25372 26298 25424
rect 13170 25344 13176 25356
rect 12360 25316 13176 25344
rect 9677 25279 9735 25285
rect 9677 25245 9689 25279
rect 9723 25276 9735 25279
rect 9766 25276 9772 25288
rect 9723 25248 9772 25276
rect 9723 25245 9735 25248
rect 9677 25239 9735 25245
rect 9766 25236 9772 25248
rect 9824 25236 9830 25288
rect 9858 25236 9864 25288
rect 9916 25276 9922 25288
rect 10229 25279 10287 25285
rect 10229 25276 10241 25279
rect 9916 25248 10241 25276
rect 9916 25236 9922 25248
rect 10229 25245 10241 25248
rect 10275 25245 10287 25279
rect 10229 25239 10287 25245
rect 10383 25279 10441 25285
rect 10383 25245 10395 25279
rect 10429 25276 10441 25279
rect 10686 25276 10692 25288
rect 10429 25248 10692 25276
rect 10429 25245 10441 25248
rect 10383 25239 10441 25245
rect 10244 25208 10272 25239
rect 10686 25236 10692 25248
rect 10744 25236 10750 25288
rect 10870 25236 10876 25288
rect 10928 25236 10934 25288
rect 12360 25285 12388 25316
rect 13170 25304 13176 25316
rect 13228 25304 13234 25356
rect 12345 25279 12403 25285
rect 12345 25245 12357 25279
rect 12391 25245 12403 25279
rect 12345 25239 12403 25245
rect 12434 25236 12440 25288
rect 12492 25236 12498 25288
rect 12618 25236 12624 25288
rect 12676 25236 12682 25288
rect 12710 25236 12716 25288
rect 12768 25236 12774 25288
rect 15562 25236 15568 25288
rect 15620 25236 15626 25288
rect 15654 25236 15660 25288
rect 15712 25236 15718 25288
rect 15749 25279 15807 25285
rect 15749 25245 15761 25279
rect 15795 25276 15807 25279
rect 15930 25276 15936 25288
rect 15795 25248 15936 25276
rect 15795 25245 15807 25248
rect 15749 25239 15807 25245
rect 15930 25236 15936 25248
rect 15988 25236 15994 25288
rect 22002 25236 22008 25288
rect 22060 25236 22066 25288
rect 25314 25236 25320 25288
rect 25372 25276 25378 25288
rect 25593 25279 25651 25285
rect 25593 25276 25605 25279
rect 25372 25248 25605 25276
rect 25372 25236 25378 25248
rect 25593 25245 25605 25248
rect 25639 25245 25651 25279
rect 25593 25239 25651 25245
rect 25869 25279 25927 25285
rect 25869 25245 25881 25279
rect 25915 25245 25927 25279
rect 25869 25239 25927 25245
rect 11054 25208 11060 25220
rect 10244 25180 11060 25208
rect 11054 25168 11060 25180
rect 11112 25168 11118 25220
rect 12897 25211 12955 25217
rect 12897 25177 12909 25211
rect 12943 25177 12955 25211
rect 15580 25208 15608 25236
rect 16114 25208 16120 25220
rect 15580 25180 16120 25208
rect 12897 25171 12955 25177
rect 9858 25100 9864 25152
rect 9916 25100 9922 25152
rect 10597 25143 10655 25149
rect 10597 25109 10609 25143
rect 10643 25140 10655 25143
rect 10686 25140 10692 25152
rect 10643 25112 10692 25140
rect 10643 25109 10655 25112
rect 10597 25103 10655 25109
rect 10686 25100 10692 25112
rect 10744 25100 10750 25152
rect 10873 25143 10931 25149
rect 10873 25109 10885 25143
rect 10919 25140 10931 25143
rect 10962 25140 10968 25152
rect 10919 25112 10968 25140
rect 10919 25109 10931 25112
rect 10873 25103 10931 25109
rect 10962 25100 10968 25112
rect 11020 25100 11026 25152
rect 11882 25100 11888 25152
rect 11940 25140 11946 25152
rect 12161 25143 12219 25149
rect 12161 25140 12173 25143
rect 11940 25112 12173 25140
rect 11940 25100 11946 25112
rect 12161 25109 12173 25112
rect 12207 25109 12219 25143
rect 12161 25103 12219 25109
rect 12434 25100 12440 25152
rect 12492 25140 12498 25152
rect 12912 25140 12940 25171
rect 16114 25168 16120 25180
rect 16172 25168 16178 25220
rect 16761 25211 16819 25217
rect 16761 25177 16773 25211
rect 16807 25208 16819 25211
rect 17586 25208 17592 25220
rect 16807 25180 17592 25208
rect 16807 25177 16819 25180
rect 16761 25171 16819 25177
rect 17586 25168 17592 25180
rect 17644 25168 17650 25220
rect 22186 25168 22192 25220
rect 22244 25168 22250 25220
rect 25884 25208 25912 25239
rect 27522 25236 27528 25288
rect 27580 25236 27586 25288
rect 25608 25180 25912 25208
rect 26053 25211 26111 25217
rect 25608 25152 25636 25180
rect 26053 25177 26065 25211
rect 26099 25208 26111 25211
rect 26145 25211 26203 25217
rect 26145 25208 26157 25211
rect 26099 25180 26157 25208
rect 26099 25177 26111 25180
rect 26053 25171 26111 25177
rect 26145 25177 26157 25180
rect 26191 25177 26203 25211
rect 26145 25171 26203 25177
rect 26326 25168 26332 25220
rect 26384 25168 26390 25220
rect 27157 25211 27215 25217
rect 27157 25177 27169 25211
rect 27203 25208 27215 25211
rect 27430 25208 27436 25220
rect 27203 25180 27436 25208
rect 27203 25177 27215 25180
rect 27157 25171 27215 25177
rect 27430 25168 27436 25180
rect 27488 25168 27494 25220
rect 12492 25112 12940 25140
rect 12492 25100 12498 25112
rect 16942 25100 16948 25152
rect 17000 25149 17006 25152
rect 17000 25143 17019 25149
rect 17007 25109 17019 25143
rect 17000 25103 17019 25109
rect 17000 25100 17006 25103
rect 17126 25100 17132 25152
rect 17184 25100 17190 25152
rect 25590 25100 25596 25152
rect 25648 25100 25654 25152
rect 27062 25100 27068 25152
rect 27120 25100 27126 25152
rect 27706 25100 27712 25152
rect 27764 25100 27770 25152
rect 1104 25050 28152 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 28152 25050
rect 1104 24976 28152 24998
rect 10870 24896 10876 24948
rect 10928 24896 10934 24948
rect 10962 24896 10968 24948
rect 11020 24896 11026 24948
rect 11054 24896 11060 24948
rect 11112 24936 11118 24948
rect 14921 24939 14979 24945
rect 14921 24936 14933 24939
rect 11112 24908 14933 24936
rect 11112 24896 11118 24908
rect 14921 24905 14933 24908
rect 14967 24905 14979 24939
rect 14921 24899 14979 24905
rect 2866 24828 2872 24880
rect 2924 24868 2930 24880
rect 4890 24868 4896 24880
rect 2924 24840 3280 24868
rect 2924 24828 2930 24840
rect 842 24760 848 24812
rect 900 24800 906 24812
rect 1397 24803 1455 24809
rect 1397 24800 1409 24803
rect 900 24772 1409 24800
rect 900 24760 906 24772
rect 1397 24769 1409 24772
rect 1443 24769 1455 24803
rect 1397 24763 1455 24769
rect 2498 24760 2504 24812
rect 2556 24760 2562 24812
rect 2682 24760 2688 24812
rect 2740 24760 2746 24812
rect 2976 24809 3004 24840
rect 2777 24803 2835 24809
rect 2777 24769 2789 24803
rect 2823 24800 2835 24803
rect 2961 24803 3019 24809
rect 2823 24772 2857 24800
rect 2823 24769 2835 24772
rect 2777 24763 2835 24769
rect 2961 24769 2973 24803
rect 3007 24769 3019 24803
rect 2961 24763 3019 24769
rect 3145 24803 3203 24809
rect 3145 24769 3157 24803
rect 3191 24769 3203 24803
rect 3252 24786 3280 24840
rect 4632 24840 4896 24868
rect 3145 24763 3203 24769
rect 2593 24735 2651 24741
rect 2593 24701 2605 24735
rect 2639 24732 2651 24735
rect 2792 24732 2820 24763
rect 3160 24732 3188 24763
rect 4062 24760 4068 24812
rect 4120 24800 4126 24812
rect 4632 24809 4660 24840
rect 4890 24828 4896 24840
rect 4948 24868 4954 24880
rect 4948 24840 5488 24868
rect 4948 24828 4954 24840
rect 5460 24812 5488 24840
rect 9858 24828 9864 24880
rect 9916 24868 9922 24880
rect 10137 24871 10195 24877
rect 10137 24868 10149 24871
rect 9916 24840 10149 24868
rect 9916 24828 9922 24840
rect 10137 24837 10149 24840
rect 10183 24837 10195 24871
rect 10888 24868 10916 24896
rect 10137 24831 10195 24837
rect 10612 24840 10916 24868
rect 10980 24868 11008 24896
rect 12066 24877 12072 24880
rect 11793 24871 11851 24877
rect 10980 24840 11192 24868
rect 4433 24803 4491 24809
rect 4433 24800 4445 24803
rect 4120 24772 4445 24800
rect 4120 24760 4126 24772
rect 4433 24769 4445 24772
rect 4479 24769 4491 24803
rect 4433 24763 4491 24769
rect 4617 24803 4675 24809
rect 4617 24769 4629 24803
rect 4663 24769 4675 24803
rect 4617 24763 4675 24769
rect 5074 24760 5080 24812
rect 5132 24760 5138 24812
rect 5258 24760 5264 24812
rect 5316 24760 5322 24812
rect 5350 24760 5356 24812
rect 5408 24760 5414 24812
rect 5442 24760 5448 24812
rect 5500 24760 5506 24812
rect 7650 24760 7656 24812
rect 7708 24800 7714 24812
rect 8205 24803 8263 24809
rect 8205 24800 8217 24803
rect 7708 24772 8217 24800
rect 7708 24760 7714 24772
rect 8205 24769 8217 24772
rect 8251 24769 8263 24803
rect 8205 24763 8263 24769
rect 2639 24704 3188 24732
rect 4157 24735 4215 24741
rect 2639 24701 2651 24704
rect 2593 24695 2651 24701
rect 4157 24701 4169 24735
rect 4203 24732 4215 24735
rect 4706 24732 4712 24744
rect 4203 24704 4712 24732
rect 4203 24701 4215 24704
rect 4157 24695 4215 24701
rect 4706 24692 4712 24704
rect 4764 24692 4770 24744
rect 8220 24732 8248 24763
rect 8386 24760 8392 24812
rect 8444 24760 8450 24812
rect 8662 24760 8668 24812
rect 8720 24800 8726 24812
rect 10612 24809 10640 24840
rect 9033 24803 9091 24809
rect 9033 24800 9045 24803
rect 8720 24772 9045 24800
rect 8720 24760 8726 24772
rect 9033 24769 9045 24772
rect 9079 24769 9091 24803
rect 9033 24763 9091 24769
rect 10321 24803 10379 24809
rect 10321 24769 10333 24803
rect 10367 24769 10379 24803
rect 10321 24763 10379 24769
rect 10597 24803 10655 24809
rect 10597 24769 10609 24803
rect 10643 24769 10655 24803
rect 10597 24763 10655 24769
rect 9125 24735 9183 24741
rect 9125 24732 9137 24735
rect 8220 24704 9137 24732
rect 9125 24701 9137 24704
rect 9171 24701 9183 24735
rect 9125 24695 9183 24701
rect 9217 24735 9275 24741
rect 9217 24701 9229 24735
rect 9263 24701 9275 24735
rect 10336 24732 10364 24763
rect 10686 24760 10692 24812
rect 10744 24800 10750 24812
rect 10781 24803 10839 24809
rect 10781 24800 10793 24803
rect 10744 24772 10793 24800
rect 10744 24760 10750 24772
rect 10781 24769 10793 24772
rect 10827 24769 10839 24803
rect 10781 24763 10839 24769
rect 10870 24760 10876 24812
rect 10928 24760 10934 24812
rect 10965 24803 11023 24809
rect 10965 24769 10977 24803
rect 11011 24800 11023 24803
rect 11011 24772 11100 24800
rect 11011 24769 11023 24772
rect 10965 24763 11023 24769
rect 10336 24704 11008 24732
rect 9217 24695 9275 24701
rect 5169 24667 5227 24673
rect 5169 24633 5181 24667
rect 5215 24664 5227 24667
rect 5902 24664 5908 24676
rect 5215 24636 5908 24664
rect 5215 24633 5227 24636
rect 5169 24627 5227 24633
rect 5902 24624 5908 24636
rect 5960 24624 5966 24676
rect 8386 24624 8392 24676
rect 8444 24664 8450 24676
rect 9232 24664 9260 24695
rect 10980 24676 11008 24704
rect 8444 24636 9260 24664
rect 8444 24624 8450 24636
rect 10962 24624 10968 24676
rect 11020 24624 11026 24676
rect 1581 24599 1639 24605
rect 1581 24565 1593 24599
rect 1627 24596 1639 24599
rect 2130 24596 2136 24608
rect 1627 24568 2136 24596
rect 1627 24565 1639 24568
rect 1581 24559 1639 24565
rect 2130 24556 2136 24568
rect 2188 24556 2194 24608
rect 2958 24556 2964 24608
rect 3016 24556 3022 24608
rect 4525 24599 4583 24605
rect 4525 24565 4537 24599
rect 4571 24596 4583 24599
rect 4614 24596 4620 24608
rect 4571 24568 4620 24596
rect 4571 24565 4583 24568
rect 4525 24559 4583 24565
rect 4614 24556 4620 24568
rect 4672 24556 4678 24608
rect 8849 24599 8907 24605
rect 8849 24565 8861 24599
rect 8895 24596 8907 24599
rect 9306 24596 9312 24608
rect 8895 24568 9312 24596
rect 8895 24565 8907 24568
rect 8849 24559 8907 24565
rect 9306 24556 9312 24568
rect 9364 24556 9370 24608
rect 9398 24556 9404 24608
rect 9456 24556 9462 24608
rect 10410 24556 10416 24608
rect 10468 24596 10474 24608
rect 10505 24599 10563 24605
rect 10505 24596 10517 24599
rect 10468 24568 10517 24596
rect 10468 24556 10474 24568
rect 10505 24565 10517 24568
rect 10551 24596 10563 24599
rect 11072 24596 11100 24772
rect 11164 24664 11192 24840
rect 11793 24837 11805 24871
rect 11839 24837 11851 24871
rect 11793 24831 11851 24837
rect 12009 24871 12072 24877
rect 12009 24837 12021 24871
rect 12055 24837 12072 24871
rect 12009 24831 12072 24837
rect 11808 24800 11836 24831
rect 12066 24828 12072 24831
rect 12124 24828 12130 24880
rect 14936 24868 14964 24899
rect 15654 24896 15660 24948
rect 15712 24936 15718 24948
rect 15712 24908 16436 24936
rect 15712 24896 15718 24908
rect 15930 24868 15936 24880
rect 14936 24840 15936 24868
rect 15930 24828 15936 24840
rect 15988 24868 15994 24880
rect 16408 24877 16436 24908
rect 16850 24896 16856 24948
rect 16908 24896 16914 24948
rect 17402 24896 17408 24948
rect 17460 24896 17466 24948
rect 21545 24939 21603 24945
rect 21545 24905 21557 24939
rect 21591 24936 21603 24939
rect 22002 24936 22008 24948
rect 21591 24908 22008 24936
rect 21591 24905 21603 24908
rect 21545 24899 21603 24905
rect 22002 24896 22008 24908
rect 22060 24896 22066 24948
rect 25869 24939 25927 24945
rect 25869 24905 25881 24939
rect 25915 24936 25927 24939
rect 26326 24936 26332 24948
rect 25915 24908 26332 24936
rect 25915 24905 25927 24908
rect 25869 24899 25927 24905
rect 26326 24896 26332 24908
rect 26384 24936 26390 24948
rect 27173 24939 27231 24945
rect 27173 24936 27185 24939
rect 26384 24908 27185 24936
rect 26384 24896 26390 24908
rect 27173 24905 27185 24908
rect 27219 24905 27231 24939
rect 27173 24899 27231 24905
rect 16209 24871 16267 24877
rect 16209 24868 16221 24871
rect 15988 24840 16221 24868
rect 15988 24828 15994 24840
rect 16209 24837 16221 24840
rect 16255 24837 16267 24871
rect 16209 24831 16267 24837
rect 16393 24871 16451 24877
rect 16393 24837 16405 24871
rect 16439 24837 16451 24871
rect 19150 24868 19156 24880
rect 16393 24831 16451 24837
rect 17144 24840 19156 24868
rect 11808 24772 12020 24800
rect 11992 24744 12020 24772
rect 14826 24760 14832 24812
rect 14884 24760 14890 24812
rect 15105 24803 15163 24809
rect 15105 24769 15117 24803
rect 15151 24800 15163 24803
rect 15381 24803 15439 24809
rect 15381 24800 15393 24803
rect 15151 24772 15393 24800
rect 15151 24769 15163 24772
rect 15105 24763 15163 24769
rect 15381 24769 15393 24772
rect 15427 24800 15439 24803
rect 15562 24800 15568 24812
rect 15427 24772 15568 24800
rect 15427 24769 15439 24772
rect 15381 24763 15439 24769
rect 11974 24692 11980 24744
rect 12032 24692 12038 24744
rect 12342 24692 12348 24744
rect 12400 24732 12406 24744
rect 12526 24732 12532 24744
rect 12400 24704 12532 24732
rect 12400 24692 12406 24704
rect 12526 24692 12532 24704
rect 12584 24692 12590 24744
rect 15120 24664 15148 24763
rect 15562 24760 15568 24772
rect 15620 24760 15626 24812
rect 15654 24760 15660 24812
rect 15712 24800 15718 24812
rect 15826 24803 15884 24809
rect 15826 24800 15838 24803
rect 15712 24772 15838 24800
rect 15712 24760 15718 24772
rect 15826 24769 15838 24772
rect 15872 24769 15884 24803
rect 15826 24763 15884 24769
rect 16114 24760 16120 24812
rect 16172 24760 16178 24812
rect 17144 24809 17172 24840
rect 19150 24828 19156 24840
rect 19208 24828 19214 24880
rect 22186 24828 22192 24880
rect 22244 24868 22250 24880
rect 23750 24868 23756 24880
rect 22244 24840 23756 24868
rect 22244 24828 22250 24840
rect 16669 24803 16727 24809
rect 16669 24769 16681 24803
rect 16715 24769 16727 24803
rect 16669 24763 16727 24769
rect 16761 24803 16819 24809
rect 16761 24769 16773 24803
rect 16807 24769 16819 24803
rect 16761 24763 16819 24769
rect 17129 24803 17187 24809
rect 17129 24769 17141 24803
rect 17175 24769 17187 24803
rect 17129 24763 17187 24769
rect 17313 24803 17371 24809
rect 17313 24769 17325 24803
rect 17359 24769 17371 24803
rect 17313 24763 17371 24769
rect 15749 24735 15807 24741
rect 15749 24701 15761 24735
rect 15795 24732 15807 24735
rect 15930 24732 15936 24744
rect 15795 24704 15936 24732
rect 15795 24701 15807 24704
rect 15749 24695 15807 24701
rect 15930 24692 15936 24704
rect 15988 24692 15994 24744
rect 16684 24732 16712 24763
rect 16040 24704 16712 24732
rect 11164 24636 15148 24664
rect 15289 24667 15347 24673
rect 15289 24633 15301 24667
rect 15335 24664 15347 24667
rect 16040 24664 16068 24704
rect 15335 24636 16068 24664
rect 15335 24633 15347 24636
rect 15289 24627 15347 24633
rect 15856 24608 15884 24636
rect 16114 24624 16120 24676
rect 16172 24664 16178 24676
rect 16301 24667 16359 24673
rect 16301 24664 16313 24667
rect 16172 24636 16313 24664
rect 16172 24624 16178 24636
rect 16301 24633 16313 24636
rect 16347 24664 16359 24667
rect 16776 24664 16804 24763
rect 16942 24692 16948 24744
rect 17000 24732 17006 24744
rect 17328 24732 17356 24763
rect 17586 24760 17592 24812
rect 17644 24760 17650 24812
rect 19886 24760 19892 24812
rect 19944 24800 19950 24812
rect 21453 24803 21511 24809
rect 21453 24800 21465 24803
rect 19944 24772 21465 24800
rect 19944 24760 19950 24772
rect 21453 24769 21465 24772
rect 21499 24769 21511 24803
rect 21453 24763 21511 24769
rect 22002 24760 22008 24812
rect 22060 24760 22066 24812
rect 22296 24809 22324 24840
rect 23750 24828 23756 24840
rect 23808 24828 23814 24880
rect 25792 24840 26004 24868
rect 25792 24812 25820 24840
rect 22281 24803 22339 24809
rect 22281 24769 22293 24803
rect 22327 24769 22339 24803
rect 22281 24763 22339 24769
rect 22557 24803 22615 24809
rect 22557 24769 22569 24803
rect 22603 24800 22615 24803
rect 22603 24772 22784 24800
rect 22603 24769 22615 24772
rect 22557 24763 22615 24769
rect 17000 24704 17356 24732
rect 17000 24692 17006 24704
rect 16347 24636 16804 24664
rect 16347 24633 16359 24636
rect 16301 24627 16359 24633
rect 10551 24568 11100 24596
rect 11241 24599 11299 24605
rect 10551 24565 10563 24568
rect 10505 24559 10563 24565
rect 11241 24565 11253 24599
rect 11287 24596 11299 24599
rect 11698 24596 11704 24608
rect 11287 24568 11704 24596
rect 11287 24565 11299 24568
rect 11241 24559 11299 24565
rect 11698 24556 11704 24568
rect 11756 24596 11762 24608
rect 11977 24599 12035 24605
rect 11977 24596 11989 24599
rect 11756 24568 11989 24596
rect 11756 24556 11762 24568
rect 11977 24565 11989 24568
rect 12023 24565 12035 24599
rect 11977 24559 12035 24565
rect 12161 24599 12219 24605
rect 12161 24565 12173 24599
rect 12207 24596 12219 24599
rect 12986 24596 12992 24608
rect 12207 24568 12992 24596
rect 12207 24565 12219 24568
rect 12161 24559 12219 24565
rect 12986 24556 12992 24568
rect 13044 24556 13050 24608
rect 15838 24556 15844 24608
rect 15896 24556 15902 24608
rect 16025 24599 16083 24605
rect 16025 24565 16037 24599
rect 16071 24596 16083 24599
rect 16960 24596 16988 24692
rect 18046 24664 18052 24676
rect 17052 24636 18052 24664
rect 17052 24605 17080 24636
rect 18046 24624 18052 24636
rect 18104 24624 18110 24676
rect 21450 24624 21456 24676
rect 21508 24664 21514 24676
rect 22756 24664 22784 24772
rect 22922 24760 22928 24812
rect 22980 24760 22986 24812
rect 23106 24760 23112 24812
rect 23164 24760 23170 24812
rect 23201 24803 23259 24809
rect 23201 24769 23213 24803
rect 23247 24769 23259 24803
rect 23201 24763 23259 24769
rect 22833 24735 22891 24741
rect 22833 24701 22845 24735
rect 22879 24732 22891 24735
rect 23124 24732 23152 24760
rect 22879 24704 23152 24732
rect 22879 24701 22891 24704
rect 22833 24695 22891 24701
rect 22925 24667 22983 24673
rect 22925 24664 22937 24667
rect 21508 24636 22692 24664
rect 22756 24636 22937 24664
rect 21508 24624 21514 24636
rect 16071 24568 16988 24596
rect 17037 24599 17095 24605
rect 16071 24565 16083 24568
rect 16025 24559 16083 24565
rect 17037 24565 17049 24599
rect 17083 24565 17095 24599
rect 17037 24559 17095 24565
rect 17129 24599 17187 24605
rect 17129 24565 17141 24599
rect 17175 24596 17187 24599
rect 17218 24596 17224 24608
rect 17175 24568 17224 24596
rect 17175 24565 17187 24568
rect 17129 24559 17187 24565
rect 17218 24556 17224 24568
rect 17276 24556 17282 24608
rect 17773 24599 17831 24605
rect 17773 24565 17785 24599
rect 17819 24596 17831 24599
rect 17862 24596 17868 24608
rect 17819 24568 17868 24596
rect 17819 24565 17831 24568
rect 17773 24559 17831 24565
rect 17862 24556 17868 24568
rect 17920 24556 17926 24608
rect 21358 24556 21364 24608
rect 21416 24596 21422 24608
rect 21821 24599 21879 24605
rect 21821 24596 21833 24599
rect 21416 24568 21833 24596
rect 21416 24556 21422 24568
rect 21821 24565 21833 24568
rect 21867 24565 21879 24599
rect 21821 24559 21879 24565
rect 22186 24556 22192 24608
rect 22244 24556 22250 24608
rect 22370 24556 22376 24608
rect 22428 24556 22434 24608
rect 22664 24596 22692 24636
rect 22925 24633 22937 24636
rect 22971 24633 22983 24667
rect 22925 24627 22983 24633
rect 22741 24599 22799 24605
rect 22741 24596 22753 24599
rect 22664 24568 22753 24596
rect 22741 24565 22753 24568
rect 22787 24596 22799 24599
rect 23216 24596 23244 24763
rect 25222 24760 25228 24812
rect 25280 24800 25286 24812
rect 25774 24800 25780 24812
rect 25280 24772 25780 24800
rect 25280 24760 25286 24772
rect 25774 24760 25780 24772
rect 25832 24760 25838 24812
rect 25866 24760 25872 24812
rect 25924 24760 25930 24812
rect 25976 24809 26004 24840
rect 26234 24828 26240 24880
rect 26292 24868 26298 24880
rect 26973 24871 27031 24877
rect 26973 24868 26985 24871
rect 26292 24840 26985 24868
rect 26292 24828 26298 24840
rect 26973 24837 26985 24840
rect 27019 24837 27031 24871
rect 26973 24831 27031 24837
rect 25961 24803 26019 24809
rect 25961 24769 25973 24803
rect 26007 24769 26019 24803
rect 25961 24763 26019 24769
rect 26421 24803 26479 24809
rect 26421 24769 26433 24803
rect 26467 24800 26479 24803
rect 27525 24803 27583 24809
rect 27525 24800 27537 24803
rect 26467 24772 27200 24800
rect 26467 24769 26479 24772
rect 26421 24763 26479 24769
rect 25038 24692 25044 24744
rect 25096 24732 25102 24744
rect 25590 24732 25596 24744
rect 25096 24704 25596 24732
rect 25096 24692 25102 24704
rect 25590 24692 25596 24704
rect 25648 24732 25654 24744
rect 26237 24735 26295 24741
rect 26237 24732 26249 24735
rect 25648 24704 26249 24732
rect 25648 24692 25654 24704
rect 26237 24701 26249 24704
rect 26283 24701 26295 24735
rect 26237 24695 26295 24701
rect 27172 24608 27200 24772
rect 27356 24772 27537 24800
rect 27356 24673 27384 24772
rect 27525 24769 27537 24772
rect 27571 24769 27583 24803
rect 27525 24763 27583 24769
rect 27341 24667 27399 24673
rect 27341 24633 27353 24667
rect 27387 24633 27399 24667
rect 27341 24627 27399 24633
rect 23474 24596 23480 24608
rect 22787 24568 23480 24596
rect 22787 24565 22799 24568
rect 22741 24559 22799 24565
rect 23474 24556 23480 24568
rect 23532 24556 23538 24608
rect 25866 24556 25872 24608
rect 25924 24596 25930 24608
rect 26053 24599 26111 24605
rect 26053 24596 26065 24599
rect 25924 24568 26065 24596
rect 25924 24556 25930 24568
rect 26053 24565 26065 24568
rect 26099 24565 26111 24599
rect 26053 24559 26111 24565
rect 26605 24599 26663 24605
rect 26605 24565 26617 24599
rect 26651 24596 26663 24599
rect 26878 24596 26884 24608
rect 26651 24568 26884 24596
rect 26651 24565 26663 24568
rect 26605 24559 26663 24565
rect 26878 24556 26884 24568
rect 26936 24556 26942 24608
rect 27154 24556 27160 24608
rect 27212 24556 27218 24608
rect 27706 24556 27712 24608
rect 27764 24556 27770 24608
rect 1104 24506 28152 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 28152 24506
rect 1104 24432 28152 24454
rect 2774 24392 2780 24404
rect 2746 24352 2780 24392
rect 2832 24392 2838 24404
rect 3418 24392 3424 24404
rect 2832 24364 3424 24392
rect 2832 24352 2838 24364
rect 3418 24352 3424 24364
rect 3476 24352 3482 24404
rect 7837 24395 7895 24401
rect 7837 24361 7849 24395
rect 7883 24392 7895 24395
rect 8386 24392 8392 24404
rect 7883 24364 8392 24392
rect 7883 24361 7895 24364
rect 7837 24355 7895 24361
rect 8386 24352 8392 24364
rect 8444 24352 8450 24404
rect 10229 24395 10287 24401
rect 10229 24361 10241 24395
rect 10275 24392 10287 24395
rect 14826 24392 14832 24404
rect 10275 24364 14832 24392
rect 10275 24361 10287 24364
rect 10229 24355 10287 24361
rect 14826 24352 14832 24364
rect 14884 24392 14890 24404
rect 15654 24392 15660 24404
rect 14884 24364 15660 24392
rect 14884 24352 14890 24364
rect 2746 24256 2774 24352
rect 4062 24324 4068 24336
rect 2424 24228 2774 24256
rect 2884 24296 4068 24324
rect 2424 24197 2452 24228
rect 2409 24191 2467 24197
rect 2409 24157 2421 24191
rect 2455 24157 2467 24191
rect 2409 24151 2467 24157
rect 2498 24148 2504 24200
rect 2556 24148 2562 24200
rect 2590 24148 2596 24200
rect 2648 24188 2654 24200
rect 2884 24188 2912 24296
rect 4062 24284 4068 24296
rect 4120 24324 4126 24336
rect 4709 24327 4767 24333
rect 4120 24296 4476 24324
rect 4120 24284 4126 24296
rect 2958 24216 2964 24268
rect 3016 24256 3022 24268
rect 4448 24265 4476 24296
rect 4709 24293 4721 24327
rect 4755 24324 4767 24327
rect 9585 24327 9643 24333
rect 4755 24296 5120 24324
rect 4755 24293 4767 24296
rect 4709 24287 4767 24293
rect 5092 24268 5120 24296
rect 9585 24293 9597 24327
rect 9631 24324 9643 24327
rect 10870 24324 10876 24336
rect 9631 24296 10876 24324
rect 9631 24293 9643 24296
rect 9585 24287 9643 24293
rect 4249 24259 4307 24265
rect 4249 24256 4261 24259
rect 3016 24228 4261 24256
rect 3016 24216 3022 24228
rect 4249 24225 4261 24228
rect 4295 24225 4307 24259
rect 4249 24219 4307 24225
rect 4433 24259 4491 24265
rect 4433 24225 4445 24259
rect 4479 24256 4491 24259
rect 4798 24256 4804 24268
rect 4479 24228 4804 24256
rect 4479 24225 4491 24228
rect 4433 24219 4491 24225
rect 4798 24216 4804 24228
rect 4856 24216 4862 24268
rect 5074 24216 5080 24268
rect 5132 24216 5138 24268
rect 10704 24265 10732 24296
rect 10870 24284 10876 24296
rect 10928 24284 10934 24336
rect 12621 24327 12679 24333
rect 12621 24293 12633 24327
rect 12667 24324 12679 24327
rect 12710 24324 12716 24336
rect 12667 24296 12716 24324
rect 12667 24293 12679 24296
rect 12621 24287 12679 24293
rect 12710 24284 12716 24296
rect 12768 24284 12774 24336
rect 12989 24327 13047 24333
rect 12989 24293 13001 24327
rect 13035 24324 13047 24327
rect 14182 24324 14188 24336
rect 13035 24296 14188 24324
rect 13035 24293 13047 24296
rect 12989 24287 13047 24293
rect 14182 24284 14188 24296
rect 14240 24284 14246 24336
rect 10597 24259 10655 24265
rect 10597 24256 10609 24259
rect 9876 24228 10609 24256
rect 9876 24200 9904 24228
rect 10597 24225 10609 24228
rect 10643 24225 10655 24259
rect 10597 24219 10655 24225
rect 10689 24259 10747 24265
rect 10689 24225 10701 24259
rect 10735 24225 10747 24259
rect 10689 24219 10747 24225
rect 11698 24216 11704 24268
rect 11756 24216 11762 24268
rect 2648 24160 2912 24188
rect 4341 24191 4399 24197
rect 2648 24148 2654 24160
rect 4341 24157 4353 24191
rect 4387 24157 4399 24191
rect 4341 24151 4399 24157
rect 4525 24191 4583 24197
rect 4525 24157 4537 24191
rect 4571 24188 4583 24191
rect 4706 24188 4712 24200
rect 4571 24160 4712 24188
rect 4571 24157 4583 24160
rect 4525 24151 4583 24157
rect 842 24080 848 24132
rect 900 24120 906 24132
rect 1489 24123 1547 24129
rect 1489 24120 1501 24123
rect 900 24092 1501 24120
rect 900 24080 906 24092
rect 1489 24089 1501 24092
rect 1535 24089 1547 24123
rect 1489 24083 1547 24089
rect 2130 24080 2136 24132
rect 2188 24120 2194 24132
rect 3513 24123 3571 24129
rect 3513 24120 3525 24123
rect 2188 24092 3525 24120
rect 2188 24080 2194 24092
rect 3513 24089 3525 24092
rect 3559 24089 3571 24123
rect 4356 24120 4384 24151
rect 4706 24148 4712 24160
rect 4764 24148 4770 24200
rect 5258 24148 5264 24200
rect 5316 24148 5322 24200
rect 7466 24148 7472 24200
rect 7524 24148 7530 24200
rect 7558 24148 7564 24200
rect 7616 24188 7622 24200
rect 7653 24191 7711 24197
rect 7653 24188 7665 24191
rect 7616 24160 7665 24188
rect 7616 24148 7622 24160
rect 7653 24157 7665 24160
rect 7699 24157 7711 24191
rect 7653 24151 7711 24157
rect 9398 24148 9404 24200
rect 9456 24188 9462 24200
rect 9677 24191 9735 24197
rect 9677 24188 9689 24191
rect 9456 24160 9689 24188
rect 9456 24148 9462 24160
rect 9677 24157 9689 24160
rect 9723 24157 9735 24191
rect 9677 24151 9735 24157
rect 9769 24191 9827 24197
rect 9769 24157 9781 24191
rect 9815 24188 9827 24191
rect 9858 24188 9864 24200
rect 9815 24160 9864 24188
rect 9815 24157 9827 24160
rect 9769 24151 9827 24157
rect 9858 24148 9864 24160
rect 9916 24148 9922 24200
rect 9950 24148 9956 24200
rect 10008 24148 10014 24200
rect 10045 24191 10103 24197
rect 10045 24157 10057 24191
rect 10091 24157 10103 24191
rect 10045 24151 10103 24157
rect 4430 24120 4436 24132
rect 4356 24092 4436 24120
rect 3513 24083 3571 24089
rect 1765 24055 1823 24061
rect 1765 24021 1777 24055
rect 1811 24052 1823 24055
rect 2222 24052 2228 24064
rect 1811 24024 2228 24052
rect 1811 24021 1823 24024
rect 1765 24015 1823 24021
rect 2222 24012 2228 24024
rect 2280 24012 2286 24064
rect 3053 24055 3111 24061
rect 3053 24021 3065 24055
rect 3099 24052 3111 24055
rect 3142 24052 3148 24064
rect 3099 24024 3148 24052
rect 3099 24021 3111 24024
rect 3053 24015 3111 24021
rect 3142 24012 3148 24024
rect 3200 24012 3206 24064
rect 3528 24052 3556 24083
rect 4430 24080 4436 24092
rect 4488 24120 4494 24132
rect 4890 24120 4896 24132
rect 4488 24092 4896 24120
rect 4488 24080 4494 24092
rect 4890 24080 4896 24092
rect 4948 24080 4954 24132
rect 5626 24080 5632 24132
rect 5684 24080 5690 24132
rect 9214 24080 9220 24132
rect 9272 24120 9278 24132
rect 10060 24120 10088 24151
rect 10134 24148 10140 24200
rect 10192 24188 10198 24200
rect 10321 24191 10379 24197
rect 10321 24188 10333 24191
rect 10192 24160 10333 24188
rect 10192 24148 10198 24160
rect 10321 24157 10333 24160
rect 10367 24157 10379 24191
rect 10321 24151 10379 24157
rect 10413 24191 10471 24197
rect 10413 24157 10425 24191
rect 10459 24188 10471 24191
rect 10870 24188 10876 24200
rect 10459 24160 10876 24188
rect 10459 24157 10471 24160
rect 10413 24151 10471 24157
rect 9272 24092 10088 24120
rect 10336 24120 10364 24151
rect 10870 24148 10876 24160
rect 10928 24148 10934 24200
rect 11974 24148 11980 24200
rect 12032 24148 12038 24200
rect 12066 24148 12072 24200
rect 12124 24188 12130 24200
rect 12529 24191 12587 24197
rect 12529 24188 12541 24191
rect 12124 24160 12541 24188
rect 12124 24148 12130 24160
rect 12529 24157 12541 24160
rect 12575 24157 12587 24191
rect 12728 24188 12756 24284
rect 15120 24265 15148 24364
rect 15654 24352 15660 24364
rect 15712 24352 15718 24404
rect 21453 24395 21511 24401
rect 21453 24361 21465 24395
rect 21499 24392 21511 24395
rect 22002 24392 22008 24404
rect 21499 24364 22008 24392
rect 21499 24361 21511 24364
rect 21453 24355 21511 24361
rect 22002 24352 22008 24364
rect 22060 24352 22066 24404
rect 23106 24352 23112 24404
rect 23164 24392 23170 24404
rect 23293 24395 23351 24401
rect 23293 24392 23305 24395
rect 23164 24364 23305 24392
rect 23164 24352 23170 24364
rect 23293 24361 23305 24364
rect 23339 24361 23351 24395
rect 23293 24355 23351 24361
rect 17034 24284 17040 24336
rect 17092 24324 17098 24336
rect 17405 24327 17463 24333
rect 17405 24324 17417 24327
rect 17092 24296 17417 24324
rect 17092 24284 17098 24296
rect 17405 24293 17417 24296
rect 17451 24324 17463 24327
rect 17586 24324 17592 24336
rect 17451 24296 17592 24324
rect 17451 24293 17463 24296
rect 17405 24287 17463 24293
rect 17586 24284 17592 24296
rect 17644 24284 17650 24336
rect 15105 24259 15163 24265
rect 15105 24225 15117 24259
rect 15151 24225 15163 24259
rect 15105 24219 15163 24225
rect 15473 24259 15531 24265
rect 15473 24225 15485 24259
rect 15519 24256 15531 24259
rect 18046 24256 18052 24268
rect 15519 24228 18052 24256
rect 15519 24225 15531 24228
rect 15473 24219 15531 24225
rect 18046 24216 18052 24228
rect 18104 24256 18110 24268
rect 18506 24256 18512 24268
rect 18104 24228 18512 24256
rect 18104 24216 18110 24228
rect 18506 24216 18512 24228
rect 18564 24216 18570 24268
rect 21085 24259 21143 24265
rect 21085 24225 21097 24259
rect 21131 24256 21143 24259
rect 21821 24259 21879 24265
rect 21131 24228 21588 24256
rect 21131 24225 21143 24228
rect 21085 24219 21143 24225
rect 21560 24200 21588 24228
rect 21821 24225 21833 24259
rect 21867 24256 21879 24259
rect 22370 24256 22376 24268
rect 21867 24228 22376 24256
rect 21867 24225 21879 24228
rect 21821 24219 21879 24225
rect 22370 24216 22376 24228
rect 22428 24216 22434 24268
rect 23308 24256 23336 24355
rect 23474 24352 23480 24404
rect 23532 24352 23538 24404
rect 25866 24352 25872 24404
rect 25924 24352 25930 24404
rect 26881 24395 26939 24401
rect 26881 24361 26893 24395
rect 26927 24392 26939 24395
rect 27522 24392 27528 24404
rect 26927 24364 27528 24392
rect 26927 24361 26939 24364
rect 26881 24355 26939 24361
rect 27522 24352 27528 24364
rect 27580 24352 27586 24404
rect 24670 24284 24676 24336
rect 24728 24324 24734 24336
rect 24728 24296 25268 24324
rect 24728 24284 24734 24296
rect 24765 24259 24823 24265
rect 24765 24256 24777 24259
rect 23308 24228 24777 24256
rect 24765 24225 24777 24228
rect 24811 24256 24823 24259
rect 25038 24256 25044 24268
rect 24811 24228 25044 24256
rect 24811 24225 24823 24228
rect 24765 24219 24823 24225
rect 25038 24216 25044 24228
rect 25096 24216 25102 24268
rect 12805 24191 12863 24197
rect 12805 24188 12817 24191
rect 12728 24160 12817 24188
rect 12529 24151 12587 24157
rect 12805 24157 12817 24160
rect 12851 24157 12863 24191
rect 12805 24151 12863 24157
rect 12986 24148 12992 24200
rect 13044 24148 13050 24200
rect 14277 24191 14335 24197
rect 14277 24157 14289 24191
rect 14323 24188 14335 24191
rect 14366 24188 14372 24200
rect 14323 24160 14372 24188
rect 14323 24157 14335 24160
rect 14277 24151 14335 24157
rect 14366 24148 14372 24160
rect 14424 24148 14430 24200
rect 15289 24191 15347 24197
rect 15289 24157 15301 24191
rect 15335 24157 15347 24191
rect 15289 24151 15347 24157
rect 10594 24120 10600 24132
rect 10336 24092 10600 24120
rect 9272 24080 9278 24092
rect 10594 24080 10600 24092
rect 10652 24080 10658 24132
rect 10781 24123 10839 24129
rect 10781 24089 10793 24123
rect 10827 24120 10839 24123
rect 15304 24120 15332 24151
rect 15654 24148 15660 24200
rect 15712 24148 15718 24200
rect 17957 24191 18015 24197
rect 17957 24157 17969 24191
rect 18003 24188 18015 24191
rect 18003 24160 19104 24188
rect 18003 24157 18015 24160
rect 17957 24151 18015 24157
rect 10827 24092 15332 24120
rect 10827 24089 10839 24092
rect 10781 24083 10839 24089
rect 15930 24080 15936 24132
rect 15988 24080 15994 24132
rect 16390 24080 16396 24132
rect 16448 24080 16454 24132
rect 19076 24064 19104 24160
rect 21266 24148 21272 24200
rect 21324 24148 21330 24200
rect 21450 24148 21456 24200
rect 21508 24148 21514 24200
rect 21542 24148 21548 24200
rect 21600 24148 21606 24200
rect 23661 24191 23719 24197
rect 23661 24188 23673 24191
rect 23124 24160 23673 24188
rect 20346 24080 20352 24132
rect 20404 24120 20410 24132
rect 20404 24092 20484 24120
rect 20404 24080 20410 24092
rect 12434 24052 12440 24064
rect 3528 24024 12440 24052
rect 12434 24012 12440 24024
rect 12492 24012 12498 24064
rect 13538 24012 13544 24064
rect 13596 24052 13602 24064
rect 14185 24055 14243 24061
rect 14185 24052 14197 24055
rect 13596 24024 14197 24052
rect 13596 24012 13602 24024
rect 14185 24021 14197 24024
rect 14231 24021 14243 24055
rect 14185 24015 14243 24021
rect 17494 24012 17500 24064
rect 17552 24052 17558 24064
rect 17589 24055 17647 24061
rect 17589 24052 17601 24055
rect 17552 24024 17601 24052
rect 17552 24012 17558 24024
rect 17589 24021 17601 24024
rect 17635 24021 17647 24055
rect 17589 24015 17647 24021
rect 19058 24012 19064 24064
rect 19116 24052 19122 24064
rect 19337 24055 19395 24061
rect 19337 24052 19349 24055
rect 19116 24024 19349 24052
rect 19116 24012 19122 24024
rect 19337 24021 19349 24024
rect 19383 24021 19395 24055
rect 20456 24052 20484 24092
rect 20530 24080 20536 24132
rect 20588 24120 20594 24132
rect 20809 24123 20867 24129
rect 20809 24120 20821 24123
rect 20588 24092 20821 24120
rect 20588 24080 20594 24092
rect 20809 24089 20821 24092
rect 20855 24089 20867 24123
rect 20809 24083 20867 24089
rect 22066 24092 22310 24120
rect 22066 24064 22094 24092
rect 22002 24052 22008 24064
rect 20456 24024 22008 24052
rect 19337 24015 19395 24021
rect 22002 24012 22008 24024
rect 22060 24024 22094 24064
rect 22060 24012 22066 24024
rect 22186 24012 22192 24064
rect 22244 24052 22250 24064
rect 23124 24052 23152 24160
rect 23661 24157 23673 24160
rect 23707 24157 23719 24191
rect 23661 24151 23719 24157
rect 23750 24148 23756 24200
rect 23808 24148 23814 24200
rect 24673 24191 24731 24197
rect 24673 24157 24685 24191
rect 24719 24188 24731 24191
rect 24946 24188 24952 24200
rect 24719 24160 24952 24188
rect 24719 24157 24731 24160
rect 24673 24151 24731 24157
rect 24946 24148 24952 24160
rect 25004 24148 25010 24200
rect 25130 24148 25136 24200
rect 25188 24148 25194 24200
rect 25041 24123 25099 24129
rect 25041 24120 25053 24123
rect 24780 24092 25053 24120
rect 24780 24064 24808 24092
rect 25041 24089 25053 24092
rect 25087 24089 25099 24123
rect 25240 24120 25268 24296
rect 26326 24284 26332 24336
rect 26384 24324 26390 24336
rect 26421 24327 26479 24333
rect 26421 24324 26433 24327
rect 26384 24296 26433 24324
rect 26384 24284 26390 24296
rect 26421 24293 26433 24296
rect 26467 24293 26479 24327
rect 26421 24287 26479 24293
rect 25590 24216 25596 24268
rect 25648 24256 25654 24268
rect 25869 24259 25927 24265
rect 25869 24256 25881 24259
rect 25648 24228 25881 24256
rect 25648 24216 25654 24228
rect 25869 24225 25881 24228
rect 25915 24225 25927 24259
rect 25869 24219 25927 24225
rect 25958 24216 25964 24268
rect 26016 24256 26022 24268
rect 26237 24259 26295 24265
rect 26237 24256 26249 24259
rect 26016 24228 26249 24256
rect 26016 24216 26022 24228
rect 26237 24225 26249 24228
rect 26283 24256 26295 24259
rect 26789 24259 26847 24265
rect 26789 24256 26801 24259
rect 26283 24228 26801 24256
rect 26283 24225 26295 24228
rect 26237 24219 26295 24225
rect 26789 24225 26801 24228
rect 26835 24256 26847 24259
rect 27154 24256 27160 24268
rect 26835 24228 27160 24256
rect 26835 24225 26847 24228
rect 26789 24219 26847 24225
rect 27154 24216 27160 24228
rect 27212 24216 27218 24268
rect 26878 24148 26884 24200
rect 26936 24148 26942 24200
rect 27062 24148 27068 24200
rect 27120 24148 27126 24200
rect 27338 24148 27344 24200
rect 27396 24188 27402 24200
rect 27525 24191 27583 24197
rect 27525 24188 27537 24191
rect 27396 24160 27537 24188
rect 27396 24148 27402 24160
rect 27525 24157 27537 24160
rect 27571 24157 27583 24191
rect 27525 24151 27583 24157
rect 25866 24120 25872 24132
rect 25240 24092 25872 24120
rect 25041 24083 25099 24089
rect 25866 24080 25872 24092
rect 25924 24120 25930 24132
rect 25924 24092 26372 24120
rect 25924 24080 25930 24092
rect 22244 24024 23152 24052
rect 22244 24012 22250 24024
rect 24486 24012 24492 24064
rect 24544 24012 24550 24064
rect 24762 24012 24768 24064
rect 24820 24012 24826 24064
rect 24854 24012 24860 24064
rect 24912 24012 24918 24064
rect 26050 24012 26056 24064
rect 26108 24012 26114 24064
rect 26344 24061 26372 24092
rect 26329 24055 26387 24061
rect 26329 24021 26341 24055
rect 26375 24052 26387 24055
rect 27062 24052 27068 24064
rect 26375 24024 27068 24052
rect 26375 24021 26387 24024
rect 26329 24015 26387 24021
rect 27062 24012 27068 24024
rect 27120 24012 27126 24064
rect 27706 24012 27712 24064
rect 27764 24012 27770 24064
rect 1104 23962 28152 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 28152 23962
rect 1104 23888 28152 23910
rect 4798 23808 4804 23860
rect 4856 23848 4862 23860
rect 4856 23820 6132 23848
rect 4856 23808 4862 23820
rect 2498 23740 2504 23792
rect 2556 23740 2562 23792
rect 4614 23780 4620 23792
rect 4540 23752 4620 23780
rect 2590 23712 2596 23724
rect 2438 23684 2596 23712
rect 2590 23672 2596 23684
rect 2648 23672 2654 23724
rect 4540 23721 4568 23752
rect 4614 23740 4620 23752
rect 4672 23740 4678 23792
rect 5626 23740 5632 23792
rect 5684 23740 5690 23792
rect 4525 23715 4583 23721
rect 4525 23681 4537 23715
rect 4571 23681 4583 23715
rect 4525 23675 4583 23681
rect 4706 23672 4712 23724
rect 4764 23672 4770 23724
rect 5537 23715 5595 23721
rect 5537 23681 5549 23715
rect 5583 23712 5595 23715
rect 5644 23712 5672 23740
rect 5583 23684 5672 23712
rect 5583 23681 5595 23684
rect 5537 23675 5595 23681
rect 5902 23672 5908 23724
rect 5960 23721 5966 23724
rect 5960 23715 5997 23721
rect 5985 23681 5997 23715
rect 6104 23712 6132 23820
rect 9214 23808 9220 23860
rect 9272 23808 9278 23860
rect 15654 23848 15660 23860
rect 13372 23820 15660 23848
rect 9398 23740 9404 23792
rect 9456 23740 9462 23792
rect 9769 23783 9827 23789
rect 9769 23749 9781 23783
rect 9815 23780 9827 23783
rect 10045 23783 10103 23789
rect 10045 23780 10057 23783
rect 9815 23752 10057 23780
rect 9815 23749 9827 23752
rect 9769 23743 9827 23749
rect 10045 23749 10057 23752
rect 10091 23780 10103 23783
rect 10870 23780 10876 23792
rect 10091 23752 10876 23780
rect 10091 23749 10103 23752
rect 10045 23743 10103 23749
rect 10870 23740 10876 23752
rect 10928 23740 10934 23792
rect 13372 23780 13400 23820
rect 15654 23808 15660 23820
rect 15712 23808 15718 23860
rect 18049 23851 18107 23857
rect 18049 23817 18061 23851
rect 18095 23848 18107 23851
rect 18230 23848 18236 23860
rect 18095 23820 18236 23848
rect 18095 23817 18107 23820
rect 18049 23811 18107 23817
rect 18230 23808 18236 23820
rect 18288 23808 18294 23860
rect 18877 23851 18935 23857
rect 18877 23817 18889 23851
rect 18923 23848 18935 23851
rect 20530 23848 20536 23860
rect 18923 23820 20536 23848
rect 18923 23817 18935 23820
rect 18877 23811 18935 23817
rect 20530 23808 20536 23820
rect 20588 23808 20594 23860
rect 21542 23808 21548 23860
rect 21600 23848 21606 23860
rect 23474 23848 23480 23860
rect 21600 23820 23480 23848
rect 21600 23808 21606 23820
rect 23474 23808 23480 23820
rect 23532 23808 23538 23860
rect 26142 23848 26148 23860
rect 25792 23820 26148 23848
rect 13280 23752 13400 23780
rect 7285 23715 7343 23721
rect 7285 23712 7297 23715
rect 6104 23684 7297 23712
rect 5960 23675 5997 23681
rect 7285 23681 7297 23684
rect 7331 23712 7343 23715
rect 7466 23712 7472 23724
rect 7331 23684 7472 23712
rect 7331 23681 7343 23684
rect 7285 23675 7343 23681
rect 5960 23672 5966 23675
rect 7466 23672 7472 23684
rect 7524 23672 7530 23724
rect 9030 23672 9036 23724
rect 9088 23712 9094 23724
rect 9125 23715 9183 23721
rect 9125 23712 9137 23715
rect 9088 23684 9137 23712
rect 9088 23672 9094 23684
rect 9125 23681 9137 23684
rect 9171 23681 9183 23715
rect 9125 23675 9183 23681
rect 9306 23672 9312 23724
rect 9364 23712 9370 23724
rect 9585 23715 9643 23721
rect 9585 23712 9597 23715
rect 9364 23684 9597 23712
rect 9364 23672 9370 23684
rect 9585 23681 9597 23684
rect 9631 23681 9643 23715
rect 9585 23675 9643 23681
rect 10226 23672 10232 23724
rect 10284 23672 10290 23724
rect 12253 23715 12311 23721
rect 12253 23681 12265 23715
rect 12299 23712 12311 23715
rect 12710 23712 12716 23724
rect 12299 23684 12716 23712
rect 12299 23681 12311 23684
rect 12253 23675 12311 23681
rect 12710 23672 12716 23684
rect 12768 23672 12774 23724
rect 12894 23672 12900 23724
rect 12952 23672 12958 23724
rect 13280 23721 13308 23752
rect 13538 23740 13544 23792
rect 13596 23740 13602 23792
rect 16390 23780 16396 23792
rect 14766 23766 16396 23780
rect 14752 23752 16396 23766
rect 13265 23715 13323 23721
rect 13265 23681 13277 23715
rect 13311 23681 13323 23715
rect 13265 23675 13323 23681
rect 1946 23604 1952 23656
rect 2004 23604 2010 23656
rect 5169 23647 5227 23653
rect 5169 23613 5181 23647
rect 5215 23644 5227 23647
rect 5258 23644 5264 23656
rect 5215 23616 5264 23644
rect 5215 23613 5227 23616
rect 5169 23607 5227 23613
rect 5258 23604 5264 23616
rect 5316 23604 5322 23656
rect 5629 23647 5687 23653
rect 5629 23613 5641 23647
rect 5675 23613 5687 23647
rect 5629 23607 5687 23613
rect 7377 23647 7435 23653
rect 7377 23613 7389 23647
rect 7423 23644 7435 23647
rect 7558 23644 7564 23656
rect 7423 23616 7564 23644
rect 7423 23613 7435 23616
rect 7377 23607 7435 23613
rect 1964 23576 1992 23604
rect 2774 23576 2780 23588
rect 1964 23548 2780 23576
rect 2774 23536 2780 23548
rect 2832 23536 2838 23588
rect 5534 23536 5540 23588
rect 5592 23576 5598 23588
rect 5644 23576 5672 23607
rect 7558 23604 7564 23616
rect 7616 23604 7622 23656
rect 9858 23604 9864 23656
rect 9916 23644 9922 23656
rect 11885 23647 11943 23653
rect 11885 23644 11897 23647
rect 9916 23616 11897 23644
rect 9916 23604 9922 23616
rect 11885 23613 11897 23616
rect 11931 23644 11943 23647
rect 12342 23644 12348 23656
rect 11931 23616 12348 23644
rect 11931 23613 11943 23616
rect 11885 23607 11943 23613
rect 12342 23604 12348 23616
rect 12400 23604 12406 23656
rect 12621 23647 12679 23653
rect 12621 23613 12633 23647
rect 12667 23644 12679 23647
rect 12802 23644 12808 23656
rect 12667 23616 12808 23644
rect 12667 23613 12679 23616
rect 12621 23607 12679 23613
rect 12802 23604 12808 23616
rect 12860 23604 12866 23656
rect 13538 23604 13544 23656
rect 13596 23644 13602 23656
rect 14752 23644 14780 23752
rect 16390 23740 16396 23752
rect 16448 23740 16454 23792
rect 17494 23740 17500 23792
rect 17552 23780 17558 23792
rect 18141 23783 18199 23789
rect 18141 23780 18153 23783
rect 17552 23752 18153 23780
rect 17552 23740 17558 23752
rect 18141 23749 18153 23752
rect 18187 23780 18199 23783
rect 18477 23783 18535 23789
rect 18477 23780 18489 23783
rect 18187 23752 18489 23780
rect 18187 23749 18199 23752
rect 18141 23743 18199 23749
rect 18477 23749 18489 23752
rect 18523 23749 18535 23783
rect 18477 23743 18535 23749
rect 18693 23783 18751 23789
rect 18693 23749 18705 23783
rect 18739 23749 18751 23783
rect 18693 23743 18751 23749
rect 15838 23672 15844 23724
rect 15896 23712 15902 23724
rect 15933 23715 15991 23721
rect 15933 23712 15945 23715
rect 15896 23684 15945 23712
rect 15896 23672 15902 23684
rect 15933 23681 15945 23684
rect 15979 23681 15991 23715
rect 15933 23675 15991 23681
rect 16114 23672 16120 23724
rect 16172 23672 16178 23724
rect 16761 23715 16819 23721
rect 16761 23681 16773 23715
rect 16807 23712 16819 23715
rect 17034 23712 17040 23724
rect 16807 23684 17040 23712
rect 16807 23681 16819 23684
rect 16761 23675 16819 23681
rect 17034 23672 17040 23684
rect 17092 23672 17098 23724
rect 17126 23672 17132 23724
rect 17184 23672 17190 23724
rect 17218 23672 17224 23724
rect 17276 23672 17282 23724
rect 17405 23715 17463 23721
rect 17405 23681 17417 23715
rect 17451 23681 17463 23715
rect 17405 23675 17463 23681
rect 17589 23715 17647 23721
rect 17589 23681 17601 23715
rect 17635 23712 17647 23715
rect 18046 23712 18052 23724
rect 17635 23684 18052 23712
rect 17635 23681 17647 23684
rect 17589 23675 17647 23681
rect 13596 23616 14780 23644
rect 17420 23644 17448 23675
rect 18046 23672 18052 23684
rect 18104 23672 18110 23724
rect 18233 23715 18291 23721
rect 18233 23681 18245 23715
rect 18279 23712 18291 23715
rect 18598 23712 18604 23724
rect 18279 23684 18604 23712
rect 18279 23681 18291 23684
rect 18233 23675 18291 23681
rect 18598 23672 18604 23684
rect 18656 23672 18662 23724
rect 17862 23644 17868 23656
rect 17420 23616 17868 23644
rect 13596 23604 13602 23616
rect 17862 23604 17868 23616
rect 17920 23644 17926 23656
rect 18708 23644 18736 23743
rect 19150 23740 19156 23792
rect 19208 23740 19214 23792
rect 20346 23740 20352 23792
rect 20404 23740 20410 23792
rect 21358 23740 21364 23792
rect 21416 23740 21422 23792
rect 22002 23740 22008 23792
rect 22060 23780 22066 23792
rect 25498 23780 25504 23792
rect 22060 23766 22126 23780
rect 22060 23752 22140 23766
rect 25254 23752 25504 23780
rect 22060 23740 22066 23752
rect 18782 23672 18788 23724
rect 18840 23672 18846 23724
rect 19058 23672 19064 23724
rect 19116 23672 19122 23724
rect 17920 23616 18736 23644
rect 17920 23604 17926 23616
rect 19886 23604 19892 23656
rect 19944 23604 19950 23656
rect 21634 23604 21640 23656
rect 21692 23604 21698 23656
rect 22112 23644 22140 23752
rect 25498 23740 25504 23752
rect 25556 23740 25562 23792
rect 25590 23672 25596 23724
rect 25648 23672 25654 23724
rect 25792 23721 25820 23820
rect 26142 23808 26148 23820
rect 26200 23808 26206 23860
rect 26237 23851 26295 23857
rect 26237 23817 26249 23851
rect 26283 23848 26295 23851
rect 26418 23848 26424 23860
rect 26283 23820 26424 23848
rect 26283 23817 26295 23820
rect 26237 23811 26295 23817
rect 26418 23808 26424 23820
rect 26476 23808 26482 23860
rect 25866 23740 25872 23792
rect 25924 23740 25930 23792
rect 25958 23740 25964 23792
rect 26016 23740 26022 23792
rect 25741 23715 25820 23721
rect 25741 23681 25753 23715
rect 25787 23684 25820 23715
rect 25787 23681 25799 23684
rect 25741 23675 25799 23681
rect 22554 23644 22560 23656
rect 22112 23616 22560 23644
rect 22554 23604 22560 23616
rect 22612 23604 22618 23656
rect 23290 23604 23296 23656
rect 23348 23604 23354 23656
rect 23566 23604 23572 23656
rect 23624 23644 23630 23656
rect 23753 23647 23811 23653
rect 23753 23644 23765 23647
rect 23624 23616 23765 23644
rect 23624 23604 23630 23616
rect 23753 23613 23765 23616
rect 23799 23613 23811 23647
rect 23753 23607 23811 23613
rect 24026 23604 24032 23656
rect 24084 23604 24090 23656
rect 25038 23604 25044 23656
rect 25096 23644 25102 23656
rect 25406 23644 25412 23656
rect 25096 23616 25412 23644
rect 25096 23604 25102 23616
rect 25406 23604 25412 23616
rect 25464 23644 25470 23656
rect 25501 23647 25559 23653
rect 25501 23644 25513 23647
rect 25464 23616 25513 23644
rect 25464 23604 25470 23616
rect 25501 23613 25513 23616
rect 25547 23644 25559 23647
rect 25976 23644 26004 23740
rect 26050 23672 26056 23724
rect 26108 23721 26114 23724
rect 26108 23712 26116 23721
rect 26108 23684 26153 23712
rect 26108 23675 26116 23684
rect 26108 23672 26114 23675
rect 26970 23672 26976 23724
rect 27028 23712 27034 23724
rect 27525 23715 27583 23721
rect 27525 23712 27537 23715
rect 27028 23684 27537 23712
rect 27028 23672 27034 23684
rect 27525 23681 27537 23684
rect 27571 23681 27583 23715
rect 27525 23675 27583 23681
rect 25547 23616 26004 23644
rect 25547 23613 25559 23616
rect 25501 23607 25559 23613
rect 5592 23548 5672 23576
rect 6181 23579 6239 23585
rect 5592 23536 5598 23548
rect 6181 23545 6193 23579
rect 6227 23576 6239 23579
rect 6914 23576 6920 23588
rect 6227 23548 6920 23576
rect 6227 23545 6239 23548
rect 6181 23539 6239 23545
rect 6914 23536 6920 23548
rect 6972 23536 6978 23588
rect 7653 23579 7711 23585
rect 7653 23545 7665 23579
rect 7699 23576 7711 23579
rect 8110 23576 8116 23588
rect 7699 23548 8116 23576
rect 7699 23545 7711 23548
rect 7653 23539 7711 23545
rect 8110 23536 8116 23548
rect 8168 23536 8174 23588
rect 13170 23536 13176 23588
rect 13228 23536 13234 23588
rect 16850 23536 16856 23588
rect 16908 23576 16914 23588
rect 17402 23576 17408 23588
rect 16908 23548 17408 23576
rect 16908 23536 16914 23548
rect 17402 23536 17408 23548
rect 17460 23536 17466 23588
rect 18230 23536 18236 23588
rect 18288 23576 18294 23588
rect 18288 23548 18552 23576
rect 18288 23536 18294 23548
rect 10413 23511 10471 23517
rect 10413 23477 10425 23511
rect 10459 23508 10471 23511
rect 10502 23508 10508 23520
rect 10459 23480 10508 23508
rect 10459 23477 10471 23480
rect 10413 23471 10471 23477
rect 10502 23468 10508 23480
rect 10560 23468 10566 23520
rect 15010 23468 15016 23520
rect 15068 23468 15074 23520
rect 15746 23468 15752 23520
rect 15804 23508 15810 23520
rect 16025 23511 16083 23517
rect 16025 23508 16037 23511
rect 15804 23480 16037 23508
rect 15804 23468 15810 23480
rect 16025 23477 16037 23480
rect 16071 23477 16083 23511
rect 16025 23471 16083 23477
rect 17126 23468 17132 23520
rect 17184 23508 17190 23520
rect 17773 23511 17831 23517
rect 17773 23508 17785 23511
rect 17184 23480 17785 23508
rect 17184 23468 17190 23480
rect 17773 23477 17785 23480
rect 17819 23477 17831 23511
rect 17773 23471 17831 23477
rect 17954 23468 17960 23520
rect 18012 23468 18018 23520
rect 18322 23468 18328 23520
rect 18380 23468 18386 23520
rect 18524 23517 18552 23548
rect 18509 23511 18567 23517
rect 18509 23477 18521 23511
rect 18555 23477 18567 23511
rect 18509 23471 18567 23477
rect 21821 23511 21879 23517
rect 21821 23477 21833 23511
rect 21867 23508 21879 23511
rect 21910 23508 21916 23520
rect 21867 23480 21916 23508
rect 21867 23477 21879 23480
rect 21821 23471 21879 23477
rect 21910 23468 21916 23480
rect 21968 23468 21974 23520
rect 27522 23468 27528 23520
rect 27580 23508 27586 23520
rect 27709 23511 27767 23517
rect 27709 23508 27721 23511
rect 27580 23480 27721 23508
rect 27580 23468 27586 23480
rect 27709 23477 27721 23480
rect 27755 23477 27767 23511
rect 27709 23471 27767 23477
rect 1104 23418 28152 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 28152 23418
rect 1104 23344 28152 23366
rect 7834 23264 7840 23316
rect 7892 23304 7898 23316
rect 8573 23307 8631 23313
rect 8573 23304 8585 23307
rect 7892 23276 8585 23304
rect 7892 23264 7898 23276
rect 8573 23273 8585 23276
rect 8619 23273 8631 23307
rect 9858 23304 9864 23316
rect 8573 23267 8631 23273
rect 9600 23276 9864 23304
rect 9600 23236 9628 23276
rect 9858 23264 9864 23276
rect 9916 23264 9922 23316
rect 9953 23307 10011 23313
rect 9953 23273 9965 23307
rect 9999 23304 10011 23307
rect 11974 23304 11980 23316
rect 9999 23276 11980 23304
rect 9999 23273 10011 23276
rect 9953 23267 10011 23273
rect 11974 23264 11980 23276
rect 12032 23264 12038 23316
rect 12253 23307 12311 23313
rect 12253 23273 12265 23307
rect 12299 23304 12311 23307
rect 12710 23304 12716 23316
rect 12299 23276 12716 23304
rect 12299 23273 12311 23276
rect 12253 23267 12311 23273
rect 12710 23264 12716 23276
rect 12768 23304 12774 23316
rect 12805 23307 12863 23313
rect 12805 23304 12817 23307
rect 12768 23276 12817 23304
rect 12768 23264 12774 23276
rect 12805 23273 12817 23276
rect 12851 23273 12863 23307
rect 12805 23267 12863 23273
rect 18046 23264 18052 23316
rect 18104 23304 18110 23316
rect 19245 23307 19303 23313
rect 19245 23304 19257 23307
rect 18104 23276 19257 23304
rect 18104 23264 18110 23276
rect 19245 23273 19257 23276
rect 19291 23273 19303 23307
rect 19245 23267 19303 23273
rect 22189 23307 22247 23313
rect 22189 23273 22201 23307
rect 22235 23273 22247 23307
rect 22189 23267 22247 23273
rect 2608 23208 9628 23236
rect 9677 23239 9735 23245
rect 842 23060 848 23112
rect 900 23100 906 23112
rect 2608 23109 2636 23208
rect 9677 23205 9689 23239
rect 9723 23236 9735 23239
rect 11425 23239 11483 23245
rect 9723 23208 10732 23236
rect 9723 23205 9735 23208
rect 9677 23199 9735 23205
rect 2682 23128 2688 23180
rect 2740 23168 2746 23180
rect 2740 23140 4200 23168
rect 2740 23128 2746 23140
rect 2976 23109 3004 23140
rect 1489 23103 1547 23109
rect 1489 23100 1501 23103
rect 900 23072 1501 23100
rect 900 23060 906 23072
rect 1489 23069 1501 23072
rect 1535 23069 1547 23103
rect 1489 23063 1547 23069
rect 1673 23103 1731 23109
rect 1673 23069 1685 23103
rect 1719 23100 1731 23103
rect 2593 23103 2651 23109
rect 2593 23100 2605 23103
rect 1719 23072 2605 23100
rect 1719 23069 1731 23072
rect 1673 23063 1731 23069
rect 2593 23069 2605 23072
rect 2639 23069 2651 23103
rect 2593 23063 2651 23069
rect 2777 23103 2835 23109
rect 2777 23069 2789 23103
rect 2823 23069 2835 23103
rect 2777 23063 2835 23069
rect 2961 23103 3019 23109
rect 2961 23069 2973 23103
rect 3007 23069 3019 23103
rect 2961 23063 3019 23069
rect 3053 23103 3111 23109
rect 3053 23069 3065 23103
rect 3099 23069 3111 23103
rect 3053 23063 3111 23069
rect 2130 22992 2136 23044
rect 2188 23032 2194 23044
rect 2792 23032 2820 23063
rect 2188 23004 2820 23032
rect 2869 23035 2927 23041
rect 2188 22992 2194 23004
rect 2869 23001 2881 23035
rect 2915 23032 2927 23035
rect 3068 23032 3096 23063
rect 3142 23060 3148 23112
rect 3200 23100 3206 23112
rect 3237 23103 3295 23109
rect 3237 23100 3249 23103
rect 3200 23072 3249 23100
rect 3200 23060 3206 23072
rect 3237 23069 3249 23072
rect 3283 23069 3295 23103
rect 3237 23063 3295 23069
rect 2915 23004 3096 23032
rect 2915 23001 2927 23004
rect 2869 22995 2927 23001
rect 2976 22976 3004 23004
rect 2314 22924 2320 22976
rect 2372 22964 2378 22976
rect 2682 22964 2688 22976
rect 2372 22936 2688 22964
rect 2372 22924 2378 22936
rect 2682 22924 2688 22936
rect 2740 22924 2746 22976
rect 2958 22924 2964 22976
rect 3016 22924 3022 22976
rect 3145 22967 3203 22973
rect 3145 22933 3157 22967
rect 3191 22964 3203 22967
rect 3786 22964 3792 22976
rect 3191 22936 3792 22964
rect 3191 22933 3203 22936
rect 3145 22927 3203 22933
rect 3786 22924 3792 22936
rect 3844 22924 3850 22976
rect 4172 22964 4200 23140
rect 4614 23128 4620 23180
rect 4672 23128 4678 23180
rect 4985 23171 5043 23177
rect 4985 23137 4997 23171
rect 5031 23168 5043 23171
rect 5445 23171 5503 23177
rect 5445 23168 5457 23171
rect 5031 23140 5457 23168
rect 5031 23137 5043 23140
rect 4985 23131 5043 23137
rect 5445 23137 5457 23140
rect 5491 23168 5503 23171
rect 5534 23168 5540 23180
rect 5491 23140 5540 23168
rect 5491 23137 5503 23140
rect 5445 23131 5503 23137
rect 5534 23128 5540 23140
rect 5592 23128 5598 23180
rect 9306 23128 9312 23180
rect 9364 23168 9370 23180
rect 10704 23168 10732 23208
rect 11425 23205 11437 23239
rect 11471 23236 11483 23239
rect 16850 23236 16856 23248
rect 11471 23208 16856 23236
rect 11471 23205 11483 23208
rect 11425 23199 11483 23205
rect 16850 23196 16856 23208
rect 16908 23196 16914 23248
rect 16945 23239 17003 23245
rect 16945 23205 16957 23239
rect 16991 23236 17003 23239
rect 18230 23236 18236 23248
rect 16991 23208 18236 23236
rect 16991 23205 17003 23208
rect 16945 23199 17003 23205
rect 18230 23196 18236 23208
rect 18288 23196 18294 23248
rect 22204 23236 22232 23267
rect 22278 23264 22284 23316
rect 22336 23304 22342 23316
rect 22373 23307 22431 23313
rect 22373 23304 22385 23307
rect 22336 23276 22385 23304
rect 22336 23264 22342 23276
rect 22373 23273 22385 23276
rect 22419 23273 22431 23307
rect 22373 23267 22431 23273
rect 22741 23307 22799 23313
rect 22741 23273 22753 23307
rect 22787 23304 22799 23307
rect 23290 23304 23296 23316
rect 22787 23276 23296 23304
rect 22787 23273 22799 23276
rect 22741 23267 22799 23273
rect 22204 23208 22324 23236
rect 22296 23180 22324 23208
rect 9364 23140 10180 23168
rect 9364 23128 9370 23140
rect 4632 23100 4660 23128
rect 4893 23103 4951 23109
rect 4893 23100 4905 23103
rect 4632 23072 4905 23100
rect 4893 23069 4905 23072
rect 4939 23069 4951 23103
rect 4893 23063 4951 23069
rect 5077 23103 5135 23109
rect 5077 23069 5089 23103
rect 5123 23069 5135 23103
rect 5077 23063 5135 23069
rect 4246 22992 4252 23044
rect 4304 23032 4310 23044
rect 4614 23032 4620 23044
rect 4304 23004 4620 23032
rect 4304 22992 4310 23004
rect 4614 22992 4620 23004
rect 4672 23032 4678 23044
rect 5092 23032 5120 23063
rect 5626 23060 5632 23112
rect 5684 23060 5690 23112
rect 6086 23060 6092 23112
rect 6144 23100 6150 23112
rect 6825 23103 6883 23109
rect 6144 23072 6776 23100
rect 6144 23060 6150 23072
rect 6748 23044 6776 23072
rect 6825 23069 6837 23103
rect 6871 23100 6883 23103
rect 6914 23100 6920 23112
rect 6871 23072 6920 23100
rect 6871 23069 6883 23072
rect 6825 23063 6883 23069
rect 6914 23060 6920 23072
rect 6972 23060 6978 23112
rect 7009 23103 7067 23109
rect 7009 23069 7021 23103
rect 7055 23069 7067 23103
rect 7009 23063 7067 23069
rect 4672 23004 5120 23032
rect 4672 22992 4678 23004
rect 6270 22992 6276 23044
rect 6328 22992 6334 23044
rect 6730 22992 6736 23044
rect 6788 23032 6794 23044
rect 7024 23032 7052 23063
rect 9030 23060 9036 23112
rect 9088 23100 9094 23112
rect 10152 23109 10180 23140
rect 10704 23140 11468 23168
rect 9585 23103 9643 23109
rect 9585 23100 9597 23103
rect 9088 23072 9597 23100
rect 9088 23060 9094 23072
rect 9585 23069 9597 23072
rect 9631 23069 9643 23103
rect 9585 23063 9643 23069
rect 10137 23103 10195 23109
rect 10137 23069 10149 23103
rect 10183 23069 10195 23103
rect 10137 23063 10195 23069
rect 10229 23103 10287 23109
rect 10229 23069 10241 23103
rect 10275 23069 10287 23103
rect 10229 23063 10287 23069
rect 6788 23004 7052 23032
rect 6788 22992 6794 23004
rect 7650 22992 7656 23044
rect 7708 22992 7714 23044
rect 8386 22992 8392 23044
rect 8444 22992 8450 23044
rect 10244 23032 10272 23063
rect 10410 23060 10416 23112
rect 10468 23060 10474 23112
rect 10502 23060 10508 23112
rect 10560 23060 10566 23112
rect 10594 23060 10600 23112
rect 10652 23060 10658 23112
rect 10704 23109 10732 23140
rect 10689 23103 10747 23109
rect 10689 23069 10701 23103
rect 10735 23069 10747 23103
rect 10689 23063 10747 23069
rect 10870 23060 10876 23112
rect 10928 23100 10934 23112
rect 11440 23109 11468 23140
rect 12158 23128 12164 23180
rect 12216 23168 12222 23180
rect 12216 23140 12756 23168
rect 12216 23128 12222 23140
rect 12728 23109 12756 23140
rect 12894 23128 12900 23180
rect 12952 23168 12958 23180
rect 12989 23171 13047 23177
rect 12989 23168 13001 23171
rect 12952 23140 13001 23168
rect 12952 23128 12958 23140
rect 12989 23137 13001 23140
rect 13035 23137 13047 23171
rect 12989 23131 13047 23137
rect 14182 23128 14188 23180
rect 14240 23168 14246 23180
rect 14550 23168 14556 23180
rect 14240 23140 14556 23168
rect 14240 23128 14246 23140
rect 14550 23128 14556 23140
rect 14608 23128 14614 23180
rect 22278 23128 22284 23180
rect 22336 23128 22342 23180
rect 11149 23103 11207 23109
rect 11149 23100 11161 23103
rect 10928 23072 11161 23100
rect 10928 23060 10934 23072
rect 11149 23069 11161 23072
rect 11195 23069 11207 23103
rect 11149 23063 11207 23069
rect 11425 23103 11483 23109
rect 11425 23069 11437 23103
rect 11471 23069 11483 23103
rect 11425 23063 11483 23069
rect 12437 23103 12495 23109
rect 12437 23069 12449 23103
rect 12483 23069 12495 23103
rect 12437 23063 12495 23069
rect 12713 23103 12771 23109
rect 12713 23069 12725 23103
rect 12759 23069 12771 23103
rect 12713 23063 12771 23069
rect 9600 23004 10272 23032
rect 10612 23032 10640 23060
rect 11333 23035 11391 23041
rect 11333 23032 11345 23035
rect 10612 23004 11345 23032
rect 9600 22976 9628 23004
rect 11333 23001 11345 23004
rect 11379 23001 11391 23035
rect 12452 23032 12480 23063
rect 12912 23032 12940 23128
rect 14277 23103 14335 23109
rect 14277 23069 14289 23103
rect 14323 23100 14335 23103
rect 15010 23100 15016 23112
rect 14323 23072 15016 23100
rect 14323 23069 14335 23072
rect 14277 23063 14335 23069
rect 15010 23060 15016 23072
rect 15068 23060 15074 23112
rect 15746 23060 15752 23112
rect 15804 23100 15810 23112
rect 16853 23103 16911 23109
rect 16853 23100 16865 23103
rect 15804 23072 16865 23100
rect 15804 23060 15810 23072
rect 16853 23069 16865 23072
rect 16899 23069 16911 23103
rect 16853 23063 16911 23069
rect 17034 23060 17040 23112
rect 17092 23060 17098 23112
rect 19426 23060 19432 23112
rect 19484 23060 19490 23112
rect 19705 23103 19763 23109
rect 19705 23069 19717 23103
rect 19751 23100 19763 23103
rect 21174 23100 21180 23112
rect 19751 23072 21180 23100
rect 19751 23069 19763 23072
rect 19705 23063 19763 23069
rect 21174 23060 21180 23072
rect 21232 23060 21238 23112
rect 21910 23060 21916 23112
rect 21968 23060 21974 23112
rect 22388 23100 22416 23267
rect 23290 23264 23296 23276
rect 23348 23264 23354 23316
rect 24026 23264 24032 23316
rect 24084 23304 24090 23316
rect 24121 23307 24179 23313
rect 24121 23304 24133 23307
rect 24084 23276 24133 23304
rect 24084 23264 24090 23276
rect 24121 23273 24133 23276
rect 24167 23273 24179 23307
rect 24121 23267 24179 23273
rect 25774 23264 25780 23316
rect 25832 23304 25838 23316
rect 26789 23307 26847 23313
rect 26789 23304 26801 23307
rect 25832 23276 26801 23304
rect 25832 23264 25838 23276
rect 26789 23273 26801 23276
rect 26835 23273 26847 23307
rect 26789 23267 26847 23273
rect 22649 23239 22707 23245
rect 22649 23205 22661 23239
rect 22695 23236 22707 23239
rect 22833 23239 22891 23245
rect 22833 23236 22845 23239
rect 22695 23208 22845 23236
rect 22695 23205 22707 23208
rect 22649 23199 22707 23205
rect 22833 23205 22845 23208
rect 22879 23205 22891 23239
rect 25590 23236 25596 23248
rect 22833 23199 22891 23205
rect 24872 23208 25596 23236
rect 22465 23171 22523 23177
rect 22465 23137 22477 23171
rect 22511 23168 22523 23171
rect 22922 23168 22928 23180
rect 22511 23140 22928 23168
rect 22511 23137 22523 23140
rect 22465 23131 22523 23137
rect 22922 23128 22928 23140
rect 22980 23168 22986 23180
rect 24397 23171 24455 23177
rect 22980 23140 23980 23168
rect 22980 23128 22986 23140
rect 22741 23103 22799 23109
rect 22741 23100 22753 23103
rect 22388 23072 22753 23100
rect 22741 23069 22753 23072
rect 22787 23069 22799 23103
rect 22020 23044 22140 23066
rect 22741 23063 22799 23069
rect 23106 23060 23112 23112
rect 23164 23060 23170 23112
rect 23952 23109 23980 23140
rect 24397 23137 24409 23171
rect 24443 23168 24455 23171
rect 24486 23168 24492 23180
rect 24443 23140 24492 23168
rect 24443 23137 24455 23140
rect 24397 23131 24455 23137
rect 24486 23128 24492 23140
rect 24544 23128 24550 23180
rect 24762 23128 24768 23180
rect 24820 23128 24826 23180
rect 24872 23177 24900 23208
rect 25590 23196 25596 23208
rect 25648 23196 25654 23248
rect 26804 23236 26832 23267
rect 26970 23264 26976 23316
rect 27028 23264 27034 23316
rect 27249 23239 27307 23245
rect 27249 23236 27261 23239
rect 26804 23208 27261 23236
rect 27249 23205 27261 23208
rect 27295 23205 27307 23239
rect 27249 23199 27307 23205
rect 24857 23171 24915 23177
rect 24857 23137 24869 23171
rect 24903 23137 24915 23171
rect 24857 23131 24915 23137
rect 26234 23128 26240 23180
rect 26292 23168 26298 23180
rect 26602 23168 26608 23180
rect 26292 23140 26608 23168
rect 26292 23128 26298 23140
rect 26602 23128 26608 23140
rect 26660 23168 26666 23180
rect 27065 23171 27123 23177
rect 27065 23168 27077 23171
rect 26660 23140 27077 23168
rect 26660 23128 26666 23140
rect 27065 23137 27077 23140
rect 27111 23137 27123 23171
rect 27065 23131 27123 23137
rect 23937 23103 23995 23109
rect 23937 23069 23949 23103
rect 23983 23100 23995 23103
rect 24121 23103 24179 23109
rect 23983 23072 24072 23100
rect 23983 23069 23995 23072
rect 23937 23063 23995 23069
rect 12452 23004 12940 23032
rect 11333 22995 11391 23001
rect 22002 22992 22008 23044
rect 22060 23038 22140 23044
rect 22060 22992 22066 23038
rect 22112 23032 22140 23038
rect 22646 23032 22652 23044
rect 22112 23004 22652 23032
rect 22646 22992 22652 23004
rect 22704 23032 22710 23044
rect 22833 23035 22891 23041
rect 22833 23032 22845 23035
rect 22704 23004 22845 23032
rect 22704 22992 22710 23004
rect 22833 23001 22845 23004
rect 22879 23001 22891 23035
rect 23124 23032 23152 23060
rect 22833 22995 22891 23001
rect 22940 23004 23152 23032
rect 6362 22964 6368 22976
rect 4172 22936 6368 22964
rect 6362 22924 6368 22936
rect 6420 22924 6426 22976
rect 8110 22924 8116 22976
rect 8168 22964 8174 22976
rect 8589 22967 8647 22973
rect 8589 22964 8601 22967
rect 8168 22936 8601 22964
rect 8168 22924 8174 22936
rect 8589 22933 8601 22936
rect 8635 22933 8647 22967
rect 8589 22927 8647 22933
rect 8757 22967 8815 22973
rect 8757 22933 8769 22967
rect 8803 22964 8815 22967
rect 8846 22964 8852 22976
rect 8803 22936 8852 22964
rect 8803 22933 8815 22936
rect 8757 22927 8815 22933
rect 8846 22924 8852 22936
rect 8904 22924 8910 22976
rect 9582 22924 9588 22976
rect 9640 22924 9646 22976
rect 11054 22924 11060 22976
rect 11112 22924 11118 22976
rect 12618 22924 12624 22976
rect 12676 22924 12682 22976
rect 12710 22924 12716 22976
rect 12768 22964 12774 22976
rect 12989 22967 13047 22973
rect 12989 22964 13001 22967
rect 12768 22936 13001 22964
rect 12768 22924 12774 22936
rect 12989 22933 13001 22936
rect 13035 22933 13047 22967
rect 12989 22927 13047 22933
rect 14642 22924 14648 22976
rect 14700 22924 14706 22976
rect 18414 22924 18420 22976
rect 18472 22964 18478 22976
rect 18874 22964 18880 22976
rect 18472 22936 18880 22964
rect 18472 22924 18478 22936
rect 18874 22924 18880 22936
rect 18932 22924 18938 22976
rect 19334 22924 19340 22976
rect 19392 22964 19398 22976
rect 19613 22967 19671 22973
rect 19613 22964 19625 22967
rect 19392 22936 19625 22964
rect 19392 22924 19398 22936
rect 19613 22933 19625 22936
rect 19659 22933 19671 22967
rect 19613 22927 19671 22933
rect 21729 22967 21787 22973
rect 21729 22933 21741 22967
rect 21775 22964 21787 22967
rect 22094 22964 22100 22976
rect 21775 22936 22100 22964
rect 21775 22933 21787 22936
rect 21729 22927 21787 22933
rect 22094 22924 22100 22936
rect 22152 22924 22158 22976
rect 22215 22967 22273 22973
rect 22215 22933 22227 22967
rect 22261 22964 22273 22967
rect 22940 22964 22968 23004
rect 22261 22936 22968 22964
rect 22261 22933 22273 22936
rect 22215 22927 22273 22933
rect 23014 22924 23020 22976
rect 23072 22924 23078 22976
rect 24044 22964 24072 23072
rect 24121 23069 24133 23103
rect 24167 23069 24179 23103
rect 24121 23063 24179 23069
rect 24136 23032 24164 23063
rect 24210 23060 24216 23112
rect 24268 23100 24274 23112
rect 24780 23100 24808 23128
rect 24268 23072 24808 23100
rect 24268 23060 24274 23072
rect 25406 23060 25412 23112
rect 25464 23060 25470 23112
rect 25593 23103 25651 23109
rect 25593 23069 25605 23103
rect 25639 23100 25651 23103
rect 26050 23100 26056 23112
rect 25639 23072 26056 23100
rect 25639 23069 25651 23072
rect 25593 23063 25651 23069
rect 26050 23060 26056 23072
rect 26108 23100 26114 23112
rect 27341 23103 27399 23109
rect 26108 23072 27200 23100
rect 26108 23060 26114 23072
rect 27172 23044 27200 23072
rect 27341 23069 27353 23103
rect 27387 23069 27399 23103
rect 27341 23063 27399 23069
rect 25041 23035 25099 23041
rect 25041 23032 25053 23035
rect 24136 23004 25053 23032
rect 25041 23001 25053 23004
rect 25087 23001 25099 23035
rect 25041 22995 25099 23001
rect 26602 22992 26608 23044
rect 26660 22992 26666 23044
rect 27154 22992 27160 23044
rect 27212 23032 27218 23044
rect 27356 23032 27384 23063
rect 27430 23060 27436 23112
rect 27488 23100 27494 23112
rect 27617 23103 27675 23109
rect 27617 23100 27629 23103
rect 27488 23072 27629 23100
rect 27488 23060 27494 23072
rect 27617 23069 27629 23072
rect 27663 23069 27675 23103
rect 27617 23063 27675 23069
rect 27212 23004 27384 23032
rect 27212 22992 27218 23004
rect 24854 22964 24860 22976
rect 24044 22936 24860 22964
rect 24854 22924 24860 22936
rect 24912 22924 24918 22976
rect 25406 22924 25412 22976
rect 25464 22924 25470 22976
rect 26142 22924 26148 22976
rect 26200 22964 26206 22976
rect 26805 22967 26863 22973
rect 26805 22964 26817 22967
rect 26200 22936 26817 22964
rect 26200 22924 26206 22936
rect 26805 22933 26817 22936
rect 26851 22933 26863 22967
rect 26805 22927 26863 22933
rect 27338 22924 27344 22976
rect 27396 22924 27402 22976
rect 27433 22967 27491 22973
rect 27433 22933 27445 22967
rect 27479 22964 27491 22967
rect 27522 22964 27528 22976
rect 27479 22936 27528 22964
rect 27479 22933 27491 22936
rect 27433 22927 27491 22933
rect 27522 22924 27528 22936
rect 27580 22924 27586 22976
rect 1104 22874 28152 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 28152 22874
rect 1104 22800 28152 22822
rect 2501 22763 2559 22769
rect 2501 22729 2513 22763
rect 2547 22760 2559 22763
rect 2866 22760 2872 22772
rect 2547 22732 2872 22760
rect 2547 22729 2559 22732
rect 2501 22723 2559 22729
rect 2866 22720 2872 22732
rect 2924 22720 2930 22772
rect 3973 22763 4031 22769
rect 3973 22729 3985 22763
rect 4019 22729 4031 22763
rect 3973 22723 4031 22729
rect 3786 22652 3792 22704
rect 3844 22652 3850 22704
rect 3988 22692 4016 22723
rect 4062 22720 4068 22772
rect 4120 22760 4126 22772
rect 6917 22763 6975 22769
rect 4120 22732 4384 22760
rect 4120 22720 4126 22732
rect 4246 22692 4252 22704
rect 3988 22664 4252 22692
rect 4246 22652 4252 22664
rect 4304 22652 4310 22704
rect 4356 22692 4384 22732
rect 6917 22729 6929 22763
rect 6963 22760 6975 22763
rect 7929 22763 7987 22769
rect 7929 22760 7941 22763
rect 6963 22732 7941 22760
rect 6963 22729 6975 22732
rect 6917 22723 6975 22729
rect 7929 22729 7941 22732
rect 7975 22760 7987 22763
rect 8386 22760 8392 22772
rect 7975 22732 8392 22760
rect 7975 22729 7987 22732
rect 7929 22723 7987 22729
rect 8386 22720 8392 22732
rect 8444 22720 8450 22772
rect 9582 22720 9588 22772
rect 9640 22760 9646 22772
rect 9677 22763 9735 22769
rect 9677 22760 9689 22763
rect 9640 22732 9689 22760
rect 9640 22720 9646 22732
rect 9677 22729 9689 22732
rect 9723 22729 9735 22763
rect 9677 22723 9735 22729
rect 10045 22763 10103 22769
rect 10045 22729 10057 22763
rect 10091 22760 10103 22763
rect 10594 22760 10600 22772
rect 10091 22732 10600 22760
rect 10091 22729 10103 22732
rect 10045 22723 10103 22729
rect 10594 22720 10600 22732
rect 10652 22720 10658 22772
rect 18414 22720 18420 22772
rect 18472 22720 18478 22772
rect 18874 22720 18880 22772
rect 18932 22720 18938 22772
rect 22278 22720 22284 22772
rect 22336 22760 22342 22772
rect 23014 22760 23020 22772
rect 22336 22732 23020 22760
rect 22336 22720 22342 22732
rect 23014 22720 23020 22732
rect 23072 22760 23078 22772
rect 25130 22760 25136 22772
rect 23072 22732 25136 22760
rect 23072 22720 23078 22732
rect 25130 22720 25136 22732
rect 25188 22720 25194 22772
rect 25317 22763 25375 22769
rect 25317 22760 25329 22763
rect 25240 22732 25329 22760
rect 7561 22695 7619 22701
rect 4356 22664 7512 22692
rect 7484 22636 7512 22664
rect 7561 22661 7573 22695
rect 7607 22692 7619 22695
rect 7607 22664 7880 22692
rect 7607 22661 7619 22664
rect 7561 22655 7619 22661
rect 7852 22636 7880 22664
rect 8110 22652 8116 22704
rect 8168 22652 8174 22704
rect 8846 22652 8852 22704
rect 8904 22652 8910 22704
rect 9217 22695 9275 22701
rect 9217 22661 9229 22695
rect 9263 22692 9275 22695
rect 9263 22664 9904 22692
rect 9263 22661 9275 22664
rect 9217 22655 9275 22661
rect 1857 22627 1915 22633
rect 1857 22593 1869 22627
rect 1903 22624 1915 22627
rect 2314 22624 2320 22636
rect 1903 22596 2320 22624
rect 1903 22593 1915 22596
rect 1857 22587 1915 22593
rect 2314 22584 2320 22596
rect 2372 22584 2378 22636
rect 3142 22584 3148 22636
rect 3200 22584 3206 22636
rect 4157 22627 4215 22633
rect 4157 22624 4169 22627
rect 3620 22596 4169 22624
rect 3620 22568 3648 22596
rect 4157 22593 4169 22596
rect 4203 22593 4215 22627
rect 4157 22587 4215 22593
rect 6730 22584 6736 22636
rect 6788 22584 6794 22636
rect 6914 22584 6920 22636
rect 6972 22584 6978 22636
rect 7466 22584 7472 22636
rect 7524 22584 7530 22636
rect 7650 22584 7656 22636
rect 7708 22584 7714 22636
rect 7834 22584 7840 22636
rect 7892 22584 7898 22636
rect 9030 22624 9036 22636
rect 8128 22596 9036 22624
rect 1949 22559 2007 22565
rect 1949 22525 1961 22559
rect 1995 22556 2007 22559
rect 2130 22556 2136 22568
rect 1995 22528 2136 22556
rect 1995 22525 2007 22528
rect 1949 22519 2007 22525
rect 2130 22516 2136 22528
rect 2188 22516 2194 22568
rect 2869 22559 2927 22565
rect 2869 22525 2881 22559
rect 2915 22556 2927 22559
rect 2958 22556 2964 22568
rect 2915 22528 2964 22556
rect 2915 22525 2927 22528
rect 2869 22519 2927 22525
rect 2958 22516 2964 22528
rect 3016 22516 3022 22568
rect 3602 22516 3608 22568
rect 3660 22516 3666 22568
rect 4341 22491 4399 22497
rect 4341 22457 4353 22491
rect 4387 22488 4399 22491
rect 4798 22488 4804 22500
rect 4387 22460 4804 22488
rect 4387 22457 4399 22460
rect 4341 22451 4399 22457
rect 4798 22448 4804 22460
rect 4856 22448 4862 22500
rect 8128 22497 8156 22596
rect 9030 22584 9036 22596
rect 9088 22584 9094 22636
rect 9306 22584 9312 22636
rect 9364 22624 9370 22636
rect 9876 22633 9904 22664
rect 11054 22652 11060 22704
rect 11112 22692 11118 22704
rect 18432 22692 18460 22720
rect 18601 22695 18659 22701
rect 18601 22692 18613 22695
rect 11112 22664 18613 22692
rect 11112 22652 11118 22664
rect 9585 22627 9643 22633
rect 9585 22624 9597 22627
rect 9364 22596 9597 22624
rect 9364 22584 9370 22596
rect 9585 22593 9597 22596
rect 9631 22593 9643 22627
rect 9585 22587 9643 22593
rect 9861 22627 9919 22633
rect 9861 22593 9873 22627
rect 9907 22624 9919 22627
rect 10226 22624 10232 22636
rect 9907 22596 10232 22624
rect 9907 22593 9919 22596
rect 9861 22587 9919 22593
rect 10226 22584 10232 22596
rect 10284 22584 10290 22636
rect 12618 22584 12624 22636
rect 12676 22584 12682 22636
rect 12805 22627 12863 22633
rect 12805 22593 12817 22627
rect 12851 22624 12863 22627
rect 13170 22624 13176 22636
rect 12851 22596 13176 22624
rect 12851 22593 12863 22596
rect 12805 22587 12863 22593
rect 13170 22584 13176 22596
rect 13228 22584 13234 22636
rect 18156 22633 18184 22664
rect 18601 22661 18613 22664
rect 18647 22661 18659 22695
rect 18601 22655 18659 22661
rect 18690 22652 18696 22704
rect 18748 22652 18754 22704
rect 19337 22695 19395 22701
rect 19337 22661 19349 22695
rect 19383 22692 19395 22695
rect 20257 22695 20315 22701
rect 20257 22692 20269 22695
rect 19383 22664 20269 22692
rect 19383 22661 19395 22664
rect 19337 22655 19395 22661
rect 20257 22661 20269 22664
rect 20303 22661 20315 22695
rect 20257 22655 20315 22661
rect 22002 22652 22008 22704
rect 22060 22692 22066 22704
rect 22189 22695 22247 22701
rect 22189 22692 22201 22695
rect 22060 22664 22201 22692
rect 22060 22652 22066 22664
rect 22189 22661 22201 22664
rect 22235 22661 22247 22695
rect 22189 22655 22247 22661
rect 22370 22652 22376 22704
rect 22428 22652 22434 22704
rect 25240 22701 25268 22732
rect 25317 22729 25329 22732
rect 25363 22760 25375 22763
rect 25590 22760 25596 22772
rect 25363 22732 25596 22760
rect 25363 22729 25375 22732
rect 25317 22723 25375 22729
rect 25590 22720 25596 22732
rect 25648 22720 25654 22772
rect 26142 22720 26148 22772
rect 26200 22760 26206 22772
rect 26237 22763 26295 22769
rect 26237 22760 26249 22763
rect 26200 22732 26249 22760
rect 26200 22720 26206 22732
rect 26237 22729 26249 22732
rect 26283 22729 26295 22763
rect 26237 22723 26295 22729
rect 27154 22720 27160 22772
rect 27212 22720 27218 22772
rect 27522 22760 27528 22772
rect 27264 22732 27528 22760
rect 25225 22695 25283 22701
rect 25225 22661 25237 22695
rect 25271 22661 25283 22695
rect 25225 22655 25283 22661
rect 25485 22695 25543 22701
rect 25485 22661 25497 22695
rect 25531 22692 25543 22695
rect 25531 22664 25636 22692
rect 25531 22661 25543 22664
rect 25485 22655 25543 22661
rect 18691 22649 18749 22652
rect 18141 22627 18199 22633
rect 18141 22593 18153 22627
rect 18187 22593 18199 22627
rect 18141 22587 18199 22593
rect 18325 22627 18383 22633
rect 18325 22593 18337 22627
rect 18371 22624 18383 22627
rect 18417 22627 18475 22633
rect 18417 22624 18429 22627
rect 18371 22596 18429 22624
rect 18371 22593 18383 22596
rect 18325 22587 18383 22593
rect 18417 22593 18429 22596
rect 18463 22593 18475 22627
rect 18691 22615 18703 22649
rect 18737 22615 18749 22649
rect 18691 22609 18749 22615
rect 18785 22633 18843 22639
rect 18785 22599 18797 22633
rect 18831 22622 18843 22633
rect 18874 22622 18880 22636
rect 18831 22599 18880 22622
rect 18785 22594 18880 22599
rect 18785 22593 18843 22594
rect 18417 22587 18475 22593
rect 12529 22559 12587 22565
rect 12529 22556 12541 22559
rect 12406 22528 12541 22556
rect 8113 22491 8171 22497
rect 8113 22457 8125 22491
rect 8159 22457 8171 22491
rect 8113 22451 8171 22457
rect 3878 22380 3884 22432
rect 3936 22420 3942 22432
rect 12406 22420 12434 22528
rect 12529 22525 12541 22528
rect 12575 22525 12587 22559
rect 12529 22519 12587 22525
rect 16850 22516 16856 22568
rect 16908 22556 16914 22568
rect 18340 22556 18368 22587
rect 18874 22584 18880 22594
rect 18932 22584 18938 22636
rect 18966 22584 18972 22636
rect 19024 22624 19030 22636
rect 19061 22627 19119 22633
rect 19061 22624 19073 22627
rect 19024 22596 19073 22624
rect 19024 22584 19030 22596
rect 19061 22593 19073 22596
rect 19107 22624 19119 22627
rect 19518 22624 19524 22636
rect 19107 22596 19524 22624
rect 19107 22593 19119 22596
rect 19061 22587 19119 22593
rect 19518 22584 19524 22596
rect 19576 22584 19582 22636
rect 20165 22627 20223 22633
rect 20165 22593 20177 22627
rect 20211 22593 20223 22627
rect 20165 22587 20223 22593
rect 20349 22627 20407 22633
rect 20349 22593 20361 22627
rect 20395 22624 20407 22627
rect 20714 22624 20720 22636
rect 20395 22596 20720 22624
rect 20395 22593 20407 22596
rect 20349 22587 20407 22593
rect 16908 22528 18368 22556
rect 20180 22556 20208 22587
rect 20714 22584 20720 22596
rect 20772 22584 20778 22636
rect 25608 22624 25636 22664
rect 25682 22652 25688 22704
rect 25740 22692 25746 22704
rect 26050 22692 26056 22704
rect 25740 22664 26056 22692
rect 25740 22652 25746 22664
rect 26050 22652 26056 22664
rect 26108 22652 26114 22704
rect 25958 22624 25964 22636
rect 25608 22596 25964 22624
rect 25958 22584 25964 22596
rect 26016 22624 26022 22636
rect 26160 22624 26188 22720
rect 27172 22692 27200 22720
rect 26344 22664 27200 22692
rect 26344 22633 26372 22664
rect 26016 22596 26188 22624
rect 26329 22627 26387 22633
rect 26016 22584 26022 22596
rect 26329 22593 26341 22627
rect 26375 22593 26387 22627
rect 26329 22587 26387 22593
rect 27062 22584 27068 22636
rect 27120 22624 27126 22636
rect 27157 22627 27215 22633
rect 27157 22624 27169 22627
rect 27120 22596 27169 22624
rect 27120 22584 27126 22596
rect 27157 22593 27169 22596
rect 27203 22593 27215 22627
rect 27157 22587 27215 22593
rect 21174 22556 21180 22568
rect 20180 22528 21180 22556
rect 16908 22516 16914 22528
rect 18340 22488 18368 22528
rect 21174 22516 21180 22528
rect 21232 22516 21238 22568
rect 23106 22516 23112 22568
rect 23164 22556 23170 22568
rect 24765 22559 24823 22565
rect 24765 22556 24777 22559
rect 23164 22528 24777 22556
rect 23164 22516 23170 22528
rect 24765 22525 24777 22528
rect 24811 22556 24823 22559
rect 25590 22556 25596 22568
rect 24811 22528 25596 22556
rect 24811 22525 24823 22528
rect 24765 22519 24823 22525
rect 25590 22516 25596 22528
rect 25648 22516 25654 22568
rect 26142 22516 26148 22568
rect 26200 22556 26206 22568
rect 26973 22559 27031 22565
rect 26973 22556 26985 22559
rect 26200 22528 26985 22556
rect 26200 22516 26206 22528
rect 26973 22525 26985 22528
rect 27019 22556 27031 22559
rect 27264 22556 27292 22732
rect 27522 22720 27528 22732
rect 27580 22720 27586 22772
rect 27338 22584 27344 22636
rect 27396 22624 27402 22636
rect 27525 22627 27583 22633
rect 27525 22624 27537 22627
rect 27396 22596 27537 22624
rect 27396 22584 27402 22596
rect 27525 22593 27537 22596
rect 27571 22593 27583 22627
rect 27525 22587 27583 22593
rect 27019 22528 27292 22556
rect 27019 22525 27031 22528
rect 26973 22519 27031 22525
rect 18874 22488 18880 22500
rect 18340 22460 18880 22488
rect 18874 22448 18880 22460
rect 18932 22448 18938 22500
rect 19061 22491 19119 22497
rect 19061 22457 19073 22491
rect 19107 22488 19119 22491
rect 19426 22488 19432 22500
rect 19107 22460 19432 22488
rect 19107 22457 19119 22460
rect 19061 22451 19119 22457
rect 19426 22448 19432 22460
rect 19484 22488 19490 22500
rect 19705 22491 19763 22497
rect 19705 22488 19717 22491
rect 19484 22460 19717 22488
rect 19484 22448 19490 22460
rect 19705 22457 19717 22460
rect 19751 22457 19763 22491
rect 19705 22451 19763 22457
rect 24670 22448 24676 22500
rect 24728 22488 24734 22500
rect 24728 22460 24900 22488
rect 24728 22448 24734 22460
rect 3936 22392 12434 22420
rect 12989 22423 13047 22429
rect 3936 22380 3942 22392
rect 12989 22389 13001 22423
rect 13035 22420 13047 22423
rect 14182 22420 14188 22432
rect 13035 22392 14188 22420
rect 13035 22389 13047 22392
rect 12989 22383 13047 22389
rect 14182 22380 14188 22392
rect 14240 22380 14246 22432
rect 18230 22380 18236 22432
rect 18288 22380 18294 22432
rect 18414 22380 18420 22432
rect 18472 22420 18478 22432
rect 18509 22423 18567 22429
rect 18509 22420 18521 22423
rect 18472 22392 18521 22420
rect 18472 22380 18478 22392
rect 18509 22389 18521 22392
rect 18555 22389 18567 22423
rect 18509 22383 18567 22389
rect 18598 22380 18604 22432
rect 18656 22420 18662 22432
rect 19153 22423 19211 22429
rect 19153 22420 19165 22423
rect 18656 22392 19165 22420
rect 18656 22380 18662 22392
rect 19153 22389 19165 22392
rect 19199 22389 19211 22423
rect 19153 22383 19211 22389
rect 19334 22380 19340 22432
rect 19392 22380 19398 22432
rect 24872 22420 24900 22460
rect 24946 22448 24952 22500
rect 25004 22448 25010 22500
rect 25222 22448 25228 22500
rect 25280 22488 25286 22500
rect 25682 22488 25688 22500
rect 25280 22460 25688 22488
rect 25280 22448 25286 22460
rect 25682 22448 25688 22460
rect 25740 22448 25746 22500
rect 27706 22448 27712 22500
rect 27764 22448 27770 22500
rect 25501 22423 25559 22429
rect 25501 22420 25513 22423
rect 24872 22392 25513 22420
rect 25501 22389 25513 22392
rect 25547 22420 25559 22423
rect 25774 22420 25780 22432
rect 25547 22392 25780 22420
rect 25547 22389 25559 22392
rect 25501 22383 25559 22389
rect 25774 22380 25780 22392
rect 25832 22420 25838 22432
rect 26050 22420 26056 22432
rect 25832 22392 26056 22420
rect 25832 22380 25838 22392
rect 26050 22380 26056 22392
rect 26108 22380 26114 22432
rect 27341 22423 27399 22429
rect 27341 22389 27353 22423
rect 27387 22420 27399 22423
rect 27522 22420 27528 22432
rect 27387 22392 27528 22420
rect 27387 22389 27399 22392
rect 27341 22383 27399 22389
rect 27522 22380 27528 22392
rect 27580 22380 27586 22432
rect 1104 22330 28152 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 28152 22330
rect 1104 22256 28152 22278
rect 12618 22176 12624 22228
rect 12676 22176 12682 22228
rect 14274 22176 14280 22228
rect 14332 22216 14338 22228
rect 14645 22219 14703 22225
rect 14645 22216 14657 22219
rect 14332 22188 14657 22216
rect 14332 22176 14338 22188
rect 14645 22185 14657 22188
rect 14691 22185 14703 22219
rect 14645 22179 14703 22185
rect 17129 22219 17187 22225
rect 17129 22185 17141 22219
rect 17175 22216 17187 22219
rect 17218 22216 17224 22228
rect 17175 22188 17224 22216
rect 17175 22185 17187 22188
rect 17129 22179 17187 22185
rect 17218 22176 17224 22188
rect 17276 22176 17282 22228
rect 21174 22176 21180 22228
rect 21232 22176 21238 22228
rect 24029 22219 24087 22225
rect 24029 22185 24041 22219
rect 24075 22216 24087 22219
rect 24210 22216 24216 22228
rect 24075 22188 24216 22216
rect 24075 22185 24087 22188
rect 24029 22179 24087 22185
rect 24210 22176 24216 22188
rect 24268 22176 24274 22228
rect 25222 22216 25228 22228
rect 24412 22188 25228 22216
rect 4062 22148 4068 22160
rect 2516 22120 4068 22148
rect 2314 22040 2320 22092
rect 2372 22080 2378 22092
rect 2516 22080 2544 22120
rect 4062 22108 4068 22120
rect 4120 22108 4126 22160
rect 10796 22120 20944 22148
rect 3053 22083 3111 22089
rect 3053 22080 3065 22083
rect 2372 22052 2544 22080
rect 2372 22040 2378 22052
rect 1394 21972 1400 22024
rect 1452 21972 1458 22024
rect 2516 21998 2544 22052
rect 2700 22052 3065 22080
rect 2700 22024 2728 22052
rect 3053 22049 3065 22052
rect 3099 22080 3111 22083
rect 9493 22083 9551 22089
rect 3099 22052 4384 22080
rect 3099 22049 3111 22052
rect 3053 22043 3111 22049
rect 2682 21972 2688 22024
rect 2740 21972 2746 22024
rect 2866 21972 2872 22024
rect 2924 21972 2930 22024
rect 3973 22015 4031 22021
rect 3973 21981 3985 22015
rect 4019 21981 4031 22015
rect 3973 21975 4031 21981
rect 1949 21947 2007 21953
rect 1949 21913 1961 21947
rect 1995 21944 2007 21947
rect 2130 21944 2136 21956
rect 1995 21916 2136 21944
rect 1995 21913 2007 21916
rect 1949 21907 2007 21913
rect 2130 21904 2136 21916
rect 2188 21904 2194 21956
rect 3988 21944 4016 21975
rect 4062 21972 4068 22024
rect 4120 22012 4126 22024
rect 4356 22021 4384 22052
rect 9493 22049 9505 22083
rect 9539 22080 9551 22083
rect 9861 22083 9919 22089
rect 9861 22080 9873 22083
rect 9539 22052 9873 22080
rect 9539 22049 9551 22052
rect 9493 22043 9551 22049
rect 9861 22049 9873 22052
rect 9907 22049 9919 22083
rect 9861 22043 9919 22049
rect 10689 22083 10747 22089
rect 10689 22049 10701 22083
rect 10735 22080 10747 22083
rect 10796 22080 10824 22120
rect 10735 22052 10824 22080
rect 11900 22052 12480 22080
rect 10735 22049 10747 22052
rect 10689 22043 10747 22049
rect 11900 22024 11928 22052
rect 4167 22015 4225 22021
rect 4167 22012 4179 22015
rect 4120 21984 4179 22012
rect 4120 21972 4126 21984
rect 4167 21981 4179 21984
rect 4213 21981 4225 22015
rect 4167 21975 4225 21981
rect 4341 22015 4399 22021
rect 4341 21981 4353 22015
rect 4387 21981 4399 22015
rect 4341 21975 4399 21981
rect 4798 21972 4804 22024
rect 4856 21972 4862 22024
rect 5258 21972 5264 22024
rect 5316 21972 5322 22024
rect 9306 21972 9312 22024
rect 9364 22012 9370 22024
rect 9401 22015 9459 22021
rect 9401 22012 9413 22015
rect 9364 21984 9413 22012
rect 9364 21972 9370 21984
rect 9401 21981 9413 21984
rect 9447 21981 9459 22015
rect 9401 21975 9459 21981
rect 9582 21972 9588 22024
rect 9640 21972 9646 22024
rect 10137 22015 10195 22021
rect 10137 21981 10149 22015
rect 10183 22012 10195 22015
rect 10226 22012 10232 22024
rect 10183 21984 10232 22012
rect 10183 21981 10195 21984
rect 10137 21975 10195 21981
rect 10226 21972 10232 21984
rect 10284 21972 10290 22024
rect 11609 22015 11667 22021
rect 11609 21981 11621 22015
rect 11655 21981 11667 22015
rect 11609 21975 11667 21981
rect 11793 22015 11851 22021
rect 11793 21981 11805 22015
rect 11839 22012 11851 22015
rect 11882 22012 11888 22024
rect 11839 21984 11888 22012
rect 11839 21981 11851 21984
rect 11793 21975 11851 21981
rect 3988 21916 4476 21944
rect 1581 21879 1639 21885
rect 1581 21845 1593 21879
rect 1627 21876 1639 21879
rect 3050 21876 3056 21888
rect 1627 21848 3056 21876
rect 1627 21845 1639 21848
rect 1581 21839 1639 21845
rect 3050 21836 3056 21848
rect 3108 21876 3114 21888
rect 3878 21876 3884 21888
rect 3108 21848 3884 21876
rect 3108 21836 3114 21848
rect 3878 21836 3884 21848
rect 3936 21836 3942 21888
rect 3970 21836 3976 21888
rect 4028 21836 4034 21888
rect 4448 21885 4476 21916
rect 6086 21904 6092 21956
rect 6144 21904 6150 21956
rect 11624 21944 11652 21975
rect 11882 21972 11888 21984
rect 11940 21972 11946 22024
rect 12158 21972 12164 22024
rect 12216 21972 12222 22024
rect 12452 22021 12480 22052
rect 14366 22040 14372 22092
rect 14424 22080 14430 22092
rect 14734 22080 14740 22092
rect 14424 22052 14740 22080
rect 14424 22040 14430 22052
rect 14734 22040 14740 22052
rect 14792 22040 14798 22092
rect 16206 22040 16212 22092
rect 16264 22080 16270 22092
rect 16264 22052 17080 22080
rect 16264 22040 16270 22052
rect 12437 22015 12495 22021
rect 12437 21981 12449 22015
rect 12483 21981 12495 22015
rect 12437 21975 12495 21981
rect 12526 21972 12532 22024
rect 12584 22012 12590 22024
rect 12713 22015 12771 22021
rect 12713 22012 12725 22015
rect 12584 21984 12725 22012
rect 12584 21972 12590 21984
rect 12713 21981 12725 21984
rect 12759 21981 12771 22015
rect 12713 21975 12771 21981
rect 14921 22015 14979 22021
rect 14921 21981 14933 22015
rect 14967 22012 14979 22015
rect 15010 22012 15016 22024
rect 14967 21984 15016 22012
rect 14967 21981 14979 21984
rect 14921 21975 14979 21981
rect 15010 21972 15016 21984
rect 15068 21972 15074 22024
rect 15105 22015 15163 22021
rect 15105 21981 15117 22015
rect 15151 22012 15163 22015
rect 15286 22012 15292 22024
rect 15151 21984 15292 22012
rect 15151 21981 15163 21984
rect 15105 21975 15163 21981
rect 15286 21972 15292 21984
rect 15344 22012 15350 22024
rect 15344 21984 16988 22012
rect 15344 21972 15350 21984
rect 12345 21947 12403 21953
rect 11624 21916 12020 21944
rect 4433 21879 4491 21885
rect 4433 21845 4445 21879
rect 4479 21876 4491 21879
rect 4614 21876 4620 21888
rect 4479 21848 4620 21876
rect 4479 21845 4491 21848
rect 4433 21839 4491 21845
rect 4614 21836 4620 21848
rect 4672 21836 4678 21888
rect 11698 21836 11704 21888
rect 11756 21836 11762 21888
rect 11992 21885 12020 21916
rect 12345 21913 12357 21947
rect 12391 21944 12403 21947
rect 14274 21944 14280 21956
rect 12391 21916 14280 21944
rect 12391 21913 12403 21916
rect 12345 21907 12403 21913
rect 14274 21904 14280 21916
rect 14332 21904 14338 21956
rect 14461 21947 14519 21953
rect 14461 21944 14473 21947
rect 14384 21916 14473 21944
rect 11977 21879 12035 21885
rect 11977 21845 11989 21879
rect 12023 21876 12035 21879
rect 12710 21876 12716 21888
rect 12023 21848 12716 21876
rect 12023 21845 12035 21848
rect 11977 21839 12035 21845
rect 12710 21836 12716 21848
rect 12768 21836 12774 21888
rect 12989 21879 13047 21885
rect 12989 21845 13001 21879
rect 13035 21876 13047 21879
rect 14090 21876 14096 21888
rect 13035 21848 14096 21876
rect 13035 21845 13047 21848
rect 12989 21839 13047 21845
rect 14090 21836 14096 21848
rect 14148 21876 14154 21888
rect 14384 21876 14412 21916
rect 14461 21913 14473 21916
rect 14507 21913 14519 21947
rect 14461 21907 14519 21913
rect 14642 21904 14648 21956
rect 14700 21953 14706 21956
rect 14700 21947 14719 21953
rect 14707 21913 14719 21947
rect 14700 21907 14719 21913
rect 14752 21916 15056 21944
rect 14700 21904 14706 21907
rect 14148 21848 14412 21876
rect 14148 21836 14154 21848
rect 14550 21836 14556 21888
rect 14608 21876 14614 21888
rect 14752 21876 14780 21916
rect 14608 21848 14780 21876
rect 14608 21836 14614 21848
rect 14826 21836 14832 21888
rect 14884 21836 14890 21888
rect 15028 21885 15056 21916
rect 16960 21888 16988 21984
rect 17052 21944 17080 22052
rect 17218 22040 17224 22092
rect 17276 22080 17282 22092
rect 19058 22080 19064 22092
rect 17276 22052 19064 22080
rect 17276 22040 17282 22052
rect 19058 22040 19064 22052
rect 19116 22040 19122 22092
rect 20714 22040 20720 22092
rect 20772 22040 20778 22092
rect 20916 22021 20944 22120
rect 21085 22083 21143 22089
rect 21085 22049 21097 22083
rect 21131 22080 21143 22083
rect 24412 22080 24440 22188
rect 25222 22176 25228 22188
rect 25280 22176 25286 22228
rect 25314 22176 25320 22228
rect 25372 22216 25378 22228
rect 25501 22219 25559 22225
rect 25501 22216 25513 22219
rect 25372 22188 25513 22216
rect 25372 22176 25378 22188
rect 25501 22185 25513 22188
rect 25547 22216 25559 22219
rect 25777 22219 25835 22225
rect 25777 22216 25789 22219
rect 25547 22188 25789 22216
rect 25547 22185 25559 22188
rect 25501 22179 25559 22185
rect 25777 22185 25789 22188
rect 25823 22185 25835 22219
rect 25777 22179 25835 22185
rect 25406 22148 25412 22160
rect 21131 22052 21404 22080
rect 21131 22049 21143 22052
rect 21085 22043 21143 22049
rect 21376 22021 21404 22052
rect 23952 22052 24440 22080
rect 24504 22120 25412 22148
rect 20901 22015 20959 22021
rect 20901 21981 20913 22015
rect 20947 22012 20959 22015
rect 21177 22015 21235 22021
rect 21177 22012 21189 22015
rect 20947 21984 21189 22012
rect 20947 21981 20959 21984
rect 20901 21975 20959 21981
rect 21100 21956 21128 21984
rect 21177 21981 21189 21984
rect 21223 21981 21235 22015
rect 21177 21975 21235 21981
rect 21361 22015 21419 22021
rect 21361 21981 21373 22015
rect 21407 22012 21419 22015
rect 22186 22012 22192 22024
rect 21407 21984 22192 22012
rect 21407 21981 21419 21984
rect 21361 21975 21419 21981
rect 22186 21972 22192 21984
rect 22244 21972 22250 22024
rect 17108 21947 17166 21953
rect 17108 21944 17120 21947
rect 17052 21916 17120 21944
rect 17108 21913 17120 21916
rect 17154 21944 17166 21947
rect 17154 21916 17264 21944
rect 17154 21913 17166 21916
rect 17108 21907 17166 21913
rect 15013 21879 15071 21885
rect 15013 21845 15025 21879
rect 15059 21845 15071 21879
rect 15013 21839 15071 21845
rect 16942 21836 16948 21888
rect 17000 21836 17006 21888
rect 17236 21876 17264 21916
rect 17310 21904 17316 21956
rect 17368 21904 17374 21956
rect 21082 21904 21088 21956
rect 21140 21904 21146 21956
rect 23845 21947 23903 21953
rect 23845 21913 23857 21947
rect 23891 21944 23903 21947
rect 23952 21944 23980 22052
rect 24504 21944 24532 22120
rect 25406 22108 25412 22120
rect 25464 22148 25470 22160
rect 25869 22151 25927 22157
rect 25464 22120 25820 22148
rect 25464 22108 25470 22120
rect 25682 22080 25688 22092
rect 24964 22052 25688 22080
rect 24578 21972 24584 22024
rect 24636 21972 24642 22024
rect 24670 21972 24676 22024
rect 24728 21972 24734 22024
rect 24854 21972 24860 22024
rect 24912 22012 24918 22024
rect 24964 22012 24992 22052
rect 25682 22040 25688 22052
rect 25740 22040 25746 22092
rect 25792 22080 25820 22120
rect 25869 22117 25881 22151
rect 25915 22148 25927 22151
rect 26421 22151 26479 22157
rect 26421 22148 26433 22151
rect 25915 22120 26433 22148
rect 25915 22117 25927 22120
rect 25869 22111 25927 22117
rect 26421 22117 26433 22120
rect 26467 22117 26479 22151
rect 26421 22111 26479 22117
rect 25792 22052 26188 22080
rect 24912 21984 24992 22012
rect 24912 21972 24918 21984
rect 25590 21972 25596 22024
rect 25648 22012 25654 22024
rect 25777 22015 25835 22021
rect 25777 22012 25789 22015
rect 25648 21984 25789 22012
rect 25648 21972 25654 21984
rect 25777 21981 25789 21984
rect 25823 21981 25835 22015
rect 25777 21975 25835 21981
rect 25866 21972 25872 22024
rect 25924 22012 25930 22024
rect 26160 22021 26188 22052
rect 26053 22015 26111 22021
rect 26053 22012 26065 22015
rect 25924 21984 26065 22012
rect 25924 21972 25930 21984
rect 26053 21981 26065 21984
rect 26099 21981 26111 22015
rect 26053 21975 26111 21981
rect 26145 22015 26203 22021
rect 26145 21981 26157 22015
rect 26191 21981 26203 22015
rect 26145 21975 26203 21981
rect 26234 21972 26240 22024
rect 26292 22012 26298 22024
rect 26421 22015 26479 22021
rect 26421 22012 26433 22015
rect 26292 21984 26433 22012
rect 26292 21972 26298 21984
rect 26421 21981 26433 21984
rect 26467 21981 26479 22015
rect 26421 21975 26479 21981
rect 27522 21972 27528 22024
rect 27580 21972 27586 22024
rect 23891 21916 23980 21944
rect 24044 21916 24532 21944
rect 25317 21947 25375 21953
rect 23891 21913 23903 21916
rect 23845 21907 23903 21913
rect 19426 21876 19432 21888
rect 17236 21848 19432 21876
rect 19426 21836 19432 21848
rect 19484 21836 19490 21888
rect 24044 21885 24072 21916
rect 25317 21913 25329 21947
rect 25363 21944 25375 21947
rect 25958 21944 25964 21956
rect 25363 21916 25964 21944
rect 25363 21913 25375 21916
rect 25317 21907 25375 21913
rect 25958 21904 25964 21916
rect 26016 21904 26022 21956
rect 24044 21879 24113 21885
rect 24044 21848 24067 21879
rect 24055 21845 24067 21848
rect 24101 21845 24113 21879
rect 24055 21839 24113 21845
rect 24213 21879 24271 21885
rect 24213 21845 24225 21879
rect 24259 21876 24271 21879
rect 24578 21876 24584 21888
rect 24259 21848 24584 21876
rect 24259 21845 24271 21848
rect 24213 21839 24271 21845
rect 24578 21836 24584 21848
rect 24636 21836 24642 21888
rect 24762 21836 24768 21888
rect 24820 21876 24826 21888
rect 25041 21879 25099 21885
rect 25041 21876 25053 21879
rect 24820 21848 25053 21876
rect 24820 21836 24826 21848
rect 25041 21845 25053 21848
rect 25087 21845 25099 21879
rect 25041 21839 25099 21845
rect 25130 21836 25136 21888
rect 25188 21876 25194 21888
rect 25517 21879 25575 21885
rect 25517 21876 25529 21879
rect 25188 21848 25529 21876
rect 25188 21836 25194 21848
rect 25517 21845 25529 21848
rect 25563 21845 25575 21879
rect 25517 21839 25575 21845
rect 25682 21836 25688 21888
rect 25740 21836 25746 21888
rect 25866 21836 25872 21888
rect 25924 21876 25930 21888
rect 26237 21879 26295 21885
rect 26237 21876 26249 21879
rect 25924 21848 26249 21876
rect 25924 21836 25930 21848
rect 26237 21845 26249 21848
rect 26283 21845 26295 21879
rect 26237 21839 26295 21845
rect 27706 21836 27712 21888
rect 27764 21836 27770 21888
rect 1104 21786 28152 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 28152 21786
rect 1104 21712 28152 21734
rect 14274 21632 14280 21684
rect 14332 21632 14338 21684
rect 14461 21675 14519 21681
rect 14461 21641 14473 21675
rect 14507 21641 14519 21675
rect 14461 21635 14519 21641
rect 1302 21564 1308 21616
rect 1360 21604 1366 21616
rect 2501 21607 2559 21613
rect 2501 21604 2513 21607
rect 1360 21576 2513 21604
rect 1360 21564 1366 21576
rect 2501 21573 2513 21576
rect 2547 21573 2559 21607
rect 2501 21567 2559 21573
rect 2869 21607 2927 21613
rect 2869 21573 2881 21607
rect 2915 21604 2927 21607
rect 2958 21604 2964 21616
rect 2915 21576 2964 21604
rect 2915 21573 2927 21576
rect 2869 21567 2927 21573
rect 2958 21564 2964 21576
rect 3016 21564 3022 21616
rect 7466 21564 7472 21616
rect 7524 21604 7530 21616
rect 7524 21576 7788 21604
rect 7524 21564 7530 21576
rect 1394 21496 1400 21548
rect 1452 21496 1458 21548
rect 2225 21539 2283 21545
rect 2225 21505 2237 21539
rect 2271 21536 2283 21539
rect 2314 21536 2320 21548
rect 2271 21508 2320 21536
rect 2271 21505 2283 21508
rect 2225 21499 2283 21505
rect 2314 21496 2320 21508
rect 2372 21496 2378 21548
rect 3602 21496 3608 21548
rect 3660 21496 3666 21548
rect 3970 21496 3976 21548
rect 4028 21496 4034 21548
rect 4798 21496 4804 21548
rect 4856 21536 4862 21548
rect 4893 21539 4951 21545
rect 4893 21536 4905 21539
rect 4856 21508 4905 21536
rect 4856 21496 4862 21508
rect 4893 21505 4905 21508
rect 4939 21505 4951 21539
rect 4893 21499 4951 21505
rect 5077 21539 5135 21545
rect 5077 21505 5089 21539
rect 5123 21536 5135 21539
rect 5258 21536 5264 21548
rect 5123 21508 5264 21536
rect 5123 21505 5135 21508
rect 5077 21499 5135 21505
rect 5258 21496 5264 21508
rect 5316 21496 5322 21548
rect 7561 21539 7619 21545
rect 7561 21505 7573 21539
rect 7607 21536 7619 21539
rect 7650 21536 7656 21548
rect 7607 21508 7656 21536
rect 7607 21505 7619 21508
rect 7561 21499 7619 21505
rect 7650 21496 7656 21508
rect 7708 21496 7714 21548
rect 7760 21545 7788 21576
rect 14090 21564 14096 21616
rect 14148 21604 14154 21616
rect 14369 21607 14427 21613
rect 14148 21576 14320 21604
rect 14148 21564 14154 21576
rect 7745 21539 7803 21545
rect 7745 21505 7757 21539
rect 7791 21505 7803 21539
rect 7745 21499 7803 21505
rect 12066 21496 12072 21548
rect 12124 21536 12130 21548
rect 14292 21536 14320 21576
rect 14369 21573 14381 21607
rect 14415 21604 14427 21607
rect 14476 21604 14504 21635
rect 15010 21632 15016 21684
rect 15068 21632 15074 21684
rect 16301 21675 16359 21681
rect 16301 21641 16313 21675
rect 16347 21672 16359 21675
rect 17218 21672 17224 21684
rect 16347 21644 17224 21672
rect 16347 21641 16359 21644
rect 16301 21635 16359 21641
rect 17218 21632 17224 21644
rect 17276 21632 17282 21684
rect 24949 21675 25007 21681
rect 24949 21641 24961 21675
rect 24995 21672 25007 21675
rect 25130 21672 25136 21684
rect 24995 21644 25136 21672
rect 24995 21641 25007 21644
rect 24949 21635 25007 21641
rect 25130 21632 25136 21644
rect 25188 21632 25194 21684
rect 25222 21632 25228 21684
rect 25280 21672 25286 21684
rect 26789 21675 26847 21681
rect 25280 21644 26648 21672
rect 25280 21632 25286 21644
rect 14415 21576 14504 21604
rect 15028 21604 15056 21632
rect 16485 21607 16543 21613
rect 15028 21576 15424 21604
rect 14415 21573 14427 21576
rect 14369 21567 14427 21573
rect 15013 21539 15071 21545
rect 15013 21536 15025 21539
rect 12124 21508 14228 21536
rect 14292 21508 15025 21536
rect 12124 21496 12130 21508
rect 4617 21471 4675 21477
rect 4617 21437 4629 21471
rect 4663 21468 4675 21471
rect 4706 21468 4712 21480
rect 4663 21440 4712 21468
rect 4663 21437 4675 21440
rect 4617 21431 4675 21437
rect 4706 21428 4712 21440
rect 4764 21428 4770 21480
rect 4985 21471 5043 21477
rect 4985 21437 4997 21471
rect 5031 21468 5043 21471
rect 5353 21471 5411 21477
rect 5353 21468 5365 21471
rect 5031 21440 5365 21468
rect 5031 21437 5043 21440
rect 4985 21431 5043 21437
rect 5353 21437 5365 21440
rect 5399 21437 5411 21471
rect 5353 21431 5411 21437
rect 5718 21428 5724 21480
rect 5776 21428 5782 21480
rect 5813 21471 5871 21477
rect 5813 21437 5825 21471
rect 5859 21468 5871 21471
rect 6086 21468 6092 21480
rect 5859 21440 6092 21468
rect 5859 21437 5871 21440
rect 5813 21431 5871 21437
rect 6086 21428 6092 21440
rect 6144 21428 6150 21480
rect 13998 21428 14004 21480
rect 14056 21428 14062 21480
rect 8570 21360 8576 21412
rect 8628 21360 8634 21412
rect 13814 21360 13820 21412
rect 13872 21400 13878 21412
rect 14093 21403 14151 21409
rect 14093 21400 14105 21403
rect 13872 21372 14105 21400
rect 13872 21360 13878 21372
rect 14093 21369 14105 21372
rect 14139 21369 14151 21403
rect 14200 21400 14228 21508
rect 15013 21505 15025 21508
rect 15059 21505 15071 21539
rect 15013 21499 15071 21505
rect 15286 21496 15292 21548
rect 15344 21496 15350 21548
rect 15396 21545 15424 21576
rect 16485 21573 16497 21607
rect 16531 21604 16543 21607
rect 17034 21604 17040 21616
rect 16531 21576 17040 21604
rect 16531 21573 16543 21576
rect 16485 21567 16543 21573
rect 17034 21564 17040 21576
rect 17092 21604 17098 21616
rect 17310 21604 17316 21616
rect 17092 21576 17316 21604
rect 17092 21564 17098 21576
rect 17310 21564 17316 21576
rect 17368 21564 17374 21616
rect 17681 21607 17739 21613
rect 17681 21573 17693 21607
rect 17727 21604 17739 21607
rect 18874 21604 18880 21616
rect 17727 21576 18880 21604
rect 17727 21573 17739 21576
rect 17681 21567 17739 21573
rect 18874 21564 18880 21576
rect 18932 21564 18938 21616
rect 19610 21604 19616 21616
rect 18984 21576 19616 21604
rect 15381 21539 15439 21545
rect 15381 21505 15393 21539
rect 15427 21536 15439 21539
rect 15565 21539 15623 21545
rect 15565 21536 15577 21539
rect 15427 21508 15577 21536
rect 15427 21505 15439 21508
rect 15381 21499 15439 21505
rect 15565 21505 15577 21508
rect 15611 21505 15623 21539
rect 15565 21499 15623 21505
rect 16206 21496 16212 21548
rect 16264 21496 16270 21548
rect 16390 21496 16396 21548
rect 16448 21536 16454 21548
rect 16945 21539 17003 21545
rect 16945 21536 16957 21539
rect 16448 21508 16957 21536
rect 16448 21496 16454 21508
rect 16945 21505 16957 21508
rect 16991 21505 17003 21539
rect 17586 21536 17592 21548
rect 16945 21499 17003 21505
rect 17144 21508 17592 21536
rect 14366 21428 14372 21480
rect 14424 21468 14430 21480
rect 14642 21468 14648 21480
rect 14424 21440 14648 21468
rect 14424 21428 14430 21440
rect 14642 21428 14648 21440
rect 14700 21468 14706 21480
rect 14737 21471 14795 21477
rect 14737 21468 14749 21471
rect 14700 21440 14749 21468
rect 14700 21428 14706 21440
rect 14737 21437 14749 21440
rect 14783 21437 14795 21471
rect 14737 21431 14795 21437
rect 14826 21428 14832 21480
rect 14884 21468 14890 21480
rect 16758 21468 16764 21480
rect 14884 21440 16764 21468
rect 14884 21428 14890 21440
rect 16758 21428 16764 21440
rect 16816 21428 16822 21480
rect 17144 21477 17172 21508
rect 17586 21496 17592 21508
rect 17644 21536 17650 21548
rect 17773 21539 17831 21545
rect 17773 21536 17785 21539
rect 17644 21508 17785 21536
rect 17644 21496 17650 21508
rect 17773 21505 17785 21508
rect 17819 21505 17831 21539
rect 17773 21499 17831 21505
rect 18138 21496 18144 21548
rect 18196 21536 18202 21548
rect 18233 21539 18291 21545
rect 18233 21536 18245 21539
rect 18196 21508 18245 21536
rect 18196 21496 18202 21508
rect 18233 21505 18245 21508
rect 18279 21536 18291 21539
rect 18322 21536 18328 21548
rect 18279 21508 18328 21536
rect 18279 21505 18291 21508
rect 18233 21499 18291 21505
rect 18322 21496 18328 21508
rect 18380 21496 18386 21548
rect 18414 21496 18420 21548
rect 18472 21536 18478 21548
rect 18598 21536 18604 21548
rect 18472 21508 18604 21536
rect 18472 21496 18478 21508
rect 18598 21496 18604 21508
rect 18656 21496 18662 21548
rect 18984 21545 19012 21576
rect 19610 21564 19616 21576
rect 19668 21564 19674 21616
rect 24670 21604 24676 21616
rect 24320 21576 24676 21604
rect 18969 21539 19027 21545
rect 18969 21505 18981 21539
rect 19015 21505 19027 21539
rect 18969 21499 19027 21505
rect 16853 21471 16911 21477
rect 16853 21437 16865 21471
rect 16899 21437 16911 21471
rect 16853 21431 16911 21437
rect 17129 21471 17187 21477
rect 17129 21437 17141 21471
rect 17175 21437 17187 21471
rect 17129 21431 17187 21437
rect 15378 21400 15384 21412
rect 14200 21372 14872 21400
rect 14093 21363 14151 21369
rect 14844 21344 14872 21372
rect 14936 21372 15384 21400
rect 5997 21335 6055 21341
rect 5997 21301 6009 21335
rect 6043 21332 6055 21335
rect 6914 21332 6920 21344
rect 6043 21304 6920 21332
rect 6043 21301 6055 21304
rect 5997 21295 6055 21301
rect 6914 21292 6920 21304
rect 6972 21292 6978 21344
rect 13906 21292 13912 21344
rect 13964 21292 13970 21344
rect 14458 21292 14464 21344
rect 14516 21332 14522 21344
rect 14734 21332 14740 21344
rect 14516 21304 14740 21332
rect 14516 21292 14522 21304
rect 14734 21292 14740 21304
rect 14792 21292 14798 21344
rect 14826 21292 14832 21344
rect 14884 21292 14890 21344
rect 14936 21341 14964 21372
rect 15378 21360 15384 21372
rect 15436 21400 15442 21412
rect 15657 21403 15715 21409
rect 15657 21400 15669 21403
rect 15436 21372 15669 21400
rect 15436 21360 15442 21372
rect 15657 21369 15669 21372
rect 15703 21369 15715 21403
rect 15657 21363 15715 21369
rect 16574 21360 16580 21412
rect 16632 21400 16638 21412
rect 16868 21400 16896 21431
rect 18046 21428 18052 21480
rect 18104 21468 18110 21480
rect 18984 21468 19012 21499
rect 19058 21496 19064 21548
rect 19116 21536 19122 21548
rect 24320 21545 24348 21576
rect 24670 21564 24676 21576
rect 24728 21564 24734 21616
rect 25314 21564 25320 21616
rect 25372 21564 25378 21616
rect 25406 21564 25412 21616
rect 25464 21604 25470 21616
rect 26620 21604 26648 21644
rect 26789 21641 26801 21675
rect 26835 21672 26847 21675
rect 27430 21672 27436 21684
rect 26835 21644 27436 21672
rect 26835 21641 26847 21644
rect 26789 21635 26847 21641
rect 27430 21632 27436 21644
rect 27488 21632 27494 21684
rect 27065 21607 27123 21613
rect 27065 21604 27077 21607
rect 25464 21576 25806 21604
rect 26620 21576 27077 21604
rect 25464 21564 25470 21576
rect 27065 21573 27077 21576
rect 27111 21573 27123 21607
rect 27065 21567 27123 21573
rect 19521 21539 19579 21545
rect 19521 21536 19533 21539
rect 19116 21508 19533 21536
rect 19116 21496 19122 21508
rect 19521 21505 19533 21508
rect 19567 21505 19579 21539
rect 19521 21499 19579 21505
rect 24305 21539 24363 21545
rect 24305 21505 24317 21539
rect 24351 21505 24363 21539
rect 24305 21499 24363 21505
rect 24489 21539 24547 21545
rect 24489 21505 24501 21539
rect 24535 21536 24547 21539
rect 24578 21536 24584 21548
rect 24535 21508 24584 21536
rect 24535 21505 24547 21508
rect 24489 21499 24547 21505
rect 18104 21440 19012 21468
rect 18104 21428 18110 21440
rect 19426 21428 19432 21480
rect 19484 21428 19490 21480
rect 16632 21372 16896 21400
rect 16632 21360 16638 21372
rect 17218 21360 17224 21412
rect 17276 21400 17282 21412
rect 17313 21403 17371 21409
rect 17313 21400 17325 21403
rect 17276 21372 17325 21400
rect 17276 21360 17282 21372
rect 17313 21369 17325 21372
rect 17359 21369 17371 21403
rect 17313 21363 17371 21369
rect 19889 21403 19947 21409
rect 19889 21369 19901 21403
rect 19935 21400 19947 21403
rect 19978 21400 19984 21412
rect 19935 21372 19984 21400
rect 19935 21369 19947 21372
rect 19889 21363 19947 21369
rect 19978 21360 19984 21372
rect 20036 21360 20042 21412
rect 24504 21400 24532 21499
rect 24578 21496 24584 21508
rect 24636 21496 24642 21548
rect 24762 21496 24768 21548
rect 24820 21496 24826 21548
rect 27798 21496 27804 21548
rect 27856 21496 27862 21548
rect 24670 21428 24676 21480
rect 24728 21468 24734 21480
rect 25041 21471 25099 21477
rect 25041 21468 25053 21471
rect 24728 21440 25053 21468
rect 24728 21428 24734 21440
rect 25041 21437 25053 21440
rect 25087 21437 25099 21471
rect 25041 21431 25099 21437
rect 26050 21428 26056 21480
rect 26108 21468 26114 21480
rect 27249 21471 27307 21477
rect 27249 21468 27261 21471
rect 26108 21440 27261 21468
rect 26108 21428 26114 21440
rect 27249 21437 27261 21440
rect 27295 21437 27307 21471
rect 27249 21431 27307 21437
rect 24946 21400 24952 21412
rect 24504 21372 24952 21400
rect 24946 21360 24952 21372
rect 25004 21360 25010 21412
rect 14921 21335 14979 21341
rect 14921 21301 14933 21335
rect 14967 21301 14979 21335
rect 14921 21295 14979 21301
rect 15010 21292 15016 21344
rect 15068 21332 15074 21344
rect 15105 21335 15163 21341
rect 15105 21332 15117 21335
rect 15068 21304 15117 21332
rect 15068 21292 15074 21304
rect 15105 21301 15117 21304
rect 15151 21301 15163 21335
rect 15105 21295 15163 21301
rect 16485 21335 16543 21341
rect 16485 21301 16497 21335
rect 16531 21332 16543 21335
rect 17034 21332 17040 21344
rect 16531 21304 17040 21332
rect 16531 21301 16543 21304
rect 16485 21295 16543 21301
rect 17034 21292 17040 21304
rect 17092 21292 17098 21344
rect 24210 21292 24216 21344
rect 24268 21332 24274 21344
rect 25866 21332 25872 21344
rect 24268 21304 25872 21332
rect 24268 21292 24274 21304
rect 25866 21292 25872 21304
rect 25924 21292 25930 21344
rect 27614 21292 27620 21344
rect 27672 21292 27678 21344
rect 1104 21242 28152 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 28152 21242
rect 1104 21168 28152 21190
rect 12158 21088 12164 21140
rect 12216 21128 12222 21140
rect 12253 21131 12311 21137
rect 12253 21128 12265 21131
rect 12216 21100 12265 21128
rect 12216 21088 12222 21100
rect 12253 21097 12265 21100
rect 12299 21097 12311 21131
rect 12253 21091 12311 21097
rect 14553 21131 14611 21137
rect 14553 21097 14565 21131
rect 14599 21128 14611 21131
rect 15102 21128 15108 21140
rect 14599 21100 15108 21128
rect 14599 21097 14611 21100
rect 14553 21091 14611 21097
rect 15102 21088 15108 21100
rect 15160 21088 15166 21140
rect 15194 21088 15200 21140
rect 15252 21128 15258 21140
rect 15252 21100 16068 21128
rect 15252 21088 15258 21100
rect 12176 21060 12204 21088
rect 11256 21032 12204 21060
rect 14093 21063 14151 21069
rect 2314 20952 2320 21004
rect 2372 20992 2378 21004
rect 2501 20995 2559 21001
rect 2501 20992 2513 20995
rect 2372 20964 2513 20992
rect 2372 20952 2378 20964
rect 2501 20961 2513 20964
rect 2547 20961 2559 20995
rect 2501 20955 2559 20961
rect 2596 20936 2648 20942
rect 4614 20884 4620 20936
rect 4672 20924 4678 20936
rect 4985 20927 5043 20933
rect 4985 20924 4997 20927
rect 4672 20896 4997 20924
rect 4672 20884 4678 20896
rect 4985 20893 4997 20896
rect 5031 20893 5043 20927
rect 4985 20887 5043 20893
rect 5258 20884 5264 20936
rect 5316 20884 5322 20936
rect 5353 20927 5411 20933
rect 5353 20893 5365 20927
rect 5399 20924 5411 20927
rect 5537 20927 5595 20933
rect 5537 20924 5549 20927
rect 5399 20896 5549 20924
rect 5399 20893 5411 20896
rect 5353 20887 5411 20893
rect 5537 20893 5549 20896
rect 5583 20924 5595 20927
rect 5718 20924 5724 20936
rect 5583 20896 5724 20924
rect 5583 20893 5595 20896
rect 5537 20887 5595 20893
rect 5718 20884 5724 20896
rect 5776 20884 5782 20936
rect 6086 20884 6092 20936
rect 6144 20884 6150 20936
rect 7098 20884 7104 20936
rect 7156 20924 7162 20936
rect 7561 20927 7619 20933
rect 7561 20924 7573 20927
rect 7156 20896 7573 20924
rect 7156 20884 7162 20896
rect 7561 20893 7573 20896
rect 7607 20893 7619 20927
rect 7561 20887 7619 20893
rect 2596 20878 2648 20884
rect 1949 20859 2007 20865
rect 1949 20825 1961 20859
rect 1995 20825 2007 20859
rect 1949 20819 2007 20825
rect 1964 20788 1992 20819
rect 6546 20816 6552 20868
rect 6604 20816 6610 20868
rect 7668 20856 7696 20910
rect 11146 20884 11152 20936
rect 11204 20884 11210 20936
rect 11256 20933 11284 21032
rect 14093 21029 14105 21063
rect 14139 21060 14151 21063
rect 15838 21060 15844 21072
rect 14139 21032 14872 21060
rect 14139 21029 14151 21032
rect 14093 21023 14151 21029
rect 11514 20952 11520 21004
rect 11572 20952 11578 21004
rect 12066 20952 12072 21004
rect 12124 20952 12130 21004
rect 12802 20952 12808 21004
rect 12860 20992 12866 21004
rect 14461 20995 14519 21001
rect 14461 20992 14473 20995
rect 12860 20964 14473 20992
rect 12860 20952 12866 20964
rect 14461 20961 14473 20964
rect 14507 20992 14519 20995
rect 14734 20992 14740 21004
rect 14507 20964 14740 20992
rect 14507 20961 14519 20964
rect 14461 20955 14519 20961
rect 14734 20952 14740 20964
rect 14792 20952 14798 21004
rect 14844 21001 14872 21032
rect 15028 21032 15844 21060
rect 15028 21001 15056 21032
rect 15838 21020 15844 21032
rect 15896 21020 15902 21072
rect 14829 20995 14887 21001
rect 14829 20961 14841 20995
rect 14875 20961 14887 20995
rect 14829 20955 14887 20961
rect 15013 20995 15071 21001
rect 15013 20961 15025 20995
rect 15059 20961 15071 20995
rect 15013 20955 15071 20961
rect 15105 20995 15163 21001
rect 15105 20961 15117 20995
rect 15151 20992 15163 20995
rect 15151 20964 15884 20992
rect 15151 20961 15163 20964
rect 15105 20955 15163 20961
rect 11241 20927 11299 20933
rect 11241 20893 11253 20927
rect 11287 20924 11299 20927
rect 11330 20924 11336 20936
rect 11287 20896 11336 20924
rect 11287 20893 11299 20896
rect 11241 20887 11299 20893
rect 11330 20884 11336 20896
rect 11388 20884 11394 20936
rect 11606 20884 11612 20936
rect 11664 20884 11670 20936
rect 12345 20927 12403 20933
rect 12345 20893 12357 20927
rect 12391 20924 12403 20927
rect 12526 20924 12532 20936
rect 12391 20896 12532 20924
rect 12391 20893 12403 20896
rect 12345 20887 12403 20893
rect 12526 20884 12532 20896
rect 12584 20884 12590 20936
rect 13170 20884 13176 20936
rect 13228 20924 13234 20936
rect 13449 20927 13507 20933
rect 13449 20924 13461 20927
rect 13228 20896 13461 20924
rect 13228 20884 13234 20896
rect 13449 20893 13461 20896
rect 13495 20924 13507 20927
rect 13538 20924 13544 20936
rect 13495 20896 13544 20924
rect 13495 20893 13507 20896
rect 13449 20887 13507 20893
rect 13538 20884 13544 20896
rect 13596 20884 13602 20936
rect 13633 20927 13691 20933
rect 13633 20893 13645 20927
rect 13679 20924 13691 20927
rect 14090 20924 14096 20936
rect 13679 20896 14096 20924
rect 13679 20893 13691 20896
rect 13633 20887 13691 20893
rect 14090 20884 14096 20896
rect 14148 20884 14154 20936
rect 14277 20927 14335 20933
rect 14277 20893 14289 20927
rect 14323 20924 14335 20927
rect 14366 20924 14372 20936
rect 14323 20896 14372 20924
rect 14323 20893 14335 20896
rect 14277 20887 14335 20893
rect 14366 20884 14372 20896
rect 14424 20884 14430 20936
rect 14550 20884 14556 20936
rect 14608 20884 14614 20936
rect 14918 20884 14924 20936
rect 14976 20884 14982 20936
rect 15856 20933 15884 20964
rect 16040 20933 16068 21100
rect 17218 21088 17224 21140
rect 17276 21088 17282 21140
rect 18322 21088 18328 21140
rect 18380 21128 18386 21140
rect 18782 21128 18788 21140
rect 18380 21100 18788 21128
rect 18380 21088 18386 21100
rect 18782 21088 18788 21100
rect 18840 21088 18846 21140
rect 19058 21088 19064 21140
rect 19116 21128 19122 21140
rect 21450 21128 21456 21140
rect 19116 21100 21456 21128
rect 19116 21088 19122 21100
rect 21450 21088 21456 21100
rect 21508 21088 21514 21140
rect 22646 21128 22652 21140
rect 21559 21100 22652 21128
rect 16485 21063 16543 21069
rect 16485 21029 16497 21063
rect 16531 21060 16543 21063
rect 16574 21060 16580 21072
rect 16531 21032 16580 21060
rect 16531 21029 16543 21032
rect 16485 21023 16543 21029
rect 16574 21020 16580 21032
rect 16632 21020 16638 21072
rect 16758 20952 16764 21004
rect 16816 20992 16822 21004
rect 16945 20995 17003 21001
rect 16945 20992 16957 20995
rect 16816 20964 16957 20992
rect 16816 20952 16822 20964
rect 16945 20961 16957 20964
rect 16991 20961 17003 20995
rect 16945 20955 17003 20961
rect 17037 20995 17095 21001
rect 17037 20961 17049 20995
rect 17083 20992 17095 20995
rect 17126 20992 17132 21004
rect 17083 20964 17132 20992
rect 17083 20961 17095 20964
rect 17037 20955 17095 20961
rect 17126 20952 17132 20964
rect 17184 20952 17190 21004
rect 17236 20992 17264 21088
rect 17313 21063 17371 21069
rect 17313 21029 17325 21063
rect 17359 21060 17371 21063
rect 17359 21032 19840 21060
rect 17359 21029 17371 21032
rect 17313 21023 17371 21029
rect 17497 20995 17555 21001
rect 17497 20992 17509 20995
rect 17236 20964 17509 20992
rect 17497 20961 17509 20964
rect 17543 20961 17555 20995
rect 17497 20955 17555 20961
rect 17586 20952 17592 21004
rect 17644 20952 17650 21004
rect 17865 20995 17923 21001
rect 17865 20961 17877 20995
rect 17911 20992 17923 20995
rect 18414 20992 18420 21004
rect 17911 20964 18420 20992
rect 17911 20961 17923 20964
rect 17865 20955 17923 20961
rect 18414 20952 18420 20964
rect 18472 20952 18478 21004
rect 19613 20995 19671 21001
rect 19613 20992 19625 20995
rect 18524 20964 19625 20992
rect 15657 20927 15715 20933
rect 15657 20924 15669 20927
rect 15580 20896 15669 20924
rect 7576 20828 7696 20856
rect 2038 20788 2044 20800
rect 1964 20760 2044 20788
rect 2038 20748 2044 20760
rect 2096 20748 2102 20800
rect 6270 20748 6276 20800
rect 6328 20788 6334 20800
rect 7576 20788 7604 20828
rect 8294 20816 8300 20868
rect 8352 20816 8358 20868
rect 11882 20816 11888 20868
rect 11940 20816 11946 20868
rect 14734 20816 14740 20868
rect 14792 20856 14798 20868
rect 15580 20856 15608 20896
rect 15657 20893 15669 20896
rect 15703 20893 15715 20927
rect 15657 20887 15715 20893
rect 15841 20927 15899 20933
rect 15841 20893 15853 20927
rect 15887 20893 15899 20927
rect 15841 20887 15899 20893
rect 16025 20927 16083 20933
rect 16025 20893 16037 20927
rect 16071 20924 16083 20927
rect 16206 20924 16212 20936
rect 16071 20896 16212 20924
rect 16071 20893 16083 20896
rect 16025 20887 16083 20893
rect 16206 20884 16212 20896
rect 16264 20884 16270 20936
rect 16301 20927 16359 20933
rect 16301 20893 16313 20927
rect 16347 20924 16359 20927
rect 17770 20924 17776 20936
rect 16347 20896 17776 20924
rect 16347 20893 16359 20896
rect 16301 20887 16359 20893
rect 17770 20884 17776 20896
rect 17828 20884 17834 20936
rect 17957 20927 18015 20933
rect 17957 20893 17969 20927
rect 18003 20924 18015 20927
rect 18046 20924 18052 20936
rect 18003 20896 18052 20924
rect 18003 20893 18015 20896
rect 17957 20887 18015 20893
rect 18046 20884 18052 20896
rect 18104 20884 18110 20936
rect 18524 20933 18552 20964
rect 19613 20961 19625 20964
rect 19659 20961 19671 20995
rect 19812 20992 19840 21032
rect 19886 21020 19892 21072
rect 19944 21020 19950 21072
rect 20438 21020 20444 21072
rect 20496 21060 20502 21072
rect 21559 21060 21587 21100
rect 22646 21088 22652 21100
rect 22704 21088 22710 21140
rect 20496 21032 21587 21060
rect 20496 21020 20502 21032
rect 22186 21020 22192 21072
rect 22244 21020 22250 21072
rect 21542 20992 21548 21004
rect 19812 20964 20300 20992
rect 19613 20955 19671 20961
rect 18233 20927 18291 20933
rect 18233 20893 18245 20927
rect 18279 20893 18291 20927
rect 18233 20887 18291 20893
rect 18509 20927 18567 20933
rect 18509 20893 18521 20927
rect 18555 20893 18567 20927
rect 18509 20887 18567 20893
rect 14792 20828 15608 20856
rect 14792 20816 14798 20828
rect 16482 20816 16488 20868
rect 16540 20816 16546 20868
rect 18138 20856 18144 20868
rect 17788 20828 18144 20856
rect 6328 20760 7604 20788
rect 6328 20748 6334 20760
rect 13538 20748 13544 20800
rect 13596 20748 13602 20800
rect 14274 20748 14280 20800
rect 14332 20788 14338 20800
rect 14458 20788 14464 20800
rect 14332 20760 14464 20788
rect 14332 20748 14338 20760
rect 14458 20748 14464 20760
rect 14516 20788 14522 20800
rect 14645 20791 14703 20797
rect 14645 20788 14657 20791
rect 14516 20760 14657 20788
rect 14516 20748 14522 20760
rect 14645 20757 14657 20760
rect 14691 20757 14703 20791
rect 14645 20751 14703 20757
rect 15194 20748 15200 20800
rect 15252 20788 15258 20800
rect 15381 20791 15439 20797
rect 15381 20788 15393 20791
rect 15252 20760 15393 20788
rect 15252 20748 15258 20760
rect 15381 20757 15393 20760
rect 15427 20757 15439 20791
rect 15381 20751 15439 20757
rect 15470 20748 15476 20800
rect 15528 20788 15534 20800
rect 17788 20797 17816 20828
rect 18138 20816 18144 20828
rect 18196 20816 18202 20868
rect 18248 20856 18276 20887
rect 18782 20884 18788 20936
rect 18840 20884 18846 20936
rect 19058 20924 19064 20936
rect 18892 20896 19064 20924
rect 18601 20859 18659 20865
rect 18601 20856 18613 20859
rect 18248 20828 18613 20856
rect 18601 20825 18613 20828
rect 18647 20825 18659 20859
rect 18601 20819 18659 20825
rect 18690 20816 18696 20868
rect 18748 20856 18754 20868
rect 18892 20856 18920 20896
rect 19058 20884 19064 20896
rect 19116 20884 19122 20936
rect 19150 20884 19156 20936
rect 19208 20884 19214 20936
rect 19521 20927 19579 20933
rect 19521 20893 19533 20927
rect 19567 20924 19579 20927
rect 19702 20924 19708 20936
rect 19567 20896 19708 20924
rect 19567 20893 19579 20896
rect 19521 20887 19579 20893
rect 19702 20884 19708 20896
rect 19760 20884 19766 20936
rect 19797 20927 19855 20933
rect 19797 20893 19809 20927
rect 19843 20924 19855 20927
rect 19886 20924 19892 20936
rect 19843 20896 19892 20924
rect 19843 20893 19855 20896
rect 19797 20887 19855 20893
rect 19886 20884 19892 20896
rect 19944 20884 19950 20936
rect 19978 20884 19984 20936
rect 20036 20884 20042 20936
rect 20070 20884 20076 20936
rect 20128 20884 20134 20936
rect 20272 20933 20300 20964
rect 20732 20964 21548 20992
rect 20257 20927 20315 20933
rect 20257 20893 20269 20927
rect 20303 20893 20315 20927
rect 20257 20887 20315 20893
rect 18748 20828 18920 20856
rect 18969 20859 19027 20865
rect 18748 20816 18754 20828
rect 18969 20825 18981 20859
rect 19015 20856 19027 20859
rect 19168 20856 19196 20884
rect 19015 20828 19196 20856
rect 19260 20828 19932 20856
rect 19015 20825 19027 20828
rect 18969 20819 19027 20825
rect 16209 20791 16267 20797
rect 16209 20788 16221 20791
rect 15528 20760 16221 20788
rect 15528 20748 15534 20760
rect 16209 20757 16221 20760
rect 16255 20757 16267 20791
rect 16209 20751 16267 20757
rect 17773 20791 17831 20797
rect 17773 20757 17785 20791
rect 17819 20757 17831 20791
rect 17773 20751 17831 20757
rect 18049 20791 18107 20797
rect 18049 20757 18061 20791
rect 18095 20788 18107 20791
rect 18322 20788 18328 20800
rect 18095 20760 18328 20788
rect 18095 20757 18107 20760
rect 18049 20751 18107 20757
rect 18322 20748 18328 20760
rect 18380 20748 18386 20800
rect 18414 20748 18420 20800
rect 18472 20748 18478 20800
rect 18782 20748 18788 20800
rect 18840 20788 18846 20800
rect 19260 20788 19288 20828
rect 18840 20760 19288 20788
rect 19337 20791 19395 20797
rect 18840 20748 18846 20760
rect 19337 20757 19349 20791
rect 19383 20788 19395 20791
rect 19794 20788 19800 20800
rect 19383 20760 19800 20788
rect 19383 20757 19395 20760
rect 19337 20751 19395 20757
rect 19794 20748 19800 20760
rect 19852 20748 19858 20800
rect 19904 20788 19932 20828
rect 20732 20788 20760 20964
rect 21542 20952 21548 20964
rect 21600 20952 21606 21004
rect 22204 20992 22232 21020
rect 22557 20995 22615 21001
rect 22557 20992 22569 20995
rect 21744 20964 22569 20992
rect 21450 20884 21456 20936
rect 21508 20924 21514 20936
rect 21744 20933 21772 20964
rect 22557 20961 22569 20964
rect 22603 20961 22615 20995
rect 22557 20955 22615 20961
rect 24949 20995 25007 21001
rect 24949 20961 24961 20995
rect 24995 20992 25007 20995
rect 25038 20992 25044 21004
rect 24995 20964 25044 20992
rect 24995 20961 25007 20964
rect 24949 20955 25007 20961
rect 25038 20952 25044 20964
rect 25096 20952 25102 21004
rect 21637 20927 21695 20933
rect 21637 20924 21649 20927
rect 21508 20896 21649 20924
rect 21508 20884 21514 20896
rect 21637 20893 21649 20896
rect 21683 20893 21695 20927
rect 21637 20887 21695 20893
rect 21729 20927 21787 20933
rect 21729 20893 21741 20927
rect 21775 20893 21787 20927
rect 21729 20887 21787 20893
rect 21818 20884 21824 20936
rect 21876 20924 21882 20936
rect 21913 20927 21971 20933
rect 21913 20924 21925 20927
rect 21876 20896 21925 20924
rect 21876 20884 21882 20896
rect 21913 20893 21925 20896
rect 21959 20893 21971 20927
rect 21913 20887 21971 20893
rect 22097 20927 22155 20933
rect 22097 20893 22109 20927
rect 22143 20924 22155 20927
rect 22189 20927 22247 20933
rect 22189 20924 22201 20927
rect 22143 20896 22201 20924
rect 22143 20893 22155 20896
rect 22097 20887 22155 20893
rect 22189 20893 22201 20896
rect 22235 20893 22247 20927
rect 22189 20887 22247 20893
rect 19904 20760 20760 20788
rect 21468 20788 21496 20884
rect 21542 20816 21548 20868
rect 21600 20856 21606 20868
rect 22112 20856 22140 20887
rect 22370 20884 22376 20936
rect 22428 20884 22434 20936
rect 22462 20884 22468 20936
rect 22520 20924 22526 20936
rect 22649 20927 22707 20933
rect 22649 20924 22661 20927
rect 22520 20896 22661 20924
rect 22520 20884 22526 20896
rect 22649 20893 22661 20896
rect 22695 20924 22707 20927
rect 23566 20924 23572 20936
rect 22695 20896 23572 20924
rect 22695 20893 22707 20896
rect 22649 20887 22707 20893
rect 23566 20884 23572 20896
rect 23624 20884 23630 20936
rect 24670 20884 24676 20936
rect 24728 20884 24734 20936
rect 21600 20828 22140 20856
rect 21600 20816 21606 20828
rect 24026 20816 24032 20868
rect 24084 20856 24090 20868
rect 25406 20856 25412 20868
rect 24084 20828 25412 20856
rect 24084 20816 24090 20828
rect 25406 20816 25412 20828
rect 25464 20816 25470 20868
rect 21910 20788 21916 20800
rect 21468 20760 21916 20788
rect 21910 20748 21916 20760
rect 21968 20748 21974 20800
rect 22094 20748 22100 20800
rect 22152 20788 22158 20800
rect 22281 20791 22339 20797
rect 22281 20788 22293 20791
rect 22152 20760 22293 20788
rect 22152 20748 22158 20760
rect 22281 20757 22293 20760
rect 22327 20757 22339 20791
rect 22281 20751 22339 20757
rect 26418 20748 26424 20800
rect 26476 20748 26482 20800
rect 1104 20698 28152 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 28152 20698
rect 1104 20624 28152 20646
rect 10781 20587 10839 20593
rect 10781 20553 10793 20587
rect 10827 20584 10839 20587
rect 11606 20584 11612 20596
rect 10827 20556 11612 20584
rect 10827 20553 10839 20556
rect 10781 20547 10839 20553
rect 11606 20544 11612 20556
rect 11664 20544 11670 20596
rect 13081 20587 13139 20593
rect 13081 20553 13093 20587
rect 13127 20584 13139 20587
rect 13814 20584 13820 20596
rect 13127 20556 13820 20584
rect 13127 20553 13139 20556
rect 13081 20547 13139 20553
rect 13814 20544 13820 20556
rect 13872 20584 13878 20596
rect 14829 20587 14887 20593
rect 13872 20556 14780 20584
rect 13872 20544 13878 20556
rect 2792 20488 3556 20516
rect 2792 20460 2820 20488
rect 2038 20408 2044 20460
rect 2096 20408 2102 20460
rect 2222 20408 2228 20460
rect 2280 20408 2286 20460
rect 2774 20408 2780 20460
rect 2832 20408 2838 20460
rect 3528 20457 3556 20488
rect 11146 20476 11152 20528
rect 11204 20516 11210 20528
rect 11204 20488 11468 20516
rect 11204 20476 11210 20488
rect 3513 20451 3571 20457
rect 3513 20417 3525 20451
rect 3559 20417 3571 20451
rect 3513 20411 3571 20417
rect 3697 20451 3755 20457
rect 3697 20417 3709 20451
rect 3743 20417 3755 20451
rect 3697 20411 3755 20417
rect 2133 20383 2191 20389
rect 2133 20349 2145 20383
rect 2179 20380 2191 20383
rect 2593 20383 2651 20389
rect 2593 20380 2605 20383
rect 2179 20352 2605 20380
rect 2179 20349 2191 20352
rect 2133 20343 2191 20349
rect 2593 20349 2605 20352
rect 2639 20380 2651 20383
rect 2639 20352 2774 20380
rect 2639 20349 2651 20352
rect 2593 20343 2651 20349
rect 2746 20312 2774 20352
rect 3418 20340 3424 20392
rect 3476 20340 3482 20392
rect 3712 20312 3740 20411
rect 6270 20408 6276 20460
rect 6328 20448 6334 20460
rect 6733 20451 6791 20457
rect 6733 20448 6745 20451
rect 6328 20420 6745 20448
rect 6328 20408 6334 20420
rect 6733 20417 6745 20420
rect 6779 20417 6791 20451
rect 6733 20411 6791 20417
rect 6914 20408 6920 20460
rect 6972 20408 6978 20460
rect 7926 20408 7932 20460
rect 7984 20408 7990 20460
rect 8205 20451 8263 20457
rect 8205 20417 8217 20451
rect 8251 20448 8263 20451
rect 8294 20448 8300 20460
rect 8251 20420 8300 20448
rect 8251 20417 8263 20420
rect 8205 20411 8263 20417
rect 8294 20408 8300 20420
rect 8352 20408 8358 20460
rect 10965 20451 11023 20457
rect 10965 20417 10977 20451
rect 11011 20417 11023 20451
rect 10965 20411 11023 20417
rect 6825 20383 6883 20389
rect 6825 20349 6837 20383
rect 6871 20380 6883 20383
rect 7193 20383 7251 20389
rect 7193 20380 7205 20383
rect 6871 20352 7205 20380
rect 6871 20349 6883 20352
rect 6825 20343 6883 20349
rect 7193 20349 7205 20352
rect 7239 20349 7251 20383
rect 10980 20380 11008 20411
rect 11054 20408 11060 20460
rect 11112 20408 11118 20460
rect 11238 20408 11244 20460
rect 11296 20408 11302 20460
rect 11330 20408 11336 20460
rect 11388 20408 11394 20460
rect 11440 20448 11468 20488
rect 11514 20476 11520 20528
rect 11572 20476 11578 20528
rect 12250 20516 12256 20528
rect 11900 20488 12256 20516
rect 11609 20451 11667 20457
rect 11609 20448 11621 20451
rect 11440 20420 11621 20448
rect 11609 20417 11621 20420
rect 11655 20448 11667 20451
rect 11790 20448 11796 20460
rect 11655 20420 11796 20448
rect 11655 20417 11667 20420
rect 11609 20411 11667 20417
rect 11790 20408 11796 20420
rect 11848 20408 11854 20460
rect 11900 20457 11928 20488
rect 12250 20476 12256 20488
rect 12308 20476 12314 20528
rect 13449 20519 13507 20525
rect 13449 20485 13461 20519
rect 13495 20516 13507 20519
rect 13538 20516 13544 20528
rect 13495 20488 13544 20516
rect 13495 20485 13507 20488
rect 13449 20479 13507 20485
rect 13538 20476 13544 20488
rect 13596 20476 13602 20528
rect 14752 20516 14780 20556
rect 14829 20553 14841 20587
rect 14875 20584 14887 20587
rect 14918 20584 14924 20596
rect 14875 20556 14924 20584
rect 14875 20553 14887 20556
rect 14829 20547 14887 20553
rect 14918 20544 14924 20556
rect 14976 20544 14982 20596
rect 15102 20544 15108 20596
rect 15160 20584 15166 20596
rect 15657 20587 15715 20593
rect 15657 20584 15669 20587
rect 15160 20556 15669 20584
rect 15160 20544 15166 20556
rect 15657 20553 15669 20556
rect 15703 20553 15715 20587
rect 15657 20547 15715 20553
rect 16942 20544 16948 20596
rect 17000 20584 17006 20596
rect 17000 20556 17540 20584
rect 17000 20544 17006 20556
rect 16574 20516 16580 20528
rect 13924 20488 14504 20516
rect 14752 20488 16580 20516
rect 11885 20451 11943 20457
rect 11885 20417 11897 20451
rect 11931 20417 11943 20451
rect 11885 20411 11943 20417
rect 12069 20451 12127 20457
rect 12069 20417 12081 20451
rect 12115 20417 12127 20451
rect 12069 20411 12127 20417
rect 12084 20380 12112 20411
rect 12342 20408 12348 20460
rect 12400 20408 12406 20460
rect 12434 20408 12440 20460
rect 12492 20408 12498 20460
rect 13262 20408 13268 20460
rect 13320 20448 13326 20460
rect 13725 20451 13783 20457
rect 13725 20448 13737 20451
rect 13320 20420 13737 20448
rect 13320 20408 13326 20420
rect 13725 20417 13737 20420
rect 13771 20417 13783 20451
rect 13725 20411 13783 20417
rect 12618 20380 12624 20392
rect 10980 20352 12624 20380
rect 7193 20343 7251 20349
rect 12618 20340 12624 20352
rect 12676 20340 12682 20392
rect 13740 20380 13768 20411
rect 13814 20408 13820 20460
rect 13872 20448 13878 20460
rect 13924 20457 13952 20488
rect 14476 20457 14504 20488
rect 16574 20476 16580 20488
rect 16632 20516 16638 20528
rect 16632 20488 16988 20516
rect 16632 20476 16638 20488
rect 13909 20451 13967 20457
rect 13909 20448 13921 20451
rect 13872 20420 13921 20448
rect 13872 20408 13878 20420
rect 13909 20417 13921 20420
rect 13955 20417 13967 20451
rect 13909 20411 13967 20417
rect 14001 20451 14059 20457
rect 14001 20417 14013 20451
rect 14047 20417 14059 20451
rect 14001 20411 14059 20417
rect 14277 20451 14335 20457
rect 14277 20417 14289 20451
rect 14323 20417 14335 20451
rect 14277 20411 14335 20417
rect 14461 20451 14519 20457
rect 14461 20417 14473 20451
rect 14507 20417 14519 20451
rect 14461 20411 14519 20417
rect 14016 20380 14044 20411
rect 13740 20352 14044 20380
rect 14292 20380 14320 20411
rect 15010 20408 15016 20460
rect 15068 20408 15074 20460
rect 15105 20451 15163 20457
rect 15105 20417 15117 20451
rect 15151 20448 15163 20451
rect 15194 20448 15200 20460
rect 15151 20420 15200 20448
rect 15151 20417 15163 20420
rect 15105 20411 15163 20417
rect 15194 20408 15200 20420
rect 15252 20408 15258 20460
rect 15286 20408 15292 20460
rect 15344 20408 15350 20460
rect 15378 20408 15384 20460
rect 15436 20408 15442 20460
rect 15470 20408 15476 20460
rect 15528 20408 15534 20460
rect 16669 20451 16727 20457
rect 16669 20417 16681 20451
rect 16715 20448 16727 20451
rect 16758 20448 16764 20460
rect 16715 20420 16764 20448
rect 16715 20417 16727 20420
rect 16669 20411 16727 20417
rect 16758 20408 16764 20420
rect 16816 20408 16822 20460
rect 16960 20457 16988 20488
rect 17034 20476 17040 20528
rect 17092 20516 17098 20528
rect 17512 20525 17540 20556
rect 18414 20544 18420 20596
rect 18472 20584 18478 20596
rect 18785 20587 18843 20593
rect 18785 20584 18797 20587
rect 18472 20556 18797 20584
rect 18472 20544 18478 20556
rect 18785 20553 18797 20556
rect 18831 20553 18843 20587
rect 18785 20547 18843 20553
rect 18874 20544 18880 20596
rect 18932 20584 18938 20596
rect 20901 20587 20959 20593
rect 18932 20556 19932 20584
rect 18932 20544 18938 20556
rect 17313 20519 17371 20525
rect 17313 20516 17325 20519
rect 17092 20488 17325 20516
rect 17092 20476 17098 20488
rect 17313 20485 17325 20488
rect 17359 20485 17371 20519
rect 17313 20479 17371 20485
rect 17497 20519 17555 20525
rect 17497 20485 17509 20519
rect 17543 20485 17555 20519
rect 19794 20516 19800 20528
rect 17497 20479 17555 20485
rect 17696 20488 19104 20516
rect 16945 20451 17003 20457
rect 16945 20417 16957 20451
rect 16991 20417 17003 20451
rect 16945 20411 17003 20417
rect 14550 20380 14556 20392
rect 14292 20352 14556 20380
rect 2746 20284 3740 20312
rect 7653 20315 7711 20321
rect 7653 20281 7665 20315
rect 7699 20312 7711 20315
rect 8386 20312 8392 20324
rect 7699 20284 8392 20312
rect 7699 20281 7711 20284
rect 7653 20275 7711 20281
rect 8386 20272 8392 20284
rect 8444 20272 8450 20324
rect 11238 20272 11244 20324
rect 11296 20312 11302 20324
rect 12158 20312 12164 20324
rect 11296 20284 12164 20312
rect 11296 20272 11302 20284
rect 12158 20272 12164 20284
rect 12216 20312 12222 20324
rect 13722 20312 13728 20324
rect 12216 20284 13728 20312
rect 12216 20272 12222 20284
rect 13722 20272 13728 20284
rect 13780 20272 13786 20324
rect 3142 20204 3148 20256
rect 3200 20244 3206 20256
rect 3513 20247 3571 20253
rect 3513 20244 3525 20247
rect 3200 20216 3525 20244
rect 3200 20204 3206 20216
rect 3513 20213 3525 20216
rect 3559 20213 3571 20247
rect 3513 20207 3571 20213
rect 11054 20204 11060 20256
rect 11112 20244 11118 20256
rect 12250 20244 12256 20256
rect 11112 20216 12256 20244
rect 11112 20204 11118 20216
rect 12250 20204 12256 20216
rect 12308 20204 12314 20256
rect 13538 20204 13544 20256
rect 13596 20204 13602 20256
rect 13909 20247 13967 20253
rect 13909 20213 13921 20247
rect 13955 20244 13967 20247
rect 14292 20244 14320 20352
rect 14550 20340 14556 20352
rect 14608 20340 14614 20392
rect 14645 20383 14703 20389
rect 14645 20349 14657 20383
rect 14691 20380 14703 20383
rect 14734 20380 14740 20392
rect 14691 20352 14740 20380
rect 14691 20349 14703 20352
rect 14645 20343 14703 20349
rect 14734 20340 14740 20352
rect 14792 20340 14798 20392
rect 16482 20340 16488 20392
rect 16540 20380 16546 20392
rect 17696 20380 17724 20488
rect 17954 20408 17960 20460
rect 18012 20408 18018 20460
rect 18049 20451 18107 20457
rect 18049 20417 18061 20451
rect 18095 20448 18107 20451
rect 18598 20448 18604 20460
rect 18095 20420 18604 20448
rect 18095 20417 18107 20420
rect 18049 20411 18107 20417
rect 18598 20408 18604 20420
rect 18656 20408 18662 20460
rect 18966 20408 18972 20460
rect 19024 20408 19030 20460
rect 19076 20457 19104 20488
rect 19260 20488 19800 20516
rect 19260 20460 19288 20488
rect 19794 20476 19800 20488
rect 19852 20476 19858 20528
rect 19061 20451 19119 20457
rect 19061 20417 19073 20451
rect 19107 20417 19119 20451
rect 19061 20411 19119 20417
rect 16540 20352 17724 20380
rect 17773 20383 17831 20389
rect 16540 20340 16546 20352
rect 17773 20349 17785 20383
rect 17819 20349 17831 20383
rect 19076 20380 19104 20411
rect 19242 20408 19248 20460
rect 19300 20408 19306 20460
rect 19334 20408 19340 20460
rect 19392 20408 19398 20460
rect 19521 20451 19579 20457
rect 19521 20417 19533 20451
rect 19567 20448 19579 20451
rect 19904 20448 19932 20556
rect 20901 20553 20913 20587
rect 20947 20584 20959 20587
rect 22370 20584 22376 20596
rect 20947 20556 22376 20584
rect 20947 20553 20959 20556
rect 20901 20547 20959 20553
rect 22370 20544 22376 20556
rect 22428 20544 22434 20596
rect 23566 20544 23572 20596
rect 23624 20544 23630 20596
rect 20070 20476 20076 20528
rect 20128 20516 20134 20528
rect 20530 20516 20536 20528
rect 20128 20488 20536 20516
rect 20128 20476 20134 20488
rect 20530 20476 20536 20488
rect 20588 20476 20594 20528
rect 20749 20519 20807 20525
rect 20749 20485 20761 20519
rect 20795 20516 20807 20519
rect 20795 20488 21220 20516
rect 20795 20485 20807 20488
rect 20749 20479 20807 20485
rect 21192 20460 21220 20488
rect 22094 20476 22100 20528
rect 22152 20476 22158 20528
rect 22554 20476 22560 20528
rect 22612 20476 22618 20528
rect 25222 20476 25228 20528
rect 25280 20516 25286 20528
rect 25501 20519 25559 20525
rect 25501 20516 25513 20519
rect 25280 20488 25513 20516
rect 25280 20476 25286 20488
rect 25501 20485 25513 20488
rect 25547 20485 25559 20519
rect 25501 20479 25559 20485
rect 25685 20519 25743 20525
rect 25685 20485 25697 20519
rect 25731 20516 25743 20519
rect 26418 20516 26424 20528
rect 25731 20488 26424 20516
rect 25731 20485 25743 20488
rect 25685 20479 25743 20485
rect 26418 20476 26424 20488
rect 26476 20476 26482 20528
rect 19567 20420 19932 20448
rect 19567 20417 19579 20420
rect 19521 20411 19579 20417
rect 21174 20408 21180 20460
rect 21232 20408 21238 20460
rect 21269 20451 21327 20457
rect 21269 20417 21281 20451
rect 21315 20417 21327 20451
rect 21269 20411 21327 20417
rect 20990 20380 20996 20392
rect 19076 20352 20996 20380
rect 17773 20343 17831 20349
rect 17221 20315 17279 20321
rect 17221 20281 17233 20315
rect 17267 20312 17279 20315
rect 17788 20312 17816 20343
rect 20990 20340 20996 20352
rect 21048 20340 21054 20392
rect 21284 20380 21312 20411
rect 21358 20408 21364 20460
rect 21416 20408 21422 20460
rect 21542 20408 21548 20460
rect 21600 20408 21606 20460
rect 21637 20451 21695 20457
rect 21637 20417 21649 20451
rect 21683 20417 21695 20451
rect 21637 20411 21695 20417
rect 21450 20380 21456 20392
rect 21284 20352 21456 20380
rect 17267 20284 17816 20312
rect 18049 20315 18107 20321
rect 17267 20281 17279 20284
rect 17221 20275 17279 20281
rect 18049 20281 18061 20315
rect 18095 20312 18107 20315
rect 19702 20312 19708 20324
rect 18095 20284 19708 20312
rect 18095 20281 18107 20284
rect 18049 20275 18107 20281
rect 19702 20272 19708 20284
rect 19760 20272 19766 20324
rect 21284 20312 21312 20352
rect 21450 20340 21456 20352
rect 21508 20340 21514 20392
rect 21652 20380 21680 20411
rect 21560 20352 21680 20380
rect 20732 20284 21312 20312
rect 13955 20216 14320 20244
rect 13955 20213 13967 20216
rect 13909 20207 13967 20213
rect 16390 20204 16396 20256
rect 16448 20244 16454 20256
rect 16761 20247 16819 20253
rect 16761 20244 16773 20247
rect 16448 20216 16773 20244
rect 16448 20204 16454 20216
rect 16761 20213 16773 20216
rect 16807 20213 16819 20247
rect 16761 20207 16819 20213
rect 17494 20204 17500 20256
rect 17552 20244 17558 20256
rect 17681 20247 17739 20253
rect 17681 20244 17693 20247
rect 17552 20216 17693 20244
rect 17552 20204 17558 20216
rect 17681 20213 17693 20216
rect 17727 20213 17739 20247
rect 17681 20207 17739 20213
rect 18966 20204 18972 20256
rect 19024 20244 19030 20256
rect 19613 20247 19671 20253
rect 19613 20244 19625 20247
rect 19024 20216 19625 20244
rect 19024 20204 19030 20216
rect 19613 20213 19625 20216
rect 19659 20244 19671 20247
rect 20622 20244 20628 20256
rect 19659 20216 20628 20244
rect 19659 20213 19671 20216
rect 19613 20207 19671 20213
rect 20622 20204 20628 20216
rect 20680 20204 20686 20256
rect 20732 20253 20760 20284
rect 20717 20247 20775 20253
rect 20717 20213 20729 20247
rect 20763 20213 20775 20247
rect 20717 20207 20775 20213
rect 20898 20204 20904 20256
rect 20956 20244 20962 20256
rect 20993 20247 21051 20253
rect 20993 20244 21005 20247
rect 20956 20216 21005 20244
rect 20956 20204 20962 20216
rect 20993 20213 21005 20216
rect 21039 20213 21051 20247
rect 20993 20207 21051 20213
rect 21082 20204 21088 20256
rect 21140 20244 21146 20256
rect 21560 20244 21588 20352
rect 21818 20340 21824 20392
rect 21876 20340 21882 20392
rect 22554 20340 22560 20392
rect 22612 20380 22618 20392
rect 24026 20380 24032 20392
rect 22612 20352 24032 20380
rect 22612 20340 22618 20352
rect 24026 20340 24032 20352
rect 24084 20340 24090 20392
rect 21140 20216 21588 20244
rect 21140 20204 21146 20216
rect 1104 20154 28152 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 28152 20154
rect 1104 20080 28152 20102
rect 12161 20043 12219 20049
rect 12161 20009 12173 20043
rect 12207 20040 12219 20043
rect 12434 20040 12440 20052
rect 12207 20012 12440 20040
rect 12207 20009 12219 20012
rect 12161 20003 12219 20009
rect 12434 20000 12440 20012
rect 12492 20000 12498 20052
rect 13262 20000 13268 20052
rect 13320 20040 13326 20052
rect 13449 20043 13507 20049
rect 13449 20040 13461 20043
rect 13320 20012 13461 20040
rect 13320 20000 13326 20012
rect 13449 20009 13461 20012
rect 13495 20009 13507 20043
rect 13449 20003 13507 20009
rect 13722 20000 13728 20052
rect 13780 20040 13786 20052
rect 15286 20040 15292 20052
rect 13780 20012 15292 20040
rect 13780 20000 13786 20012
rect 15286 20000 15292 20012
rect 15344 20040 15350 20052
rect 19334 20040 19340 20052
rect 15344 20012 19340 20040
rect 15344 20000 15350 20012
rect 19306 20000 19340 20012
rect 19392 20000 19398 20052
rect 19426 20000 19432 20052
rect 19484 20040 19490 20052
rect 19521 20043 19579 20049
rect 19521 20040 19533 20043
rect 19484 20012 19533 20040
rect 19484 20000 19490 20012
rect 19521 20009 19533 20012
rect 19567 20009 19579 20043
rect 19521 20003 19579 20009
rect 19702 20000 19708 20052
rect 19760 20040 19766 20052
rect 20622 20040 20628 20052
rect 19760 20012 20628 20040
rect 19760 20000 19766 20012
rect 20622 20000 20628 20012
rect 20680 20000 20686 20052
rect 21174 20000 21180 20052
rect 21232 20040 21238 20052
rect 22189 20043 22247 20049
rect 22189 20040 22201 20043
rect 21232 20012 22201 20040
rect 21232 20000 21238 20012
rect 22189 20009 22201 20012
rect 22235 20009 22247 20043
rect 22189 20003 22247 20009
rect 22646 20000 22652 20052
rect 22704 20040 22710 20052
rect 23290 20040 23296 20052
rect 22704 20012 23296 20040
rect 22704 20000 22710 20012
rect 23290 20000 23296 20012
rect 23348 20000 23354 20052
rect 27798 20000 27804 20052
rect 27856 20000 27862 20052
rect 2590 19932 2596 19984
rect 2648 19972 2654 19984
rect 2648 19944 5672 19972
rect 2648 19932 2654 19944
rect 2038 19864 2044 19916
rect 2096 19864 2102 19916
rect 2682 19864 2688 19916
rect 2740 19864 2746 19916
rect 3142 19864 3148 19916
rect 3200 19864 3206 19916
rect 3344 19913 3372 19944
rect 3329 19907 3387 19913
rect 3329 19873 3341 19907
rect 3375 19873 3387 19907
rect 3329 19867 3387 19873
rect 3418 19864 3424 19916
rect 3476 19864 3482 19916
rect 3605 19907 3663 19913
rect 3605 19873 3617 19907
rect 3651 19904 3663 19907
rect 3651 19876 5580 19904
rect 3651 19873 3663 19876
rect 3605 19867 3663 19873
rect 842 19796 848 19848
rect 900 19836 906 19848
rect 1397 19839 1455 19845
rect 1397 19836 1409 19839
rect 900 19808 1409 19836
rect 900 19796 906 19808
rect 1397 19805 1409 19808
rect 1443 19805 1455 19839
rect 1397 19799 1455 19805
rect 2133 19839 2191 19845
rect 2133 19805 2145 19839
rect 2179 19836 2191 19839
rect 2222 19836 2228 19848
rect 2179 19808 2228 19836
rect 2179 19805 2191 19808
rect 2133 19799 2191 19805
rect 2222 19796 2228 19808
rect 2280 19796 2286 19848
rect 4448 19845 4476 19876
rect 3237 19839 3295 19845
rect 3237 19805 3249 19839
rect 3283 19805 3295 19839
rect 3237 19799 3295 19805
rect 4433 19839 4491 19845
rect 4433 19805 4445 19839
rect 4479 19805 4491 19839
rect 4433 19799 4491 19805
rect 2958 19728 2964 19780
rect 3016 19768 3022 19780
rect 3252 19768 3280 19799
rect 4706 19796 4712 19848
rect 4764 19836 4770 19848
rect 5552 19845 5580 19876
rect 5353 19839 5411 19845
rect 5353 19836 5365 19839
rect 4764 19808 5365 19836
rect 4764 19796 4770 19808
rect 5353 19805 5365 19808
rect 5399 19805 5411 19839
rect 5353 19799 5411 19805
rect 5537 19839 5595 19845
rect 5537 19805 5549 19839
rect 5583 19805 5595 19839
rect 5644 19836 5672 19944
rect 12342 19932 12348 19984
rect 12400 19972 12406 19984
rect 12713 19975 12771 19981
rect 12713 19972 12725 19975
rect 12400 19944 12725 19972
rect 12400 19932 12406 19944
rect 12713 19941 12725 19944
rect 12759 19941 12771 19975
rect 12713 19935 12771 19941
rect 13998 19932 14004 19984
rect 14056 19972 14062 19984
rect 14093 19975 14151 19981
rect 14093 19972 14105 19975
rect 14056 19944 14105 19972
rect 14056 19932 14062 19944
rect 14093 19941 14105 19944
rect 14139 19941 14151 19975
rect 14093 19935 14151 19941
rect 15010 19932 15016 19984
rect 15068 19972 15074 19984
rect 18966 19972 18972 19984
rect 15068 19944 18972 19972
rect 15068 19932 15074 19944
rect 18966 19932 18972 19944
rect 19024 19932 19030 19984
rect 19306 19972 19334 20000
rect 22278 19972 22284 19984
rect 19306 19944 20852 19972
rect 7745 19907 7803 19913
rect 7745 19873 7757 19907
rect 7791 19904 7803 19907
rect 8294 19904 8300 19916
rect 7791 19876 8300 19904
rect 7791 19873 7803 19876
rect 7745 19867 7803 19873
rect 8294 19864 8300 19876
rect 8352 19864 8358 19916
rect 10321 19907 10379 19913
rect 10321 19873 10333 19907
rect 10367 19904 10379 19907
rect 11606 19904 11612 19916
rect 10367 19876 11612 19904
rect 10367 19873 10379 19876
rect 10321 19867 10379 19873
rect 11606 19864 11612 19876
rect 11664 19864 11670 19916
rect 12069 19907 12127 19913
rect 12069 19873 12081 19907
rect 12115 19904 12127 19907
rect 12526 19904 12532 19916
rect 12115 19876 12532 19904
rect 12115 19873 12127 19876
rect 12069 19867 12127 19873
rect 6362 19836 6368 19848
rect 5644 19808 6368 19836
rect 5537 19799 5595 19805
rect 6362 19796 6368 19808
rect 6420 19836 6426 19848
rect 7653 19839 7711 19845
rect 7653 19836 7665 19839
rect 6420 19808 7665 19836
rect 6420 19796 6426 19808
rect 7653 19805 7665 19808
rect 7699 19836 7711 19839
rect 7926 19836 7932 19848
rect 7699 19808 7932 19836
rect 7699 19805 7711 19808
rect 7653 19799 7711 19805
rect 7926 19796 7932 19808
rect 7984 19796 7990 19848
rect 12360 19845 12388 19876
rect 12526 19864 12532 19876
rect 12584 19904 12590 19916
rect 12584 19876 12664 19904
rect 12584 19864 12590 19876
rect 12636 19845 12664 19876
rect 14182 19864 14188 19916
rect 14240 19904 14246 19916
rect 14369 19907 14427 19913
rect 14369 19904 14381 19907
rect 14240 19876 14381 19904
rect 14240 19864 14246 19876
rect 14369 19873 14381 19876
rect 14415 19873 14427 19907
rect 14369 19867 14427 19873
rect 14734 19864 14740 19916
rect 14792 19904 14798 19916
rect 17954 19904 17960 19916
rect 14792 19876 17960 19904
rect 14792 19864 14798 19876
rect 17954 19864 17960 19876
rect 18012 19864 18018 19916
rect 12345 19839 12403 19845
rect 12345 19805 12357 19839
rect 12391 19805 12403 19839
rect 12345 19799 12403 19805
rect 12621 19839 12679 19845
rect 12621 19805 12633 19839
rect 12667 19805 12679 19839
rect 12621 19799 12679 19805
rect 12802 19796 12808 19848
rect 12860 19796 12866 19848
rect 13630 19796 13636 19848
rect 13688 19796 13694 19848
rect 13817 19839 13875 19845
rect 13817 19805 13829 19839
rect 13863 19805 13875 19839
rect 13817 19799 13875 19805
rect 4522 19768 4528 19780
rect 3016 19740 4528 19768
rect 3016 19728 3022 19740
rect 4522 19728 4528 19740
rect 4580 19728 4586 19780
rect 9490 19768 9496 19780
rect 5000 19740 9496 19768
rect 1581 19703 1639 19709
rect 1581 19669 1593 19703
rect 1627 19700 1639 19703
rect 2314 19700 2320 19712
rect 1627 19672 2320 19700
rect 1627 19669 1639 19672
rect 1581 19663 1639 19669
rect 2314 19660 2320 19672
rect 2372 19700 2378 19712
rect 5000 19700 5028 19740
rect 9490 19728 9496 19740
rect 9548 19728 9554 19780
rect 10597 19771 10655 19777
rect 10597 19737 10609 19771
rect 10643 19737 10655 19771
rect 12434 19768 12440 19780
rect 11822 19740 12440 19768
rect 10597 19731 10655 19737
rect 2372 19672 5028 19700
rect 5261 19703 5319 19709
rect 2372 19660 2378 19672
rect 5261 19669 5273 19703
rect 5307 19700 5319 19703
rect 5350 19700 5356 19712
rect 5307 19672 5356 19700
rect 5307 19669 5319 19672
rect 5261 19663 5319 19669
rect 5350 19660 5356 19672
rect 5408 19660 5414 19712
rect 5537 19703 5595 19709
rect 5537 19669 5549 19703
rect 5583 19700 5595 19703
rect 5994 19700 6000 19712
rect 5583 19672 6000 19700
rect 5583 19669 5595 19672
rect 5537 19663 5595 19669
rect 5994 19660 6000 19672
rect 6052 19660 6058 19712
rect 8021 19703 8079 19709
rect 8021 19669 8033 19703
rect 8067 19700 8079 19703
rect 8754 19700 8760 19712
rect 8067 19672 8760 19700
rect 8067 19669 8079 19672
rect 8021 19663 8079 19669
rect 8754 19660 8760 19672
rect 8812 19660 8818 19712
rect 10612 19700 10640 19731
rect 12434 19728 12440 19740
rect 12492 19728 12498 19780
rect 12529 19771 12587 19777
rect 12529 19737 12541 19771
rect 12575 19768 12587 19771
rect 12820 19768 12848 19796
rect 12575 19740 12848 19768
rect 13832 19768 13860 19799
rect 13906 19796 13912 19848
rect 13964 19836 13970 19848
rect 14461 19839 14519 19845
rect 14461 19836 14473 19839
rect 13964 19808 14473 19836
rect 13964 19796 13970 19808
rect 14461 19805 14473 19808
rect 14507 19805 14519 19839
rect 14461 19799 14519 19805
rect 19705 19839 19763 19845
rect 19705 19805 19717 19839
rect 19751 19805 19763 19839
rect 19705 19799 19763 19805
rect 19889 19839 19947 19845
rect 19889 19805 19901 19839
rect 19935 19836 19947 19839
rect 20714 19836 20720 19848
rect 19935 19808 20720 19836
rect 19935 19805 19947 19808
rect 19889 19799 19947 19805
rect 13998 19768 14004 19780
rect 13832 19740 14004 19768
rect 12575 19737 12587 19740
rect 12529 19731 12587 19737
rect 13998 19728 14004 19740
rect 14056 19728 14062 19780
rect 15102 19728 15108 19780
rect 15160 19768 15166 19780
rect 19720 19768 19748 19799
rect 20714 19796 20720 19808
rect 20772 19796 20778 19848
rect 20824 19836 20852 19944
rect 21284 19944 22284 19972
rect 20993 19907 21051 19913
rect 20993 19873 21005 19907
rect 21039 19904 21051 19907
rect 21082 19904 21088 19916
rect 21039 19876 21088 19904
rect 21039 19873 21051 19876
rect 20993 19867 21051 19873
rect 21082 19864 21088 19876
rect 21140 19864 21146 19916
rect 21284 19845 21312 19944
rect 22278 19932 22284 19944
rect 22336 19932 22342 19984
rect 21450 19864 21456 19916
rect 21508 19904 21514 19916
rect 21545 19907 21603 19913
rect 21545 19904 21557 19907
rect 21508 19876 21557 19904
rect 21508 19864 21514 19876
rect 21545 19873 21557 19876
rect 21591 19873 21603 19907
rect 22186 19904 22192 19916
rect 21545 19867 21603 19873
rect 21652 19876 21864 19904
rect 21177 19839 21235 19845
rect 20824 19808 21128 19836
rect 20806 19768 20812 19780
rect 15160 19740 19656 19768
rect 19720 19740 20812 19768
rect 15160 19728 15166 19740
rect 11882 19700 11888 19712
rect 10612 19672 11888 19700
rect 11882 19660 11888 19672
rect 11940 19660 11946 19712
rect 12250 19660 12256 19712
rect 12308 19700 12314 19712
rect 15194 19700 15200 19712
rect 12308 19672 15200 19700
rect 12308 19660 12314 19672
rect 15194 19660 15200 19672
rect 15252 19700 15258 19712
rect 16482 19700 16488 19712
rect 15252 19672 16488 19700
rect 15252 19660 15258 19672
rect 16482 19660 16488 19672
rect 16540 19660 16546 19712
rect 19628 19700 19656 19740
rect 20806 19728 20812 19740
rect 20864 19728 20870 19780
rect 19794 19700 19800 19712
rect 19628 19672 19800 19700
rect 19794 19660 19800 19672
rect 19852 19660 19858 19712
rect 19886 19660 19892 19712
rect 19944 19700 19950 19712
rect 20993 19703 21051 19709
rect 20993 19700 21005 19703
rect 19944 19672 21005 19700
rect 19944 19660 19950 19672
rect 20993 19669 21005 19672
rect 21039 19669 21051 19703
rect 21100 19700 21128 19808
rect 21177 19805 21189 19839
rect 21223 19805 21235 19839
rect 21177 19799 21235 19805
rect 21269 19839 21327 19845
rect 21269 19805 21281 19839
rect 21315 19805 21327 19839
rect 21269 19799 21327 19805
rect 21192 19768 21220 19799
rect 21358 19796 21364 19848
rect 21416 19836 21422 19848
rect 21652 19836 21680 19876
rect 21836 19845 21864 19876
rect 21928 19876 22192 19904
rect 21416 19808 21680 19836
rect 21729 19839 21787 19845
rect 21416 19796 21422 19808
rect 21729 19805 21741 19839
rect 21775 19805 21787 19839
rect 21729 19799 21787 19805
rect 21821 19839 21879 19845
rect 21821 19805 21833 19839
rect 21867 19805 21879 19839
rect 21821 19799 21879 19805
rect 21542 19768 21548 19780
rect 21192 19740 21548 19768
rect 21542 19728 21548 19740
rect 21600 19728 21606 19780
rect 21634 19728 21640 19780
rect 21692 19768 21698 19780
rect 21744 19768 21772 19799
rect 21928 19768 21956 19876
rect 22186 19864 22192 19876
rect 22244 19864 22250 19916
rect 22554 19864 22560 19916
rect 22612 19864 22618 19916
rect 23474 19864 23480 19916
rect 23532 19904 23538 19916
rect 24670 19904 24676 19916
rect 23532 19876 24676 19904
rect 23532 19864 23538 19876
rect 24670 19864 24676 19876
rect 24728 19904 24734 19916
rect 26053 19907 26111 19913
rect 26053 19904 26065 19907
rect 24728 19876 26065 19904
rect 24728 19864 24734 19876
rect 26053 19873 26065 19876
rect 26099 19873 26111 19907
rect 26053 19867 26111 19873
rect 22002 19796 22008 19848
rect 22060 19796 22066 19848
rect 22094 19796 22100 19848
rect 22152 19796 22158 19848
rect 22370 19796 22376 19848
rect 22428 19796 22434 19848
rect 21692 19740 21956 19768
rect 21692 19728 21698 19740
rect 22278 19728 22284 19780
rect 22336 19768 22342 19780
rect 22649 19771 22707 19777
rect 22649 19768 22661 19771
rect 22336 19740 22661 19768
rect 22336 19728 22342 19740
rect 22649 19737 22661 19740
rect 22695 19737 22707 19771
rect 22649 19731 22707 19737
rect 25682 19728 25688 19780
rect 25740 19768 25746 19780
rect 26329 19771 26387 19777
rect 26329 19768 26341 19771
rect 25740 19740 26341 19768
rect 25740 19728 25746 19740
rect 26329 19737 26341 19740
rect 26375 19737 26387 19771
rect 26329 19731 26387 19737
rect 26436 19740 26818 19768
rect 22002 19700 22008 19712
rect 21100 19672 22008 19700
rect 20993 19663 21051 19669
rect 22002 19660 22008 19672
rect 22060 19660 22066 19712
rect 22094 19660 22100 19712
rect 22152 19700 22158 19712
rect 22922 19700 22928 19712
rect 22152 19672 22928 19700
rect 22152 19660 22158 19672
rect 22922 19660 22928 19672
rect 22980 19660 22986 19712
rect 24854 19660 24860 19712
rect 24912 19700 24918 19712
rect 25498 19700 25504 19712
rect 24912 19672 25504 19700
rect 24912 19660 24918 19672
rect 25498 19660 25504 19672
rect 25556 19700 25562 19712
rect 26436 19700 26464 19740
rect 25556 19672 26464 19700
rect 25556 19660 25562 19672
rect 1104 19610 28152 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 28152 19610
rect 1104 19536 28152 19558
rect 5442 19496 5448 19508
rect 4448 19468 5448 19496
rect 2869 19431 2927 19437
rect 2869 19397 2881 19431
rect 2915 19428 2927 19431
rect 2915 19400 3372 19428
rect 2915 19397 2927 19400
rect 2869 19391 2927 19397
rect 1578 19320 1584 19372
rect 1636 19360 1642 19372
rect 2590 19360 2596 19372
rect 1636 19332 2596 19360
rect 1636 19320 1642 19332
rect 2590 19320 2596 19332
rect 2648 19360 2654 19372
rect 2777 19363 2835 19369
rect 2777 19360 2789 19363
rect 2648 19332 2789 19360
rect 2648 19320 2654 19332
rect 2777 19329 2789 19332
rect 2823 19329 2835 19363
rect 2777 19323 2835 19329
rect 2958 19320 2964 19372
rect 3016 19320 3022 19372
rect 3344 19369 3372 19400
rect 4062 19388 4068 19440
rect 4120 19428 4126 19440
rect 4448 19428 4476 19468
rect 5442 19456 5448 19468
rect 5500 19456 5506 19508
rect 8021 19499 8079 19505
rect 8021 19465 8033 19499
rect 8067 19496 8079 19499
rect 8386 19496 8392 19508
rect 8067 19468 8392 19496
rect 8067 19465 8079 19468
rect 8021 19459 8079 19465
rect 8386 19456 8392 19468
rect 8444 19456 8450 19508
rect 12618 19456 12624 19508
rect 12676 19496 12682 19508
rect 15010 19496 15016 19508
rect 12676 19468 15016 19496
rect 12676 19456 12682 19468
rect 15010 19456 15016 19468
rect 15068 19456 15074 19508
rect 18782 19496 18788 19508
rect 18432 19468 18788 19496
rect 4120 19400 4476 19428
rect 4120 19388 4126 19400
rect 4448 19369 4476 19400
rect 4522 19388 4528 19440
rect 4580 19428 4586 19440
rect 5258 19428 5264 19440
rect 4580 19400 5264 19428
rect 4580 19388 4586 19400
rect 5000 19369 5028 19400
rect 5258 19388 5264 19400
rect 5316 19388 5322 19440
rect 8404 19428 8432 19456
rect 7944 19400 8340 19428
rect 8404 19400 8800 19428
rect 3329 19363 3387 19369
rect 3329 19329 3341 19363
rect 3375 19329 3387 19363
rect 3329 19323 3387 19329
rect 4433 19363 4491 19369
rect 4433 19329 4445 19363
rect 4479 19329 4491 19363
rect 4433 19323 4491 19329
rect 4985 19363 5043 19369
rect 4985 19329 4997 19363
rect 5031 19329 5043 19363
rect 4985 19323 5043 19329
rect 5077 19363 5135 19369
rect 5077 19329 5089 19363
rect 5123 19329 5135 19363
rect 5077 19323 5135 19329
rect 3418 19252 3424 19304
rect 3476 19252 3482 19304
rect 4062 19252 4068 19304
rect 4120 19252 4126 19304
rect 4706 19252 4712 19304
rect 4764 19292 4770 19304
rect 5092 19292 5120 19323
rect 5350 19320 5356 19372
rect 5408 19360 5414 19372
rect 5445 19363 5503 19369
rect 5445 19360 5457 19363
rect 5408 19332 5457 19360
rect 5408 19320 5414 19332
rect 5445 19329 5457 19332
rect 5491 19329 5503 19363
rect 5445 19323 5503 19329
rect 5994 19320 6000 19372
rect 6052 19320 6058 19372
rect 6365 19363 6423 19369
rect 6365 19360 6377 19363
rect 6196 19332 6377 19360
rect 4764 19264 5120 19292
rect 4764 19252 4770 19264
rect 6086 19116 6092 19168
rect 6144 19156 6150 19168
rect 6196 19165 6224 19332
rect 6365 19329 6377 19332
rect 6411 19329 6423 19363
rect 6365 19323 6423 19329
rect 6546 19320 6552 19372
rect 6604 19320 6610 19372
rect 7944 19369 7972 19400
rect 7929 19363 7987 19369
rect 7929 19329 7941 19363
rect 7975 19329 7987 19363
rect 7929 19323 7987 19329
rect 8202 19320 8208 19372
rect 8260 19320 8266 19372
rect 8312 19360 8340 19400
rect 8570 19360 8576 19372
rect 8312 19332 8576 19360
rect 8570 19320 8576 19332
rect 8628 19320 8634 19372
rect 8772 19369 8800 19400
rect 12434 19388 12440 19440
rect 12492 19428 12498 19440
rect 13262 19428 13268 19440
rect 12492 19400 13268 19428
rect 12492 19388 12498 19400
rect 13262 19388 13268 19400
rect 13320 19388 13326 19440
rect 14090 19388 14096 19440
rect 14148 19428 14154 19440
rect 14366 19428 14372 19440
rect 14148 19400 14372 19428
rect 14148 19388 14154 19400
rect 14366 19388 14372 19400
rect 14424 19428 14430 19440
rect 15102 19428 15108 19440
rect 14424 19400 15108 19428
rect 14424 19388 14430 19400
rect 15102 19388 15108 19400
rect 15160 19388 15166 19440
rect 16298 19388 16304 19440
rect 16356 19428 16362 19440
rect 18432 19437 18460 19468
rect 18782 19456 18788 19468
rect 18840 19456 18846 19508
rect 20717 19499 20775 19505
rect 20717 19496 20729 19499
rect 19168 19468 20729 19496
rect 19168 19437 19196 19468
rect 20717 19465 20729 19468
rect 20763 19465 20775 19499
rect 20717 19459 20775 19465
rect 20806 19456 20812 19508
rect 20864 19496 20870 19508
rect 21634 19496 21640 19508
rect 20864 19468 21640 19496
rect 20864 19456 20870 19468
rect 21634 19456 21640 19468
rect 21692 19496 21698 19508
rect 21821 19499 21879 19505
rect 21821 19496 21833 19499
rect 21692 19468 21833 19496
rect 21692 19456 21698 19468
rect 21821 19465 21833 19468
rect 21867 19465 21879 19499
rect 21821 19459 21879 19465
rect 22066 19468 22600 19496
rect 18417 19431 18475 19437
rect 18417 19428 18429 19431
rect 16356 19400 18429 19428
rect 16356 19388 16362 19400
rect 18417 19397 18429 19400
rect 18463 19397 18475 19431
rect 18417 19391 18475 19397
rect 18601 19431 18659 19437
rect 18601 19397 18613 19431
rect 18647 19428 18659 19431
rect 19153 19431 19211 19437
rect 18647 19400 19104 19428
rect 18647 19397 18659 19400
rect 18601 19391 18659 19397
rect 8757 19363 8815 19369
rect 8757 19329 8769 19363
rect 8803 19329 8815 19363
rect 8757 19323 8815 19329
rect 12526 19320 12532 19372
rect 12584 19360 12590 19372
rect 12805 19363 12863 19369
rect 12805 19360 12817 19363
rect 12584 19332 12817 19360
rect 12584 19320 12590 19332
rect 12805 19329 12817 19332
rect 12851 19329 12863 19363
rect 12805 19323 12863 19329
rect 18046 19320 18052 19372
rect 18104 19360 18110 19372
rect 18690 19360 18696 19372
rect 18104 19332 18696 19360
rect 18104 19320 18110 19332
rect 18690 19320 18696 19332
rect 18748 19320 18754 19372
rect 18966 19320 18972 19372
rect 19024 19320 19030 19372
rect 19076 19360 19104 19400
rect 19153 19397 19165 19431
rect 19199 19397 19211 19431
rect 19153 19391 19211 19397
rect 19518 19388 19524 19440
rect 19576 19428 19582 19440
rect 19576 19400 19932 19428
rect 19576 19388 19582 19400
rect 19076 19332 19380 19360
rect 12710 19252 12716 19304
rect 12768 19252 12774 19304
rect 12897 19295 12955 19301
rect 12897 19261 12909 19295
rect 12943 19261 12955 19295
rect 12897 19255 12955 19261
rect 9766 19184 9772 19236
rect 9824 19184 9830 19236
rect 12912 19224 12940 19255
rect 12986 19252 12992 19304
rect 13044 19292 13050 19304
rect 13998 19292 14004 19304
rect 13044 19264 14004 19292
rect 13044 19252 13050 19264
rect 13998 19252 14004 19264
rect 14056 19292 14062 19304
rect 14366 19292 14372 19304
rect 14056 19264 14372 19292
rect 14056 19252 14062 19264
rect 14366 19252 14372 19264
rect 14424 19252 14430 19304
rect 19352 19292 19380 19332
rect 19426 19320 19432 19372
rect 19484 19320 19490 19372
rect 19794 19320 19800 19372
rect 19852 19320 19858 19372
rect 19518 19292 19524 19304
rect 19352 19264 19524 19292
rect 19518 19252 19524 19264
rect 19576 19252 19582 19304
rect 19705 19295 19763 19301
rect 19705 19261 19717 19295
rect 19751 19261 19763 19295
rect 19705 19255 19763 19261
rect 13722 19224 13728 19236
rect 12912 19196 13728 19224
rect 13722 19184 13728 19196
rect 13780 19184 13786 19236
rect 18785 19227 18843 19233
rect 18785 19193 18797 19227
rect 18831 19224 18843 19227
rect 19720 19224 19748 19255
rect 18831 19196 19748 19224
rect 19797 19227 19855 19233
rect 18831 19193 18843 19196
rect 18785 19187 18843 19193
rect 19797 19193 19809 19227
rect 19843 19193 19855 19227
rect 19904 19224 19932 19400
rect 21726 19388 21732 19440
rect 21784 19428 21790 19440
rect 21973 19431 22031 19437
rect 21973 19428 21985 19431
rect 21784 19400 21985 19428
rect 21784 19388 21790 19400
rect 21973 19397 21985 19400
rect 22019 19428 22031 19431
rect 22066 19428 22094 19468
rect 22019 19400 22094 19428
rect 22189 19431 22247 19437
rect 22019 19397 22031 19400
rect 21973 19391 22031 19397
rect 22189 19397 22201 19431
rect 22235 19428 22247 19431
rect 22281 19431 22339 19437
rect 22281 19428 22293 19431
rect 22235 19400 22293 19428
rect 22235 19397 22247 19400
rect 22189 19391 22247 19397
rect 22281 19397 22293 19400
rect 22327 19428 22339 19431
rect 22370 19428 22376 19440
rect 22327 19400 22376 19428
rect 22327 19397 22339 19400
rect 22281 19391 22339 19397
rect 22370 19388 22376 19400
rect 22428 19388 22434 19440
rect 20257 19363 20315 19369
rect 20257 19329 20269 19363
rect 20303 19360 20315 19363
rect 20438 19360 20444 19372
rect 20303 19332 20444 19360
rect 20303 19329 20315 19332
rect 20257 19323 20315 19329
rect 20438 19320 20444 19332
rect 20496 19320 20502 19372
rect 20533 19363 20591 19369
rect 20533 19329 20545 19363
rect 20579 19360 20591 19363
rect 20625 19363 20683 19369
rect 20625 19360 20637 19363
rect 20579 19332 20637 19360
rect 20579 19329 20591 19332
rect 20533 19323 20591 19329
rect 20625 19329 20637 19332
rect 20671 19360 20683 19363
rect 20714 19360 20720 19372
rect 20671 19332 20720 19360
rect 20671 19329 20683 19332
rect 20625 19323 20683 19329
rect 20714 19320 20720 19332
rect 20772 19320 20778 19372
rect 20806 19320 20812 19372
rect 20864 19320 20870 19372
rect 22572 19369 22600 19468
rect 22465 19363 22523 19369
rect 22465 19329 22477 19363
rect 22511 19329 22523 19363
rect 22465 19323 22523 19329
rect 22557 19363 22615 19369
rect 22557 19329 22569 19363
rect 22603 19329 22615 19363
rect 22557 19323 22615 19329
rect 20441 19227 20499 19233
rect 20441 19224 20453 19227
rect 19904 19196 20453 19224
rect 19797 19187 19855 19193
rect 20441 19193 20453 19196
rect 20487 19193 20499 19227
rect 20441 19187 20499 19193
rect 6181 19159 6239 19165
rect 6181 19156 6193 19159
rect 6144 19128 6193 19156
rect 6144 19116 6150 19128
rect 6181 19125 6193 19128
rect 6227 19125 6239 19159
rect 6181 19119 6239 19125
rect 6454 19116 6460 19168
rect 6512 19116 6518 19168
rect 8205 19159 8263 19165
rect 8205 19125 8217 19159
rect 8251 19156 8263 19159
rect 8386 19156 8392 19168
rect 8251 19128 8392 19156
rect 8251 19125 8263 19128
rect 8205 19119 8263 19125
rect 8386 19116 8392 19128
rect 8444 19116 8450 19168
rect 12526 19116 12532 19168
rect 12584 19116 12590 19168
rect 13630 19116 13636 19168
rect 13688 19156 13694 19168
rect 14458 19156 14464 19168
rect 13688 19128 14464 19156
rect 13688 19116 13694 19128
rect 14458 19116 14464 19128
rect 14516 19116 14522 19168
rect 18417 19159 18475 19165
rect 18417 19125 18429 19159
rect 18463 19156 18475 19159
rect 18690 19156 18696 19168
rect 18463 19128 18696 19156
rect 18463 19125 18475 19128
rect 18417 19119 18475 19125
rect 18690 19116 18696 19128
rect 18748 19116 18754 19168
rect 18966 19116 18972 19168
rect 19024 19156 19030 19168
rect 19812 19156 19840 19187
rect 22278 19184 22284 19236
rect 22336 19184 22342 19236
rect 19024 19128 19840 19156
rect 19024 19116 19030 19128
rect 21634 19116 21640 19168
rect 21692 19156 21698 19168
rect 22005 19159 22063 19165
rect 22005 19156 22017 19159
rect 21692 19128 22017 19156
rect 21692 19116 21698 19128
rect 22005 19125 22017 19128
rect 22051 19156 22063 19159
rect 22480 19156 22508 19323
rect 22051 19128 22508 19156
rect 22051 19125 22063 19128
rect 22005 19119 22063 19125
rect 1104 19066 28152 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 28152 19066
rect 1104 18992 28152 19014
rect 8202 18912 8208 18964
rect 8260 18912 8266 18964
rect 12989 18955 13047 18961
rect 12989 18952 13001 18955
rect 12268 18924 13001 18952
rect 8662 18776 8668 18828
rect 8720 18816 8726 18828
rect 9033 18819 9091 18825
rect 9033 18816 9045 18819
rect 8720 18788 9045 18816
rect 8720 18776 8726 18788
rect 9033 18785 9045 18788
rect 9079 18816 9091 18819
rect 9079 18788 9812 18816
rect 9079 18785 9091 18788
rect 9033 18779 9091 18785
rect 4798 18708 4804 18760
rect 4856 18748 4862 18760
rect 4893 18751 4951 18757
rect 4893 18748 4905 18751
rect 4856 18720 4905 18748
rect 4856 18708 4862 18720
rect 4893 18717 4905 18720
rect 4939 18717 4951 18751
rect 4893 18711 4951 18717
rect 5350 18708 5356 18760
rect 5408 18708 5414 18760
rect 6086 18708 6092 18760
rect 6144 18708 6150 18760
rect 6546 18708 6552 18760
rect 6604 18708 6610 18760
rect 8294 18708 8300 18760
rect 8352 18748 8358 18760
rect 8389 18751 8447 18757
rect 8389 18748 8401 18751
rect 8352 18720 8401 18748
rect 8352 18708 8358 18720
rect 8389 18717 8401 18720
rect 8435 18717 8447 18751
rect 8389 18711 8447 18717
rect 8481 18751 8539 18757
rect 8481 18717 8493 18751
rect 8527 18748 8539 18751
rect 8570 18748 8576 18760
rect 8527 18720 8576 18748
rect 8527 18717 8539 18720
rect 8481 18711 8539 18717
rect 8570 18708 8576 18720
rect 8628 18708 8634 18760
rect 8754 18708 8760 18760
rect 8812 18748 8818 18760
rect 9784 18757 9812 18788
rect 9125 18751 9183 18757
rect 9125 18748 9137 18751
rect 8812 18720 9137 18748
rect 8812 18708 8818 18720
rect 9125 18717 9137 18720
rect 9171 18748 9183 18751
rect 9585 18751 9643 18757
rect 9585 18748 9597 18751
rect 9171 18720 9597 18748
rect 9171 18717 9183 18720
rect 9125 18711 9183 18717
rect 9585 18717 9597 18720
rect 9631 18717 9643 18751
rect 9585 18711 9643 18717
rect 9769 18751 9827 18757
rect 9769 18717 9781 18751
rect 9815 18717 9827 18751
rect 12268 18748 12296 18924
rect 12989 18921 13001 18924
rect 13035 18921 13047 18955
rect 12989 18915 13047 18921
rect 12342 18844 12348 18896
rect 12400 18884 12406 18896
rect 13004 18884 13032 18915
rect 13814 18912 13820 18964
rect 13872 18952 13878 18964
rect 14093 18955 14151 18961
rect 14093 18952 14105 18955
rect 13872 18924 14105 18952
rect 13872 18912 13878 18924
rect 14093 18921 14105 18924
rect 14139 18921 14151 18955
rect 14093 18915 14151 18921
rect 24210 18912 24216 18964
rect 24268 18912 24274 18964
rect 12400 18856 12480 18884
rect 13004 18856 13860 18884
rect 12400 18844 12406 18856
rect 12452 18825 12480 18856
rect 13832 18825 13860 18856
rect 12437 18819 12495 18825
rect 12437 18785 12449 18819
rect 12483 18785 12495 18819
rect 12437 18779 12495 18785
rect 13817 18819 13875 18825
rect 13817 18785 13829 18819
rect 13863 18816 13875 18819
rect 13906 18816 13912 18828
rect 13863 18788 13912 18816
rect 13863 18785 13875 18788
rect 13817 18779 13875 18785
rect 12345 18751 12403 18757
rect 12345 18748 12357 18751
rect 12268 18720 12357 18748
rect 9769 18711 9827 18717
rect 12345 18717 12357 18720
rect 12391 18717 12403 18751
rect 12452 18748 12480 18779
rect 13906 18776 13912 18788
rect 13964 18776 13970 18828
rect 14292 18788 14780 18816
rect 12805 18751 12863 18757
rect 12805 18748 12817 18751
rect 12452 18720 12817 18748
rect 12345 18711 12403 18717
rect 12805 18717 12817 18720
rect 12851 18717 12863 18751
rect 12805 18711 12863 18717
rect 12894 18708 12900 18760
rect 12952 18708 12958 18760
rect 13722 18708 13728 18760
rect 13780 18748 13786 18760
rect 14292 18748 14320 18788
rect 13780 18720 14320 18748
rect 13780 18708 13786 18720
rect 14366 18708 14372 18760
rect 14424 18708 14430 18760
rect 14458 18708 14464 18760
rect 14516 18708 14522 18760
rect 14752 18757 14780 18788
rect 17972 18788 18736 18816
rect 14553 18751 14611 18757
rect 14553 18717 14565 18751
rect 14599 18717 14611 18751
rect 14553 18711 14611 18717
rect 14737 18751 14795 18757
rect 14737 18717 14749 18751
rect 14783 18748 14795 18751
rect 15378 18748 15384 18760
rect 14783 18720 15384 18748
rect 14783 18717 14795 18720
rect 14737 18711 14795 18717
rect 7650 18680 7656 18692
rect 7406 18652 7656 18680
rect 7650 18640 7656 18652
rect 7708 18640 7714 18692
rect 14090 18640 14096 18692
rect 14148 18680 14154 18692
rect 14568 18680 14596 18711
rect 15378 18708 15384 18720
rect 15436 18708 15442 18760
rect 17972 18757 18000 18788
rect 18708 18760 18736 18788
rect 21818 18776 21824 18828
rect 21876 18816 21882 18828
rect 22465 18819 22523 18825
rect 22465 18816 22477 18819
rect 21876 18788 22477 18816
rect 21876 18776 21882 18788
rect 22465 18785 22477 18788
rect 22511 18816 22523 18819
rect 23382 18816 23388 18828
rect 22511 18788 23388 18816
rect 22511 18785 22523 18788
rect 22465 18779 22523 18785
rect 23382 18776 23388 18788
rect 23440 18776 23446 18828
rect 17957 18751 18015 18757
rect 17957 18717 17969 18751
rect 18003 18717 18015 18751
rect 17957 18711 18015 18717
rect 18138 18708 18144 18760
rect 18196 18708 18202 18760
rect 18414 18708 18420 18760
rect 18472 18708 18478 18760
rect 18601 18751 18659 18757
rect 18601 18717 18613 18751
rect 18647 18717 18659 18751
rect 18601 18711 18659 18717
rect 18322 18689 18328 18692
rect 14148 18652 14596 18680
rect 18049 18683 18107 18689
rect 14148 18640 14154 18652
rect 18049 18649 18061 18683
rect 18095 18649 18107 18683
rect 18049 18643 18107 18649
rect 18279 18683 18328 18689
rect 18279 18649 18291 18683
rect 18325 18649 18328 18683
rect 18279 18643 18328 18649
rect 5718 18572 5724 18624
rect 5776 18572 5782 18624
rect 9214 18572 9220 18624
rect 9272 18612 9278 18624
rect 9493 18615 9551 18621
rect 9493 18612 9505 18615
rect 9272 18584 9505 18612
rect 9272 18572 9278 18584
rect 9493 18581 9505 18584
rect 9539 18581 9551 18615
rect 9493 18575 9551 18581
rect 9674 18572 9680 18624
rect 9732 18572 9738 18624
rect 12710 18572 12716 18624
rect 12768 18572 12774 18624
rect 13170 18572 13176 18624
rect 13228 18572 13234 18624
rect 17310 18572 17316 18624
rect 17368 18612 17374 18624
rect 17773 18615 17831 18621
rect 17773 18612 17785 18615
rect 17368 18584 17785 18612
rect 17368 18572 17374 18584
rect 17773 18581 17785 18584
rect 17819 18581 17831 18615
rect 18064 18612 18092 18643
rect 18322 18640 18328 18643
rect 18380 18680 18386 18692
rect 18506 18680 18512 18692
rect 18380 18652 18512 18680
rect 18380 18640 18386 18652
rect 18506 18640 18512 18652
rect 18564 18640 18570 18692
rect 18616 18680 18644 18711
rect 18690 18708 18696 18760
rect 18748 18708 18754 18760
rect 18966 18680 18972 18692
rect 18616 18652 18972 18680
rect 18616 18612 18644 18652
rect 18966 18640 18972 18652
rect 19024 18640 19030 18692
rect 19702 18640 19708 18692
rect 19760 18680 19766 18692
rect 20073 18683 20131 18689
rect 20073 18680 20085 18683
rect 19760 18652 20085 18680
rect 19760 18640 19766 18652
rect 20073 18649 20085 18652
rect 20119 18649 20131 18683
rect 20073 18643 20131 18649
rect 22738 18640 22744 18692
rect 22796 18640 22802 18692
rect 24026 18680 24032 18692
rect 23966 18652 24032 18680
rect 24026 18640 24032 18652
rect 24084 18640 24090 18692
rect 18064 18584 18644 18612
rect 18877 18615 18935 18621
rect 17773 18575 17831 18581
rect 18877 18581 18889 18615
rect 18923 18612 18935 18615
rect 19242 18612 19248 18624
rect 18923 18584 19248 18612
rect 18923 18581 18935 18584
rect 18877 18575 18935 18581
rect 19242 18572 19248 18584
rect 19300 18572 19306 18624
rect 1104 18522 28152 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 28152 18522
rect 1104 18448 28152 18470
rect 4798 18368 4804 18420
rect 4856 18408 4862 18420
rect 4985 18411 5043 18417
rect 4985 18408 4997 18411
rect 4856 18380 4997 18408
rect 4856 18368 4862 18380
rect 4985 18377 4997 18380
rect 5031 18377 5043 18411
rect 7285 18411 7343 18417
rect 4985 18371 5043 18377
rect 5092 18380 6868 18408
rect 1946 18300 1952 18352
rect 2004 18300 2010 18352
rect 2314 18300 2320 18352
rect 2372 18300 2378 18352
rect 5092 18340 5120 18380
rect 3344 18312 5120 18340
rect 1486 18232 1492 18284
rect 1544 18232 1550 18284
rect 2866 18232 2872 18284
rect 2924 18272 2930 18284
rect 3237 18275 3295 18281
rect 3237 18272 3249 18275
rect 2924 18244 3249 18272
rect 2924 18232 2930 18244
rect 3237 18241 3249 18244
rect 3283 18241 3295 18275
rect 3237 18235 3295 18241
rect 2958 18164 2964 18216
rect 3016 18164 3022 18216
rect 3053 18207 3111 18213
rect 3053 18173 3065 18207
rect 3099 18173 3111 18207
rect 3053 18167 3111 18173
rect 3068 18136 3096 18167
rect 3142 18164 3148 18216
rect 3200 18204 3206 18216
rect 3344 18204 3372 18312
rect 6454 18300 6460 18352
rect 6512 18340 6518 18352
rect 6733 18343 6791 18349
rect 6733 18340 6745 18343
rect 6512 18312 6745 18340
rect 6512 18300 6518 18312
rect 6733 18309 6745 18312
rect 6779 18309 6791 18343
rect 6733 18303 6791 18309
rect 4893 18275 4951 18281
rect 4893 18241 4905 18275
rect 4939 18241 4951 18275
rect 4893 18235 4951 18241
rect 5077 18275 5135 18281
rect 5077 18241 5089 18275
rect 5123 18272 5135 18275
rect 5258 18272 5264 18284
rect 5123 18244 5264 18272
rect 5123 18241 5135 18244
rect 5077 18235 5135 18241
rect 3200 18176 3372 18204
rect 3200 18164 3206 18176
rect 3878 18164 3884 18216
rect 3936 18204 3942 18216
rect 4706 18204 4712 18216
rect 3936 18176 4712 18204
rect 3936 18164 3942 18176
rect 4706 18164 4712 18176
rect 4764 18204 4770 18216
rect 4908 18204 4936 18235
rect 5258 18232 5264 18244
rect 5316 18232 5322 18284
rect 6362 18232 6368 18284
rect 6420 18232 6426 18284
rect 6840 18272 6868 18380
rect 7285 18377 7297 18411
rect 7331 18408 7343 18411
rect 8662 18408 8668 18420
rect 7331 18380 8668 18408
rect 7331 18377 7343 18380
rect 7285 18371 7343 18377
rect 8662 18368 8668 18380
rect 8720 18368 8726 18420
rect 12434 18368 12440 18420
rect 12492 18368 12498 18420
rect 12526 18368 12532 18420
rect 12584 18368 12590 18420
rect 12710 18368 12716 18420
rect 12768 18408 12774 18420
rect 12768 18380 15056 18408
rect 12768 18368 12774 18380
rect 9766 18340 9772 18352
rect 9416 18312 9772 18340
rect 7285 18275 7343 18281
rect 7285 18272 7297 18275
rect 6840 18244 7297 18272
rect 7285 18241 7297 18244
rect 7331 18272 7343 18275
rect 7558 18272 7564 18284
rect 7331 18244 7564 18272
rect 7331 18241 7343 18244
rect 7285 18235 7343 18241
rect 7558 18232 7564 18244
rect 7616 18232 7622 18284
rect 9214 18232 9220 18284
rect 9272 18232 9278 18284
rect 9416 18281 9444 18312
rect 9766 18300 9772 18312
rect 9824 18300 9830 18352
rect 10229 18343 10287 18349
rect 10229 18340 10241 18343
rect 9876 18312 10241 18340
rect 9876 18284 9904 18312
rect 10229 18309 10241 18312
rect 10275 18309 10287 18343
rect 13170 18340 13176 18352
rect 10229 18303 10287 18309
rect 12636 18312 13176 18340
rect 9401 18275 9459 18281
rect 9401 18241 9413 18275
rect 9447 18241 9459 18275
rect 9401 18235 9459 18241
rect 9493 18275 9551 18281
rect 9493 18241 9505 18275
rect 9539 18272 9551 18275
rect 9674 18272 9680 18284
rect 9539 18244 9680 18272
rect 9539 18241 9551 18244
rect 9493 18235 9551 18241
rect 9674 18232 9680 18244
rect 9732 18232 9738 18284
rect 9858 18232 9864 18284
rect 9916 18232 9922 18284
rect 10137 18275 10195 18281
rect 10137 18272 10149 18275
rect 9968 18244 10149 18272
rect 7377 18207 7435 18213
rect 4764 18176 6500 18204
rect 4764 18164 4770 18176
rect 3896 18136 3924 18164
rect 3068 18108 3924 18136
rect 1578 18028 1584 18080
rect 1636 18028 1642 18080
rect 3418 18028 3424 18080
rect 3476 18028 3482 18080
rect 6472 18077 6500 18176
rect 7377 18173 7389 18207
rect 7423 18204 7435 18207
rect 7650 18204 7656 18216
rect 7423 18176 7656 18204
rect 7423 18173 7435 18176
rect 7377 18167 7435 18173
rect 7650 18164 7656 18176
rect 7708 18164 7714 18216
rect 9232 18204 9260 18232
rect 9968 18204 9996 18244
rect 10137 18241 10149 18244
rect 10183 18241 10195 18275
rect 10137 18235 10195 18241
rect 11790 18232 11796 18284
rect 11848 18272 11854 18284
rect 12161 18275 12219 18281
rect 12161 18272 12173 18275
rect 11848 18244 12173 18272
rect 11848 18232 11854 18244
rect 12161 18241 12173 18244
rect 12207 18272 12219 18275
rect 12526 18272 12532 18284
rect 12207 18244 12532 18272
rect 12207 18241 12219 18244
rect 12161 18235 12219 18241
rect 12526 18232 12532 18244
rect 12584 18232 12590 18284
rect 12636 18281 12664 18312
rect 13170 18300 13176 18312
rect 13228 18300 13234 18352
rect 13906 18300 13912 18352
rect 13964 18340 13970 18352
rect 13964 18312 14688 18340
rect 13964 18300 13970 18312
rect 12621 18275 12679 18281
rect 12621 18241 12633 18275
rect 12667 18241 12679 18275
rect 12621 18235 12679 18241
rect 12710 18232 12716 18284
rect 12768 18272 12774 18284
rect 12986 18272 12992 18284
rect 12768 18244 12992 18272
rect 12768 18232 12774 18244
rect 12986 18232 12992 18244
rect 13044 18232 13050 18284
rect 14001 18275 14059 18281
rect 14001 18241 14013 18275
rect 14047 18272 14059 18275
rect 14182 18272 14188 18284
rect 14047 18244 14188 18272
rect 14047 18241 14059 18244
rect 14001 18235 14059 18241
rect 14182 18232 14188 18244
rect 14240 18232 14246 18284
rect 14660 18281 14688 18312
rect 15028 18281 15056 18380
rect 15930 18368 15936 18420
rect 15988 18368 15994 18420
rect 17034 18408 17040 18420
rect 16776 18380 17040 18408
rect 15654 18300 15660 18352
rect 15712 18340 15718 18352
rect 16776 18340 16804 18380
rect 17034 18368 17040 18380
rect 17092 18408 17098 18420
rect 18417 18411 18475 18417
rect 18417 18408 18429 18411
rect 17092 18380 18429 18408
rect 17092 18368 17098 18380
rect 18417 18377 18429 18380
rect 18463 18408 18475 18411
rect 18463 18380 20576 18408
rect 18463 18377 18475 18380
rect 18417 18371 18475 18377
rect 15712 18312 16804 18340
rect 15712 18300 15718 18312
rect 14645 18275 14703 18281
rect 14645 18241 14657 18275
rect 14691 18241 14703 18275
rect 14645 18235 14703 18241
rect 15013 18275 15071 18281
rect 15013 18241 15025 18275
rect 15059 18241 15071 18275
rect 15013 18235 15071 18241
rect 15102 18232 15108 18284
rect 15160 18272 15166 18284
rect 15197 18275 15255 18281
rect 15197 18272 15209 18275
rect 15160 18244 15209 18272
rect 15160 18232 15166 18244
rect 15197 18241 15209 18244
rect 15243 18272 15255 18275
rect 15838 18272 15844 18284
rect 15243 18244 15844 18272
rect 15243 18241 15255 18244
rect 15197 18235 15255 18241
rect 15838 18232 15844 18244
rect 15896 18232 15902 18284
rect 16114 18232 16120 18284
rect 16172 18232 16178 18284
rect 16776 18281 16804 18312
rect 17129 18343 17187 18349
rect 17129 18309 17141 18343
rect 17175 18340 17187 18343
rect 17175 18312 18920 18340
rect 17175 18309 17187 18312
rect 17129 18303 17187 18309
rect 16761 18275 16819 18281
rect 16224 18244 16712 18272
rect 9232 18176 9996 18204
rect 10042 18164 10048 18216
rect 10100 18164 10106 18216
rect 12250 18164 12256 18216
rect 12308 18164 12314 18216
rect 12805 18207 12863 18213
rect 12805 18173 12817 18207
rect 12851 18204 12863 18207
rect 12894 18204 12900 18216
rect 12851 18176 12900 18204
rect 12851 18173 12863 18176
rect 12805 18167 12863 18173
rect 12894 18164 12900 18176
rect 12952 18164 12958 18216
rect 14829 18207 14887 18213
rect 14829 18173 14841 18207
rect 14875 18173 14887 18207
rect 14829 18167 14887 18173
rect 14921 18207 14979 18213
rect 14921 18173 14933 18207
rect 14967 18173 14979 18207
rect 15856 18204 15884 18232
rect 16224 18204 16252 18244
rect 15856 18176 16252 18204
rect 16301 18207 16359 18213
rect 14921 18167 14979 18173
rect 16301 18173 16313 18207
rect 16347 18204 16359 18207
rect 16390 18204 16396 18216
rect 16347 18176 16396 18204
rect 16347 18173 16359 18176
rect 16301 18167 16359 18173
rect 9585 18139 9643 18145
rect 9585 18105 9597 18139
rect 9631 18136 9643 18139
rect 9674 18136 9680 18148
rect 9631 18108 9680 18136
rect 9631 18105 9643 18108
rect 9585 18099 9643 18105
rect 9674 18096 9680 18108
rect 9732 18096 9738 18148
rect 11790 18096 11796 18148
rect 11848 18136 11854 18148
rect 12268 18136 12296 18164
rect 11848 18108 12296 18136
rect 11848 18096 11854 18108
rect 6457 18071 6515 18077
rect 6457 18037 6469 18071
rect 6503 18068 6515 18071
rect 7006 18068 7012 18080
rect 6503 18040 7012 18068
rect 6503 18037 6515 18040
rect 6457 18031 6515 18037
rect 7006 18028 7012 18040
rect 7064 18028 7070 18080
rect 9401 18071 9459 18077
rect 9401 18037 9413 18071
rect 9447 18068 9459 18071
rect 9490 18068 9496 18080
rect 9447 18040 9496 18068
rect 9447 18037 9459 18040
rect 9401 18031 9459 18037
rect 9490 18028 9496 18040
rect 9548 18028 9554 18080
rect 11974 18028 11980 18080
rect 12032 18028 12038 18080
rect 14090 18028 14096 18080
rect 14148 18028 14154 18080
rect 14458 18028 14464 18080
rect 14516 18028 14522 18080
rect 14844 18068 14872 18167
rect 14936 18136 14964 18167
rect 16390 18164 16396 18176
rect 16448 18164 16454 18216
rect 16684 18204 16712 18244
rect 16761 18241 16773 18275
rect 16807 18241 16819 18275
rect 16761 18235 16819 18241
rect 17678 18204 17684 18216
rect 16684 18176 17684 18204
rect 17678 18164 17684 18176
rect 17736 18204 17742 18216
rect 18138 18204 18144 18216
rect 17736 18176 18144 18204
rect 17736 18164 17742 18176
rect 18138 18164 18144 18176
rect 18196 18164 18202 18216
rect 17586 18136 17592 18148
rect 14936 18108 17592 18136
rect 17586 18096 17592 18108
rect 17644 18096 17650 18148
rect 16850 18068 16856 18080
rect 14844 18040 16856 18068
rect 16850 18028 16856 18040
rect 16908 18028 16914 18080
rect 18892 18068 18920 18312
rect 18984 18281 19012 18380
rect 18969 18275 19027 18281
rect 18969 18241 18981 18275
rect 19015 18241 19027 18275
rect 18969 18235 19027 18241
rect 20346 18232 20352 18284
rect 20404 18232 20410 18284
rect 19242 18164 19248 18216
rect 19300 18164 19306 18216
rect 20548 18136 20576 18380
rect 20714 18368 20720 18420
rect 20772 18368 20778 18420
rect 21358 18368 21364 18420
rect 21416 18408 21422 18420
rect 21913 18411 21971 18417
rect 21913 18408 21925 18411
rect 21416 18380 21925 18408
rect 21416 18368 21422 18380
rect 21913 18377 21925 18380
rect 21959 18408 21971 18411
rect 22554 18408 22560 18420
rect 21959 18380 22560 18408
rect 21959 18377 21971 18380
rect 21913 18371 21971 18377
rect 22554 18368 22560 18380
rect 22612 18368 22618 18420
rect 20622 18300 20628 18352
rect 20680 18340 20686 18352
rect 22649 18343 22707 18349
rect 22649 18340 22661 18343
rect 20680 18312 22661 18340
rect 20680 18300 20686 18312
rect 22649 18309 22661 18312
rect 22695 18309 22707 18343
rect 22649 18303 22707 18309
rect 21821 18275 21879 18281
rect 21821 18241 21833 18275
rect 21867 18272 21879 18275
rect 22002 18272 22008 18284
rect 21867 18244 22008 18272
rect 21867 18241 21879 18244
rect 21821 18235 21879 18241
rect 22002 18232 22008 18244
rect 22060 18232 22066 18284
rect 22097 18275 22155 18281
rect 22097 18241 22109 18275
rect 22143 18272 22155 18275
rect 22143 18244 22968 18272
rect 22143 18241 22155 18244
rect 22097 18235 22155 18241
rect 22462 18136 22468 18148
rect 20548 18108 22468 18136
rect 22462 18096 22468 18108
rect 22520 18096 22526 18148
rect 19702 18068 19708 18080
rect 18892 18040 19708 18068
rect 19702 18028 19708 18040
rect 19760 18028 19766 18080
rect 22278 18028 22284 18080
rect 22336 18028 22342 18080
rect 22940 18077 22968 18244
rect 22925 18071 22983 18077
rect 22925 18037 22937 18071
rect 22971 18068 22983 18071
rect 23014 18068 23020 18080
rect 22971 18040 23020 18068
rect 22971 18037 22983 18040
rect 22925 18031 22983 18037
rect 23014 18028 23020 18040
rect 23072 18028 23078 18080
rect 1104 17978 28152 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 28152 17978
rect 1104 17904 28152 17926
rect 2958 17824 2964 17876
rect 3016 17864 3022 17876
rect 3237 17867 3295 17873
rect 3237 17864 3249 17867
rect 3016 17836 3249 17864
rect 3016 17824 3022 17836
rect 3237 17833 3249 17836
rect 3283 17833 3295 17867
rect 3237 17827 3295 17833
rect 9309 17867 9367 17873
rect 9309 17833 9321 17867
rect 9355 17864 9367 17867
rect 9582 17864 9588 17876
rect 9355 17836 9588 17864
rect 9355 17833 9367 17836
rect 9309 17827 9367 17833
rect 9582 17824 9588 17836
rect 9640 17824 9646 17876
rect 12158 17824 12164 17876
rect 12216 17824 12222 17876
rect 12250 17824 12256 17876
rect 12308 17824 12314 17876
rect 12526 17824 12532 17876
rect 12584 17864 12590 17876
rect 13446 17864 13452 17876
rect 12584 17836 13452 17864
rect 12584 17824 12590 17836
rect 13446 17824 13452 17836
rect 13504 17864 13510 17876
rect 16574 17864 16580 17876
rect 13504 17836 16580 17864
rect 13504 17824 13510 17836
rect 16574 17824 16580 17836
rect 16632 17864 16638 17876
rect 18046 17864 18052 17876
rect 16632 17836 18052 17864
rect 16632 17824 16638 17836
rect 18046 17824 18052 17836
rect 18104 17824 18110 17876
rect 3142 17796 3148 17808
rect 1688 17768 3148 17796
rect 1688 17737 1716 17768
rect 3142 17756 3148 17768
rect 3200 17756 3206 17808
rect 14458 17756 14464 17808
rect 14516 17796 14522 17808
rect 14737 17799 14795 17805
rect 14737 17796 14749 17799
rect 14516 17768 14749 17796
rect 14516 17756 14522 17768
rect 14737 17765 14749 17768
rect 14783 17765 14795 17799
rect 14737 17759 14795 17765
rect 15105 17799 15163 17805
rect 15105 17765 15117 17799
rect 15151 17765 15163 17799
rect 15105 17759 15163 17765
rect 1673 17731 1731 17737
rect 1673 17697 1685 17731
rect 1719 17697 1731 17731
rect 1673 17691 1731 17697
rect 1946 17688 1952 17740
rect 2004 17688 2010 17740
rect 2317 17731 2375 17737
rect 2317 17697 2329 17731
rect 2363 17728 2375 17731
rect 2406 17728 2412 17740
rect 2363 17700 2412 17728
rect 2363 17697 2375 17700
rect 2317 17691 2375 17697
rect 2406 17688 2412 17700
rect 2464 17728 2470 17740
rect 2464 17700 3464 17728
rect 2464 17688 2470 17700
rect 1578 17620 1584 17672
rect 1636 17620 1642 17672
rect 2590 17620 2596 17672
rect 2648 17620 2654 17672
rect 3436 17669 3464 17700
rect 8294 17688 8300 17740
rect 8352 17688 8358 17740
rect 10042 17688 10048 17740
rect 10100 17688 10106 17740
rect 12253 17731 12311 17737
rect 12253 17697 12265 17731
rect 12299 17728 12311 17731
rect 12802 17728 12808 17740
rect 12299 17700 12808 17728
rect 12299 17697 12311 17700
rect 12253 17691 12311 17697
rect 12802 17688 12808 17700
rect 12860 17688 12866 17740
rect 14642 17688 14648 17740
rect 14700 17728 14706 17740
rect 15120 17728 15148 17759
rect 15194 17756 15200 17808
rect 15252 17796 15258 17808
rect 15749 17799 15807 17805
rect 15749 17796 15761 17799
rect 15252 17768 15761 17796
rect 15252 17756 15258 17768
rect 15749 17765 15761 17768
rect 15795 17765 15807 17799
rect 16114 17796 16120 17808
rect 15749 17759 15807 17765
rect 16040 17768 16120 17796
rect 14700 17700 15148 17728
rect 14700 17688 14706 17700
rect 3237 17663 3295 17669
rect 3237 17660 3249 17663
rect 2806 17646 3249 17660
rect 2792 17632 3249 17646
rect 2608 17592 2636 17620
rect 2792 17592 2820 17632
rect 3237 17629 3249 17632
rect 3283 17629 3295 17663
rect 3237 17623 3295 17629
rect 3421 17663 3479 17669
rect 3421 17629 3433 17663
rect 3467 17629 3479 17663
rect 3421 17623 3479 17629
rect 7558 17620 7564 17672
rect 7616 17620 7622 17672
rect 7650 17620 7656 17672
rect 7708 17620 7714 17672
rect 8846 17620 8852 17672
rect 8904 17660 8910 17672
rect 9217 17663 9275 17669
rect 9217 17660 9229 17663
rect 8904 17632 9229 17660
rect 8904 17620 8910 17632
rect 9217 17629 9229 17632
rect 9263 17629 9275 17663
rect 9217 17623 9275 17629
rect 9401 17663 9459 17669
rect 9401 17629 9413 17663
rect 9447 17660 9459 17663
rect 9490 17660 9496 17672
rect 9447 17632 9496 17660
rect 9447 17629 9459 17632
rect 9401 17623 9459 17629
rect 9490 17620 9496 17632
rect 9548 17620 9554 17672
rect 9858 17620 9864 17672
rect 9916 17620 9922 17672
rect 14182 17620 14188 17672
rect 14240 17660 14246 17672
rect 14553 17663 14611 17669
rect 14553 17660 14565 17663
rect 14240 17632 14565 17660
rect 14240 17620 14246 17632
rect 14553 17629 14565 17632
rect 14599 17629 14611 17663
rect 14553 17623 14611 17629
rect 14826 17620 14832 17672
rect 14884 17620 14890 17672
rect 15102 17620 15108 17672
rect 15160 17620 15166 17672
rect 15289 17663 15347 17669
rect 15289 17629 15301 17663
rect 15335 17660 15347 17663
rect 15378 17660 15384 17672
rect 15335 17632 15384 17660
rect 15335 17629 15347 17632
rect 15289 17623 15347 17629
rect 15378 17620 15384 17632
rect 15436 17620 15442 17672
rect 15746 17620 15752 17672
rect 15804 17620 15810 17672
rect 16040 17669 16068 17768
rect 16114 17756 16120 17768
rect 16172 17796 16178 17808
rect 16301 17799 16359 17805
rect 16301 17796 16313 17799
rect 16172 17768 16313 17796
rect 16172 17756 16178 17768
rect 16301 17765 16313 17768
rect 16347 17765 16359 17799
rect 16301 17759 16359 17765
rect 16390 17756 16396 17808
rect 16448 17796 16454 17808
rect 16945 17799 17003 17805
rect 16945 17796 16957 17799
rect 16448 17768 16957 17796
rect 16448 17756 16454 17768
rect 16945 17765 16957 17768
rect 16991 17765 17003 17799
rect 17865 17799 17923 17805
rect 17865 17796 17877 17799
rect 16945 17759 17003 17765
rect 17604 17768 17877 17796
rect 17402 17728 17408 17740
rect 16500 17700 17408 17728
rect 16025 17663 16083 17669
rect 16025 17629 16037 17663
rect 16071 17629 16083 17663
rect 16025 17623 16083 17629
rect 2608 17564 2820 17592
rect 2869 17595 2927 17601
rect 2869 17561 2881 17595
rect 2915 17592 2927 17595
rect 2958 17592 2964 17604
rect 2915 17564 2964 17592
rect 2915 17561 2927 17564
rect 2869 17555 2927 17561
rect 2958 17552 2964 17564
rect 3016 17552 3022 17604
rect 11885 17595 11943 17601
rect 11885 17561 11897 17595
rect 11931 17592 11943 17595
rect 11931 17564 12204 17592
rect 11931 17561 11943 17564
rect 11885 17555 11943 17561
rect 10594 17484 10600 17536
rect 10652 17484 10658 17536
rect 11790 17484 11796 17536
rect 11848 17524 11854 17536
rect 11977 17527 12035 17533
rect 11977 17524 11989 17527
rect 11848 17496 11989 17524
rect 11848 17484 11854 17496
rect 11977 17493 11989 17496
rect 12023 17524 12035 17527
rect 12066 17524 12072 17536
rect 12023 17496 12072 17524
rect 12023 17493 12035 17496
rect 11977 17487 12035 17493
rect 12066 17484 12072 17496
rect 12124 17484 12130 17536
rect 12176 17524 12204 17564
rect 12526 17552 12532 17604
rect 12584 17592 12590 17604
rect 15120 17592 15148 17620
rect 12584 17564 15148 17592
rect 12584 17552 12590 17564
rect 15654 17552 15660 17604
rect 15712 17592 15718 17604
rect 16040 17592 16068 17623
rect 16298 17620 16304 17672
rect 16356 17620 16362 17672
rect 16500 17669 16528 17700
rect 16485 17663 16543 17669
rect 16485 17629 16497 17663
rect 16531 17629 16543 17663
rect 16485 17623 16543 17629
rect 16574 17620 16580 17672
rect 16632 17620 16638 17672
rect 16776 17669 16804 17700
rect 17402 17688 17408 17700
rect 17460 17688 17466 17740
rect 17494 17688 17500 17740
rect 17552 17688 17558 17740
rect 17604 17672 17632 17768
rect 17865 17765 17877 17768
rect 17911 17796 17923 17799
rect 19794 17796 19800 17808
rect 17911 17768 19800 17796
rect 17911 17765 17923 17768
rect 17865 17759 17923 17765
rect 19794 17756 19800 17768
rect 19852 17796 19858 17808
rect 20990 17796 20996 17808
rect 19852 17768 20996 17796
rect 19852 17756 19858 17768
rect 20990 17756 20996 17768
rect 21048 17756 21054 17808
rect 22388 17768 22600 17796
rect 17954 17688 17960 17740
rect 18012 17728 18018 17740
rect 18012 17700 18184 17728
rect 18012 17688 18018 17700
rect 16761 17663 16819 17669
rect 16761 17629 16773 17663
rect 16807 17629 16819 17663
rect 16761 17623 16819 17629
rect 16850 17620 16856 17672
rect 16908 17620 16914 17672
rect 17221 17663 17279 17669
rect 17221 17629 17233 17663
rect 17267 17660 17279 17663
rect 17586 17660 17592 17672
rect 17267 17632 17592 17660
rect 17267 17629 17279 17632
rect 17221 17623 17279 17629
rect 17586 17620 17592 17632
rect 17644 17620 17650 17672
rect 17678 17620 17684 17672
rect 17736 17620 17742 17672
rect 18046 17620 18052 17672
rect 18104 17620 18110 17672
rect 18156 17660 18184 17700
rect 18230 17688 18236 17740
rect 18288 17728 18294 17740
rect 18288 17700 18920 17728
rect 18288 17688 18294 17700
rect 18322 17660 18328 17672
rect 18156 17632 18328 17660
rect 18322 17620 18328 17632
rect 18380 17620 18386 17672
rect 18601 17663 18659 17669
rect 18601 17629 18613 17663
rect 18647 17660 18659 17663
rect 18690 17660 18696 17672
rect 18647 17632 18696 17660
rect 18647 17629 18659 17632
rect 18601 17623 18659 17629
rect 18690 17620 18696 17632
rect 18748 17620 18754 17672
rect 18892 17669 18920 17700
rect 19150 17688 19156 17740
rect 19208 17728 19214 17740
rect 22388 17737 22416 17768
rect 21637 17731 21695 17737
rect 21637 17728 21649 17731
rect 19208 17700 21649 17728
rect 19208 17688 19214 17700
rect 21637 17697 21649 17700
rect 21683 17728 21695 17731
rect 22373 17731 22431 17737
rect 21683 17700 22324 17728
rect 21683 17697 21695 17700
rect 21637 17691 21695 17697
rect 18877 17663 18935 17669
rect 18877 17629 18889 17663
rect 18923 17629 18935 17663
rect 18877 17623 18935 17629
rect 19334 17620 19340 17672
rect 19392 17620 19398 17672
rect 20714 17620 20720 17672
rect 20772 17620 20778 17672
rect 20898 17620 20904 17672
rect 20956 17620 20962 17672
rect 20990 17620 20996 17672
rect 21048 17620 21054 17672
rect 21085 17663 21143 17669
rect 21085 17629 21097 17663
rect 21131 17629 21143 17663
rect 21085 17623 21143 17629
rect 15712 17564 16068 17592
rect 16868 17592 16896 17620
rect 19352 17592 19380 17620
rect 16868 17564 19748 17592
rect 15712 17552 15718 17564
rect 17696 17536 17724 17564
rect 12342 17524 12348 17536
rect 12176 17496 12348 17524
rect 12342 17484 12348 17496
rect 12400 17484 12406 17536
rect 15010 17484 15016 17536
rect 15068 17484 15074 17536
rect 15838 17484 15844 17536
rect 15896 17524 15902 17536
rect 15933 17527 15991 17533
rect 15933 17524 15945 17527
rect 15896 17496 15945 17524
rect 15896 17484 15902 17496
rect 15933 17493 15945 17496
rect 15979 17524 15991 17527
rect 16390 17524 16396 17536
rect 15979 17496 16396 17524
rect 15979 17493 15991 17496
rect 15933 17487 15991 17493
rect 16390 17484 16396 17496
rect 16448 17484 16454 17536
rect 17678 17484 17684 17536
rect 17736 17484 17742 17536
rect 18693 17527 18751 17533
rect 18693 17493 18705 17527
rect 18739 17524 18751 17527
rect 18966 17524 18972 17536
rect 18739 17496 18972 17524
rect 18739 17493 18751 17496
rect 18693 17487 18751 17493
rect 18966 17484 18972 17496
rect 19024 17484 19030 17536
rect 19061 17527 19119 17533
rect 19061 17493 19073 17527
rect 19107 17524 19119 17527
rect 19334 17524 19340 17536
rect 19107 17496 19340 17524
rect 19107 17493 19119 17496
rect 19061 17487 19119 17493
rect 19334 17484 19340 17496
rect 19392 17484 19398 17536
rect 19720 17524 19748 17564
rect 21100 17524 21128 17623
rect 21266 17620 21272 17672
rect 21324 17620 21330 17672
rect 21453 17663 21511 17669
rect 21453 17629 21465 17663
rect 21499 17660 21511 17663
rect 21545 17663 21603 17669
rect 21545 17660 21557 17663
rect 21499 17632 21557 17660
rect 21499 17629 21511 17632
rect 21453 17623 21511 17629
rect 21545 17629 21557 17632
rect 21591 17629 21603 17663
rect 21545 17623 21603 17629
rect 21821 17663 21879 17669
rect 21821 17629 21833 17663
rect 21867 17660 21879 17663
rect 21910 17660 21916 17672
rect 21867 17632 21916 17660
rect 21867 17629 21879 17632
rect 21821 17623 21879 17629
rect 21910 17620 21916 17632
rect 21968 17620 21974 17672
rect 22005 17663 22063 17669
rect 22005 17629 22017 17663
rect 22051 17629 22063 17663
rect 22005 17623 22063 17629
rect 21284 17592 21312 17620
rect 22020 17592 22048 17623
rect 21284 17564 22048 17592
rect 22296 17592 22324 17700
rect 22373 17697 22385 17731
rect 22419 17697 22431 17731
rect 22373 17691 22431 17697
rect 22462 17688 22468 17740
rect 22520 17688 22526 17740
rect 22572 17728 22600 17768
rect 24486 17728 24492 17740
rect 22572 17700 24492 17728
rect 24486 17688 24492 17700
rect 24544 17688 24550 17740
rect 22741 17595 22799 17601
rect 22741 17592 22753 17595
rect 22296 17564 22753 17592
rect 22741 17561 22753 17564
rect 22787 17561 22799 17595
rect 24026 17592 24032 17604
rect 23966 17564 24032 17592
rect 22741 17555 22799 17561
rect 24026 17552 24032 17564
rect 24084 17552 24090 17604
rect 22278 17524 22284 17536
rect 19720 17496 22284 17524
rect 22278 17484 22284 17496
rect 22336 17524 22342 17536
rect 22462 17524 22468 17536
rect 22336 17496 22468 17524
rect 22336 17484 22342 17496
rect 22462 17484 22468 17496
rect 22520 17484 22526 17536
rect 24210 17484 24216 17536
rect 24268 17484 24274 17536
rect 1104 17434 28152 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 28152 17434
rect 1104 17360 28152 17382
rect 2406 17280 2412 17332
rect 2464 17280 2470 17332
rect 4062 17280 4068 17332
rect 4120 17320 4126 17332
rect 7745 17323 7803 17329
rect 4120 17292 4844 17320
rect 4120 17280 4126 17292
rect 1872 17224 2544 17252
rect 1872 17196 1900 17224
rect 1854 17144 1860 17196
rect 1912 17144 1918 17196
rect 2516 17193 2544 17224
rect 3528 17224 4660 17252
rect 2317 17187 2375 17193
rect 2317 17184 2329 17187
rect 1964 17156 2329 17184
rect 1964 17128 1992 17156
rect 2317 17153 2329 17156
rect 2363 17153 2375 17187
rect 2317 17147 2375 17153
rect 2501 17187 2559 17193
rect 2501 17153 2513 17187
rect 2547 17153 2559 17187
rect 2501 17147 2559 17153
rect 3418 17144 3424 17196
rect 3476 17184 3482 17196
rect 3528 17193 3556 17224
rect 3513 17187 3571 17193
rect 3513 17184 3525 17187
rect 3476 17156 3525 17184
rect 3476 17144 3482 17156
rect 3513 17153 3525 17156
rect 3559 17153 3571 17187
rect 3513 17147 3571 17153
rect 3881 17187 3939 17193
rect 3881 17153 3893 17187
rect 3927 17184 3939 17187
rect 4062 17184 4068 17196
rect 3927 17156 4068 17184
rect 3927 17153 3939 17156
rect 3881 17147 3939 17153
rect 4062 17144 4068 17156
rect 4120 17144 4126 17196
rect 4632 17193 4660 17224
rect 4816 17193 4844 17292
rect 7745 17289 7757 17323
rect 7791 17320 7803 17323
rect 8294 17320 8300 17332
rect 7791 17292 8300 17320
rect 7791 17289 7803 17292
rect 7745 17283 7803 17289
rect 8294 17280 8300 17292
rect 8352 17280 8358 17332
rect 9309 17323 9367 17329
rect 9309 17289 9321 17323
rect 9355 17320 9367 17323
rect 10042 17320 10048 17332
rect 9355 17292 10048 17320
rect 9355 17289 9367 17292
rect 9309 17283 9367 17289
rect 10042 17280 10048 17292
rect 10100 17280 10106 17332
rect 11348 17292 15608 17320
rect 11348 17261 11376 17292
rect 11333 17255 11391 17261
rect 11333 17221 11345 17255
rect 11379 17221 11391 17255
rect 13262 17252 13268 17264
rect 13202 17224 13268 17252
rect 11333 17215 11391 17221
rect 13262 17212 13268 17224
rect 13320 17252 13326 17264
rect 15470 17252 15476 17264
rect 13320 17224 15476 17252
rect 13320 17212 13326 17224
rect 15470 17212 15476 17224
rect 15528 17212 15534 17264
rect 4617 17187 4675 17193
rect 4617 17153 4629 17187
rect 4663 17153 4675 17187
rect 4617 17147 4675 17153
rect 4801 17187 4859 17193
rect 4801 17153 4813 17187
rect 4847 17153 4859 17187
rect 4801 17147 4859 17153
rect 7558 17144 7564 17196
rect 7616 17144 7622 17196
rect 7834 17144 7840 17196
rect 7892 17144 7898 17196
rect 8662 17144 8668 17196
rect 8720 17184 8726 17196
rect 9033 17187 9091 17193
rect 9033 17184 9045 17187
rect 8720 17156 9045 17184
rect 8720 17144 8726 17156
rect 9033 17153 9045 17156
rect 9079 17153 9091 17187
rect 9033 17147 9091 17153
rect 9674 17144 9680 17196
rect 9732 17144 9738 17196
rect 9766 17144 9772 17196
rect 9824 17184 9830 17196
rect 9861 17187 9919 17193
rect 9861 17184 9873 17187
rect 9824 17156 9873 17184
rect 9824 17144 9830 17156
rect 9861 17153 9873 17156
rect 9907 17153 9919 17187
rect 9861 17147 9919 17153
rect 11606 17144 11612 17196
rect 11664 17184 11670 17196
rect 11701 17187 11759 17193
rect 11701 17184 11713 17187
rect 11664 17156 11713 17184
rect 11664 17144 11670 17156
rect 11701 17153 11713 17156
rect 11747 17153 11759 17187
rect 11701 17147 11759 17153
rect 13633 17187 13691 17193
rect 13633 17153 13645 17187
rect 13679 17153 13691 17187
rect 13633 17147 13691 17153
rect 1946 17076 1952 17128
rect 2004 17076 2010 17128
rect 4525 17119 4583 17125
rect 4525 17085 4537 17119
rect 4571 17085 4583 17119
rect 4525 17079 4583 17085
rect 2225 17051 2283 17057
rect 2225 17017 2237 17051
rect 2271 17048 2283 17051
rect 2682 17048 2688 17060
rect 2271 17020 2688 17048
rect 2271 17017 2283 17020
rect 2225 17011 2283 17017
rect 2682 17008 2688 17020
rect 2740 17008 2746 17060
rect 4540 17048 4568 17079
rect 8846 17076 8852 17128
rect 8904 17076 8910 17128
rect 8938 17076 8944 17128
rect 8996 17076 9002 17128
rect 9125 17119 9183 17125
rect 9125 17085 9137 17119
rect 9171 17085 9183 17119
rect 9125 17079 9183 17085
rect 11977 17119 12035 17125
rect 11977 17085 11989 17119
rect 12023 17116 12035 17119
rect 12710 17116 12716 17128
rect 12023 17088 12716 17116
rect 12023 17085 12035 17088
rect 11977 17079 12035 17085
rect 4614 17048 4620 17060
rect 4540 17020 4620 17048
rect 4614 17008 4620 17020
rect 4672 17008 4678 17060
rect 7561 17051 7619 17057
rect 7561 17017 7573 17051
rect 7607 17048 7619 17051
rect 8864 17048 8892 17076
rect 7607 17020 8892 17048
rect 9140 17048 9168 17079
rect 12710 17076 12716 17088
rect 12768 17116 12774 17128
rect 13648 17116 13676 17147
rect 13814 17144 13820 17196
rect 13872 17184 13878 17196
rect 14366 17184 14372 17196
rect 13872 17156 14372 17184
rect 13872 17144 13878 17156
rect 14366 17144 14372 17156
rect 14424 17144 14430 17196
rect 14458 17144 14464 17196
rect 14516 17144 14522 17196
rect 14553 17187 14611 17193
rect 14553 17153 14565 17187
rect 14599 17184 14611 17187
rect 14642 17184 14648 17196
rect 14599 17156 14648 17184
rect 14599 17153 14611 17156
rect 14553 17147 14611 17153
rect 14642 17144 14648 17156
rect 14700 17144 14706 17196
rect 12768 17088 13676 17116
rect 14277 17119 14335 17125
rect 12768 17076 12774 17088
rect 14277 17085 14289 17119
rect 14323 17116 14335 17119
rect 14323 17088 14504 17116
rect 14323 17085 14335 17088
rect 14277 17079 14335 17085
rect 10226 17048 10232 17060
rect 9140 17020 10232 17048
rect 7607 17017 7619 17020
rect 7561 17011 7619 17017
rect 10226 17008 10232 17020
rect 10284 17008 10290 17060
rect 13262 17008 13268 17060
rect 13320 17048 13326 17060
rect 14476 17048 14504 17088
rect 13320 17020 14504 17048
rect 13320 17008 13326 17020
rect 4706 16940 4712 16992
rect 4764 16940 4770 16992
rect 12618 16940 12624 16992
rect 12676 16980 12682 16992
rect 13449 16983 13507 16989
rect 13449 16980 13461 16983
rect 12676 16952 13461 16980
rect 12676 16940 12682 16952
rect 13449 16949 13461 16952
rect 13495 16949 13507 16983
rect 13449 16943 13507 16949
rect 13633 16983 13691 16989
rect 13633 16949 13645 16983
rect 13679 16980 13691 16983
rect 13998 16980 14004 16992
rect 13679 16952 14004 16980
rect 13679 16949 13691 16952
rect 13633 16943 13691 16949
rect 13998 16940 14004 16952
rect 14056 16940 14062 16992
rect 14366 16940 14372 16992
rect 14424 16940 14430 16992
rect 14476 16980 14504 17020
rect 14550 17008 14556 17060
rect 14608 17048 14614 17060
rect 15473 17051 15531 17057
rect 15473 17048 15485 17051
rect 14608 17020 15485 17048
rect 14608 17008 14614 17020
rect 15473 17017 15485 17020
rect 15519 17017 15531 17051
rect 15580 17048 15608 17292
rect 15746 17280 15752 17332
rect 15804 17320 15810 17332
rect 15804 17292 15884 17320
rect 15804 17280 15810 17292
rect 15856 17261 15884 17292
rect 18046 17280 18052 17332
rect 18104 17320 18110 17332
rect 18690 17320 18696 17332
rect 18104 17292 18696 17320
rect 18104 17280 18110 17292
rect 18690 17280 18696 17292
rect 18748 17280 18754 17332
rect 19429 17323 19487 17329
rect 19429 17289 19441 17323
rect 19475 17320 19487 17323
rect 20806 17320 20812 17332
rect 19475 17292 20812 17320
rect 19475 17289 19487 17292
rect 19429 17283 19487 17289
rect 20806 17280 20812 17292
rect 20864 17280 20870 17332
rect 20898 17280 20904 17332
rect 20956 17320 20962 17332
rect 22373 17323 22431 17329
rect 22373 17320 22385 17323
rect 20956 17292 22385 17320
rect 20956 17280 20962 17292
rect 22373 17289 22385 17292
rect 22419 17289 22431 17323
rect 22373 17283 22431 17289
rect 15841 17255 15899 17261
rect 15841 17221 15853 17255
rect 15887 17221 15899 17255
rect 20990 17252 20996 17264
rect 15841 17215 15899 17221
rect 16132 17224 20996 17252
rect 15654 17144 15660 17196
rect 15712 17144 15718 17196
rect 15746 17144 15752 17196
rect 15804 17144 15810 17196
rect 16022 17193 16028 17196
rect 15979 17187 16028 17193
rect 15979 17153 15991 17187
rect 16025 17153 16028 17187
rect 15979 17147 16028 17153
rect 16022 17144 16028 17147
rect 16080 17144 16086 17196
rect 16132 17193 16160 17224
rect 20990 17212 20996 17224
rect 21048 17212 21054 17264
rect 22741 17255 22799 17261
rect 22741 17221 22753 17255
rect 22787 17252 22799 17255
rect 23569 17255 23627 17261
rect 23569 17252 23581 17255
rect 22787 17224 23581 17252
rect 22787 17221 22799 17224
rect 22741 17215 22799 17221
rect 23569 17221 23581 17224
rect 23615 17221 23627 17255
rect 23569 17215 23627 17221
rect 16117 17187 16175 17193
rect 16117 17153 16129 17187
rect 16163 17153 16175 17187
rect 16117 17147 16175 17153
rect 16850 17144 16856 17196
rect 16908 17144 16914 17196
rect 17037 17187 17095 17193
rect 17037 17153 17049 17187
rect 17083 17184 17095 17187
rect 17126 17184 17132 17196
rect 17083 17156 17132 17184
rect 17083 17153 17095 17156
rect 17037 17147 17095 17153
rect 17126 17144 17132 17156
rect 17184 17144 17190 17196
rect 18322 17144 18328 17196
rect 18380 17184 18386 17196
rect 19058 17184 19064 17196
rect 18380 17156 19064 17184
rect 18380 17144 18386 17156
rect 19058 17144 19064 17156
rect 19116 17144 19122 17196
rect 19334 17144 19340 17196
rect 19392 17144 19398 17196
rect 19521 17187 19579 17193
rect 19521 17153 19533 17187
rect 19567 17184 19579 17187
rect 19886 17184 19892 17196
rect 19567 17156 19892 17184
rect 19567 17153 19579 17156
rect 19521 17147 19579 17153
rect 19886 17144 19892 17156
rect 19944 17144 19950 17196
rect 20073 17187 20131 17193
rect 20073 17153 20085 17187
rect 20119 17184 20131 17187
rect 21266 17184 21272 17196
rect 20119 17156 21272 17184
rect 20119 17153 20131 17156
rect 20073 17147 20131 17153
rect 21266 17144 21272 17156
rect 21324 17144 21330 17196
rect 21361 17187 21419 17193
rect 21361 17153 21373 17187
rect 21407 17153 21419 17187
rect 21361 17147 21419 17153
rect 16945 17119 17003 17125
rect 16945 17085 16957 17119
rect 16991 17116 17003 17119
rect 16991 17088 19472 17116
rect 16991 17085 17003 17088
rect 16945 17079 17003 17085
rect 17402 17048 17408 17060
rect 15580 17020 17408 17048
rect 15473 17011 15531 17017
rect 17402 17008 17408 17020
rect 17460 17008 17466 17060
rect 17954 17008 17960 17060
rect 18012 17048 18018 17060
rect 19245 17051 19303 17057
rect 19245 17048 19257 17051
rect 18012 17020 19257 17048
rect 18012 17008 18018 17020
rect 19245 17017 19257 17020
rect 19291 17017 19303 17051
rect 19444 17048 19472 17088
rect 19794 17076 19800 17128
rect 19852 17116 19858 17128
rect 19981 17119 20039 17125
rect 19981 17116 19993 17119
rect 19852 17088 19993 17116
rect 19852 17076 19858 17088
rect 19981 17085 19993 17088
rect 20027 17085 20039 17119
rect 19981 17079 20039 17085
rect 20162 17076 20168 17128
rect 20220 17116 20226 17128
rect 21376 17116 21404 17147
rect 21726 17144 21732 17196
rect 21784 17184 21790 17196
rect 22557 17187 22615 17193
rect 22557 17184 22569 17187
rect 21784 17156 22569 17184
rect 21784 17144 21790 17156
rect 22557 17153 22569 17156
rect 22603 17184 22615 17187
rect 23017 17187 23075 17193
rect 23017 17184 23029 17187
rect 22603 17156 23029 17184
rect 22603 17153 22615 17156
rect 22557 17147 22615 17153
rect 23017 17153 23029 17156
rect 23063 17153 23075 17187
rect 23017 17147 23075 17153
rect 23201 17187 23259 17193
rect 23201 17153 23213 17187
rect 23247 17184 23259 17187
rect 23474 17184 23480 17196
rect 23247 17156 23480 17184
rect 23247 17153 23259 17156
rect 23201 17147 23259 17153
rect 23474 17144 23480 17156
rect 23532 17144 23538 17196
rect 23661 17187 23719 17193
rect 23661 17153 23673 17187
rect 23707 17184 23719 17187
rect 24210 17184 24216 17196
rect 23707 17156 24216 17184
rect 23707 17153 23719 17156
rect 23661 17147 23719 17153
rect 23385 17119 23443 17125
rect 23385 17116 23397 17119
rect 20220 17088 23397 17116
rect 20220 17076 20226 17088
rect 23385 17085 23397 17088
rect 23431 17116 23443 17119
rect 23676 17116 23704 17147
rect 24210 17144 24216 17156
rect 24268 17144 24274 17196
rect 25222 17144 25228 17196
rect 25280 17144 25286 17196
rect 23431 17088 23704 17116
rect 23431 17085 23443 17088
rect 23385 17079 23443 17085
rect 24854 17076 24860 17128
rect 24912 17116 24918 17128
rect 24949 17119 25007 17125
rect 24949 17116 24961 17119
rect 24912 17088 24961 17116
rect 24912 17076 24918 17088
rect 24949 17085 24961 17088
rect 24995 17085 25007 17119
rect 24949 17079 25007 17085
rect 22738 17048 22744 17060
rect 19444 17020 22744 17048
rect 19245 17011 19303 17017
rect 22738 17008 22744 17020
rect 22796 17008 22802 17060
rect 14826 16980 14832 16992
rect 14476 16952 14832 16980
rect 14826 16940 14832 16952
rect 14884 16980 14890 16992
rect 16298 16980 16304 16992
rect 14884 16952 16304 16980
rect 14884 16940 14890 16952
rect 16298 16940 16304 16952
rect 16356 16940 16362 16992
rect 18046 16940 18052 16992
rect 18104 16980 18110 16992
rect 19150 16980 19156 16992
rect 18104 16952 19156 16980
rect 18104 16940 18110 16952
rect 19150 16940 19156 16952
rect 19208 16980 19214 16992
rect 19705 16983 19763 16989
rect 19705 16980 19717 16983
rect 19208 16952 19717 16980
rect 19208 16940 19214 16952
rect 19705 16949 19717 16952
rect 19751 16949 19763 16983
rect 19705 16943 19763 16949
rect 20349 16983 20407 16989
rect 20349 16949 20361 16983
rect 20395 16980 20407 16983
rect 20898 16980 20904 16992
rect 20395 16952 20904 16980
rect 20395 16949 20407 16952
rect 20349 16943 20407 16949
rect 20898 16940 20904 16952
rect 20956 16940 20962 16992
rect 20990 16940 20996 16992
rect 21048 16980 21054 16992
rect 23106 16980 23112 16992
rect 21048 16952 23112 16980
rect 21048 16940 21054 16952
rect 23106 16940 23112 16952
rect 23164 16940 23170 16992
rect 1104 16890 28152 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 28152 16890
rect 1104 16816 28152 16838
rect 8662 16736 8668 16788
rect 8720 16776 8726 16788
rect 8720 16748 9536 16776
rect 8720 16736 8726 16748
rect 8386 16668 8392 16720
rect 8444 16708 8450 16720
rect 8941 16711 8999 16717
rect 8941 16708 8953 16711
rect 8444 16680 8953 16708
rect 8444 16668 8450 16680
rect 8941 16677 8953 16680
rect 8987 16677 8999 16711
rect 8941 16671 8999 16677
rect 2958 16600 2964 16652
rect 3016 16600 3022 16652
rect 3510 16600 3516 16652
rect 3568 16600 3574 16652
rect 8110 16600 8116 16652
rect 8168 16600 8174 16652
rect 9306 16600 9312 16652
rect 9364 16600 9370 16652
rect 2866 16532 2872 16584
rect 2924 16532 2930 16584
rect 4709 16575 4767 16581
rect 4709 16541 4721 16575
rect 4755 16572 4767 16575
rect 5353 16575 5411 16581
rect 4755 16544 4844 16572
rect 4755 16541 4767 16544
rect 4709 16535 4767 16541
rect 4816 16516 4844 16544
rect 5353 16541 5365 16575
rect 5399 16572 5411 16575
rect 5718 16572 5724 16584
rect 5399 16544 5724 16572
rect 5399 16541 5411 16544
rect 5353 16535 5411 16541
rect 5718 16532 5724 16544
rect 5776 16532 5782 16584
rect 7374 16532 7380 16584
rect 7432 16532 7438 16584
rect 7466 16532 7472 16584
rect 7524 16572 7530 16584
rect 7561 16575 7619 16581
rect 7561 16572 7573 16575
rect 7524 16544 7573 16572
rect 7524 16532 7530 16544
rect 7561 16541 7573 16544
rect 7607 16541 7619 16575
rect 7561 16535 7619 16541
rect 8570 16532 8576 16584
rect 8628 16572 8634 16584
rect 8938 16572 8944 16584
rect 8628 16544 8944 16572
rect 8628 16532 8634 16544
rect 8938 16532 8944 16544
rect 8996 16572 9002 16584
rect 9401 16575 9459 16581
rect 9401 16572 9413 16575
rect 8996 16544 9413 16572
rect 8996 16532 9002 16544
rect 9401 16541 9413 16544
rect 9447 16541 9459 16575
rect 9508 16572 9536 16748
rect 12342 16736 12348 16788
rect 12400 16776 12406 16788
rect 12897 16779 12955 16785
rect 12897 16776 12909 16779
rect 12400 16748 12909 16776
rect 12400 16736 12406 16748
rect 12897 16745 12909 16748
rect 12943 16745 12955 16779
rect 12897 16739 12955 16745
rect 15378 16736 15384 16788
rect 15436 16776 15442 16788
rect 15841 16779 15899 16785
rect 15841 16776 15853 16779
rect 15436 16748 15853 16776
rect 15436 16736 15442 16748
rect 15841 16745 15853 16748
rect 15887 16745 15899 16779
rect 15841 16739 15899 16745
rect 16022 16736 16028 16788
rect 16080 16736 16086 16788
rect 16114 16736 16120 16788
rect 16172 16776 16178 16788
rect 20714 16776 20720 16788
rect 16172 16748 20720 16776
rect 16172 16736 16178 16748
rect 20714 16736 20720 16748
rect 20772 16736 20778 16788
rect 20806 16736 20812 16788
rect 20864 16776 20870 16788
rect 22005 16779 22063 16785
rect 22005 16776 22017 16779
rect 20864 16748 22017 16776
rect 20864 16736 20870 16748
rect 22005 16745 22017 16748
rect 22051 16745 22063 16779
rect 22005 16739 22063 16745
rect 23106 16736 23112 16788
rect 23164 16736 23170 16788
rect 11606 16668 11612 16720
rect 11664 16708 11670 16720
rect 20441 16711 20499 16717
rect 11664 16680 14136 16708
rect 11664 16668 11670 16680
rect 11974 16600 11980 16652
rect 12032 16640 12038 16652
rect 12345 16643 12403 16649
rect 12345 16640 12357 16643
rect 12032 16612 12357 16640
rect 12032 16600 12038 16612
rect 12345 16609 12357 16612
rect 12391 16609 12403 16643
rect 12345 16603 12403 16609
rect 12710 16600 12716 16652
rect 12768 16640 12774 16652
rect 14108 16649 14136 16680
rect 20441 16677 20453 16711
rect 20487 16708 20499 16711
rect 23124 16708 23152 16736
rect 20487 16680 20576 16708
rect 20487 16677 20499 16680
rect 20441 16671 20499 16677
rect 12805 16643 12863 16649
rect 12805 16640 12817 16643
rect 12768 16612 12817 16640
rect 12768 16600 12774 16612
rect 12805 16609 12817 16612
rect 12851 16609 12863 16643
rect 12805 16603 12863 16609
rect 14093 16643 14151 16649
rect 14093 16609 14105 16643
rect 14139 16640 14151 16643
rect 20162 16640 20168 16652
rect 14139 16612 16574 16640
rect 14139 16609 14151 16612
rect 14093 16603 14151 16609
rect 9861 16575 9919 16581
rect 9861 16572 9873 16575
rect 9508 16544 9873 16572
rect 9401 16535 9459 16541
rect 9861 16541 9873 16544
rect 9907 16541 9919 16575
rect 9861 16535 9919 16541
rect 10226 16532 10232 16584
rect 10284 16532 10290 16584
rect 10597 16575 10655 16581
rect 10597 16541 10609 16575
rect 10643 16541 10655 16575
rect 10597 16535 10655 16541
rect 4798 16464 4804 16516
rect 4856 16464 4862 16516
rect 7484 16504 7512 16532
rect 6026 16476 7512 16504
rect 9490 16464 9496 16516
rect 9548 16504 9554 16516
rect 10612 16504 10640 16535
rect 11882 16532 11888 16584
rect 11940 16572 11946 16584
rect 12069 16575 12127 16581
rect 12069 16572 12081 16575
rect 11940 16544 12081 16572
rect 11940 16532 11946 16544
rect 12069 16541 12081 16544
rect 12115 16541 12127 16575
rect 12069 16535 12127 16541
rect 12250 16532 12256 16584
rect 12308 16532 12314 16584
rect 12437 16575 12495 16581
rect 12437 16541 12449 16575
rect 12483 16572 12495 16575
rect 12526 16572 12532 16584
rect 12483 16544 12532 16572
rect 12483 16541 12495 16544
rect 12437 16535 12495 16541
rect 12526 16532 12532 16544
rect 12584 16532 12590 16584
rect 12618 16532 12624 16584
rect 12676 16532 12682 16584
rect 13081 16575 13139 16581
rect 13081 16541 13093 16575
rect 13127 16541 13139 16575
rect 13081 16535 13139 16541
rect 9548 16476 10640 16504
rect 9548 16464 9554 16476
rect 12158 16464 12164 16516
rect 12216 16504 12222 16516
rect 12897 16507 12955 16513
rect 12897 16504 12909 16507
rect 12216 16476 12909 16504
rect 12216 16464 12222 16476
rect 12897 16473 12909 16476
rect 12943 16473 12955 16507
rect 13096 16504 13124 16535
rect 13170 16532 13176 16584
rect 13228 16532 13234 16584
rect 16022 16532 16028 16584
rect 16080 16572 16086 16584
rect 16117 16575 16175 16581
rect 16117 16572 16129 16575
rect 16080 16544 16129 16572
rect 16080 16532 16086 16544
rect 16117 16541 16129 16544
rect 16163 16541 16175 16575
rect 16546 16572 16574 16612
rect 19904 16612 20168 16640
rect 17034 16572 17040 16584
rect 16546 16544 17040 16572
rect 16117 16535 16175 16541
rect 17034 16532 17040 16544
rect 17092 16532 17098 16584
rect 19904 16581 19932 16612
rect 20162 16600 20168 16612
rect 20220 16600 20226 16652
rect 20548 16649 20576 16680
rect 22388 16680 23152 16708
rect 20898 16649 20904 16652
rect 20533 16643 20591 16649
rect 20533 16609 20545 16643
rect 20579 16609 20591 16643
rect 20533 16603 20591 16609
rect 20897 16603 20904 16649
rect 20956 16640 20962 16652
rect 20956 16612 20997 16640
rect 20898 16600 20904 16603
rect 20956 16600 20962 16612
rect 21082 16600 21088 16652
rect 21140 16600 21146 16652
rect 21726 16600 21732 16652
rect 21784 16600 21790 16652
rect 19889 16575 19947 16581
rect 19889 16541 19901 16575
rect 19935 16541 19947 16575
rect 19889 16535 19947 16541
rect 20303 16575 20361 16581
rect 20303 16541 20315 16575
rect 20349 16572 20361 16575
rect 20438 16572 20444 16584
rect 20349 16544 20444 16572
rect 20349 16541 20361 16544
rect 20303 16535 20361 16541
rect 20438 16532 20444 16544
rect 20496 16572 20502 16584
rect 20717 16575 20775 16581
rect 20717 16572 20729 16575
rect 20496 16544 20729 16572
rect 20496 16532 20502 16544
rect 20717 16541 20729 16544
rect 20763 16541 20775 16575
rect 20717 16535 20775 16541
rect 20809 16575 20867 16581
rect 20809 16541 20821 16575
rect 20855 16572 20867 16575
rect 21177 16575 21235 16581
rect 21177 16572 21189 16575
rect 20855 16544 21189 16572
rect 20855 16541 20867 16544
rect 20809 16535 20867 16541
rect 21177 16541 21189 16544
rect 21223 16572 21235 16575
rect 21634 16572 21640 16584
rect 21223 16544 21640 16572
rect 21223 16541 21235 16544
rect 21177 16535 21235 16541
rect 13096 16476 13492 16504
rect 12897 16467 12955 16473
rect 13354 16396 13360 16448
rect 13412 16396 13418 16448
rect 13464 16436 13492 16476
rect 14366 16464 14372 16516
rect 14424 16464 14430 16516
rect 15654 16504 15660 16516
rect 15594 16476 15660 16504
rect 15654 16464 15660 16476
rect 15712 16504 15718 16516
rect 19518 16504 19524 16516
rect 15712 16476 19524 16504
rect 15712 16464 15718 16476
rect 19518 16464 19524 16476
rect 19576 16464 19582 16516
rect 20073 16507 20131 16513
rect 20073 16504 20085 16507
rect 19904 16476 20085 16504
rect 14550 16436 14556 16448
rect 13464 16408 14556 16436
rect 14550 16396 14556 16408
rect 14608 16396 14614 16448
rect 15102 16396 15108 16448
rect 15160 16436 15166 16448
rect 19794 16436 19800 16448
rect 15160 16408 19800 16436
rect 15160 16396 15166 16408
rect 19794 16396 19800 16408
rect 19852 16436 19858 16448
rect 19904 16436 19932 16476
rect 20073 16473 20085 16476
rect 20119 16473 20131 16507
rect 20073 16467 20131 16473
rect 20162 16464 20168 16516
rect 20220 16504 20226 16516
rect 20824 16504 20852 16535
rect 21634 16532 21640 16544
rect 21692 16532 21698 16584
rect 22388 16581 22416 16680
rect 24026 16668 24032 16720
rect 24084 16708 24090 16720
rect 24857 16711 24915 16717
rect 24857 16708 24869 16711
rect 24084 16680 24869 16708
rect 24084 16668 24090 16680
rect 24857 16677 24869 16680
rect 24903 16677 24915 16711
rect 24857 16671 24915 16677
rect 23017 16643 23075 16649
rect 22572 16612 22968 16640
rect 22572 16581 22600 16612
rect 22940 16584 22968 16612
rect 23017 16609 23029 16643
rect 23063 16640 23075 16643
rect 23063 16612 23520 16640
rect 23063 16609 23075 16612
rect 23017 16603 23075 16609
rect 21913 16575 21971 16581
rect 21913 16541 21925 16575
rect 21959 16541 21971 16575
rect 21913 16535 21971 16541
rect 22097 16575 22155 16581
rect 22097 16541 22109 16575
rect 22143 16572 22155 16575
rect 22373 16575 22431 16581
rect 22143 16544 22324 16572
rect 22143 16541 22155 16544
rect 22097 16535 22155 16541
rect 20220 16476 20852 16504
rect 20220 16464 20226 16476
rect 21450 16464 21456 16516
rect 21508 16504 21514 16516
rect 21928 16504 21956 16535
rect 21508 16476 21956 16504
rect 21508 16464 21514 16476
rect 22296 16448 22324 16544
rect 22373 16541 22385 16575
rect 22419 16541 22431 16575
rect 22373 16535 22431 16541
rect 22465 16575 22523 16581
rect 22465 16541 22477 16575
rect 22511 16541 22523 16575
rect 22465 16535 22523 16541
rect 22557 16575 22615 16581
rect 22557 16541 22569 16575
rect 22603 16541 22615 16575
rect 22557 16535 22615 16541
rect 22480 16504 22508 16535
rect 22646 16532 22652 16584
rect 22704 16572 22710 16584
rect 22741 16575 22799 16581
rect 22741 16572 22753 16575
rect 22704 16544 22753 16572
rect 22704 16532 22710 16544
rect 22741 16541 22753 16544
rect 22787 16541 22799 16575
rect 22741 16535 22799 16541
rect 22830 16532 22836 16584
rect 22888 16532 22894 16584
rect 22922 16532 22928 16584
rect 22980 16532 22986 16584
rect 23492 16581 23520 16612
rect 23293 16575 23351 16581
rect 23293 16541 23305 16575
rect 23339 16541 23351 16575
rect 23293 16535 23351 16541
rect 23477 16575 23535 16581
rect 23477 16541 23489 16575
rect 23523 16541 23535 16575
rect 23477 16535 23535 16541
rect 23308 16504 23336 16535
rect 23566 16532 23572 16584
rect 23624 16532 23630 16584
rect 23842 16532 23848 16584
rect 23900 16532 23906 16584
rect 24121 16575 24179 16581
rect 24121 16541 24133 16575
rect 24167 16572 24179 16575
rect 24486 16572 24492 16584
rect 24167 16544 24492 16572
rect 24167 16541 24179 16544
rect 24121 16535 24179 16541
rect 24486 16532 24492 16544
rect 24544 16532 24550 16584
rect 23661 16507 23719 16513
rect 23661 16504 23673 16507
rect 22480 16476 23244 16504
rect 23308 16476 23673 16504
rect 23216 16448 23244 16476
rect 23661 16473 23673 16476
rect 23707 16473 23719 16507
rect 23661 16467 23719 16473
rect 24673 16507 24731 16513
rect 24673 16473 24685 16507
rect 24719 16504 24731 16507
rect 24854 16504 24860 16516
rect 24719 16476 24860 16504
rect 24719 16473 24731 16476
rect 24673 16467 24731 16473
rect 24854 16464 24860 16476
rect 24912 16464 24918 16516
rect 19852 16408 19932 16436
rect 19852 16396 19858 16408
rect 19978 16396 19984 16448
rect 20036 16436 20042 16448
rect 20533 16439 20591 16445
rect 20533 16436 20545 16439
rect 20036 16408 20545 16436
rect 20036 16396 20042 16408
rect 20533 16405 20545 16408
rect 20579 16405 20591 16439
rect 20533 16399 20591 16405
rect 20898 16396 20904 16448
rect 20956 16396 20962 16448
rect 20990 16396 20996 16448
rect 21048 16436 21054 16448
rect 21269 16439 21327 16445
rect 21269 16436 21281 16439
rect 21048 16408 21281 16436
rect 21048 16396 21054 16408
rect 21269 16405 21281 16408
rect 21315 16405 21327 16439
rect 21269 16399 21327 16405
rect 22278 16396 22284 16448
rect 22336 16396 22342 16448
rect 23198 16396 23204 16448
rect 23256 16436 23262 16448
rect 24029 16439 24087 16445
rect 24029 16436 24041 16439
rect 23256 16408 24041 16436
rect 23256 16396 23262 16408
rect 24029 16405 24041 16408
rect 24075 16405 24087 16439
rect 24029 16399 24087 16405
rect 1104 16346 28152 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 28152 16346
rect 1104 16272 28152 16294
rect 2866 16192 2872 16244
rect 2924 16232 2930 16244
rect 2961 16235 3019 16241
rect 2961 16232 2973 16235
rect 2924 16204 2973 16232
rect 2924 16192 2930 16204
rect 2961 16201 2973 16204
rect 3007 16201 3019 16235
rect 2961 16195 3019 16201
rect 7469 16235 7527 16241
rect 7469 16201 7481 16235
rect 7515 16232 7527 16235
rect 7558 16232 7564 16244
rect 7515 16204 7564 16232
rect 7515 16201 7527 16204
rect 7469 16195 7527 16201
rect 7558 16192 7564 16204
rect 7616 16192 7622 16244
rect 10226 16192 10232 16244
rect 10284 16232 10290 16244
rect 10321 16235 10379 16241
rect 10321 16232 10333 16235
rect 10284 16204 10333 16232
rect 10284 16192 10290 16204
rect 10321 16201 10333 16204
rect 10367 16201 10379 16235
rect 10321 16195 10379 16201
rect 11977 16235 12035 16241
rect 11977 16201 11989 16235
rect 12023 16232 12035 16235
rect 13170 16232 13176 16244
rect 12023 16204 13176 16232
rect 12023 16201 12035 16204
rect 11977 16195 12035 16201
rect 13170 16192 13176 16204
rect 13228 16192 13234 16244
rect 14090 16192 14096 16244
rect 14148 16232 14154 16244
rect 14461 16235 14519 16241
rect 14461 16232 14473 16235
rect 14148 16204 14473 16232
rect 14148 16192 14154 16204
rect 14461 16201 14473 16204
rect 14507 16201 14519 16235
rect 14737 16235 14795 16241
rect 14737 16232 14749 16235
rect 14461 16195 14519 16201
rect 14568 16204 14749 16232
rect 3068 16136 3924 16164
rect 842 16056 848 16108
rect 900 16096 906 16108
rect 3068 16105 3096 16136
rect 1397 16099 1455 16105
rect 1397 16096 1409 16099
rect 900 16068 1409 16096
rect 900 16056 906 16068
rect 1397 16065 1409 16068
rect 1443 16065 1455 16099
rect 1397 16059 1455 16065
rect 2869 16099 2927 16105
rect 2869 16065 2881 16099
rect 2915 16065 2927 16099
rect 2869 16059 2927 16065
rect 3053 16099 3111 16105
rect 3053 16065 3065 16099
rect 3099 16065 3111 16099
rect 3053 16059 3111 16065
rect 1673 16031 1731 16037
rect 1673 15997 1685 16031
rect 1719 16028 1731 16031
rect 1854 16028 1860 16040
rect 1719 16000 1860 16028
rect 1719 15997 1731 16000
rect 1673 15991 1731 15997
rect 1854 15988 1860 16000
rect 1912 16028 1918 16040
rect 2884 16028 2912 16059
rect 3142 16056 3148 16108
rect 3200 16056 3206 16108
rect 3620 16105 3648 16136
rect 3896 16108 3924 16136
rect 7300 16136 8340 16164
rect 3605 16099 3663 16105
rect 3605 16065 3617 16099
rect 3651 16065 3663 16099
rect 3605 16059 3663 16065
rect 3789 16099 3847 16105
rect 3789 16065 3801 16099
rect 3835 16065 3847 16099
rect 3789 16059 3847 16065
rect 3160 16028 3188 16056
rect 1912 16000 3188 16028
rect 3237 16031 3295 16037
rect 1912 15988 1918 16000
rect 3237 15997 3249 16031
rect 3283 16028 3295 16031
rect 3804 16028 3832 16059
rect 3878 16056 3884 16108
rect 3936 16056 3942 16108
rect 4249 16099 4307 16105
rect 4249 16065 4261 16099
rect 4295 16065 4307 16099
rect 4249 16059 4307 16065
rect 3970 16028 3976 16040
rect 3283 16000 3976 16028
rect 3283 15997 3295 16000
rect 3237 15991 3295 15997
rect 3970 15988 3976 16000
rect 4028 16028 4034 16040
rect 4264 16028 4292 16059
rect 4614 16056 4620 16108
rect 4672 16056 4678 16108
rect 4706 16056 4712 16108
rect 4764 16096 4770 16108
rect 5169 16099 5227 16105
rect 5169 16096 5181 16099
rect 4764 16068 5181 16096
rect 4764 16056 4770 16068
rect 5169 16065 5181 16068
rect 5215 16065 5227 16099
rect 5169 16059 5227 16065
rect 5629 16099 5687 16105
rect 5629 16065 5641 16099
rect 5675 16096 5687 16099
rect 5718 16096 5724 16108
rect 5675 16068 5724 16096
rect 5675 16065 5687 16068
rect 5629 16059 5687 16065
rect 5718 16056 5724 16068
rect 5776 16056 5782 16108
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16065 5871 16099
rect 5813 16059 5871 16065
rect 6917 16099 6975 16105
rect 6917 16065 6929 16099
rect 6963 16065 6975 16099
rect 6917 16059 6975 16065
rect 4028 16000 4292 16028
rect 4028 15988 4034 16000
rect 4632 15904 4660 16056
rect 4798 15988 4804 16040
rect 4856 16028 4862 16040
rect 5828 16028 5856 16059
rect 4856 16000 5856 16028
rect 4856 15988 4862 16000
rect 6932 15960 6960 16059
rect 7190 16056 7196 16108
rect 7248 16056 7254 16108
rect 7300 16105 7328 16136
rect 8312 16108 8340 16136
rect 9968 16136 10456 16164
rect 7285 16099 7343 16105
rect 7285 16065 7297 16099
rect 7331 16065 7343 16099
rect 7285 16059 7343 16065
rect 7653 16099 7711 16105
rect 7653 16065 7665 16099
rect 7699 16096 7711 16099
rect 7834 16096 7840 16108
rect 7699 16068 7840 16096
rect 7699 16065 7711 16068
rect 7653 16059 7711 16065
rect 7208 16028 7236 16056
rect 7668 16028 7696 16059
rect 7834 16056 7840 16068
rect 7892 16056 7898 16108
rect 8294 16056 8300 16108
rect 8352 16056 8358 16108
rect 9582 16056 9588 16108
rect 9640 16056 9646 16108
rect 9858 16056 9864 16108
rect 9916 16096 9922 16108
rect 9968 16105 9996 16136
rect 10428 16105 10456 16136
rect 11790 16124 11796 16176
rect 11848 16164 11854 16176
rect 12621 16167 12679 16173
rect 11848 16136 12296 16164
rect 11848 16124 11854 16136
rect 9953 16099 10011 16105
rect 9953 16096 9965 16099
rect 9916 16068 9965 16096
rect 9916 16056 9922 16068
rect 9953 16065 9965 16068
rect 9999 16065 10011 16099
rect 9953 16059 10011 16065
rect 10229 16099 10287 16105
rect 10229 16065 10241 16099
rect 10275 16065 10287 16099
rect 10229 16059 10287 16065
rect 10413 16099 10471 16105
rect 10413 16065 10425 16099
rect 10459 16065 10471 16099
rect 10413 16059 10471 16065
rect 7208 16000 7696 16028
rect 10042 15988 10048 16040
rect 10100 15988 10106 16040
rect 7282 15960 7288 15972
rect 6932 15932 7288 15960
rect 7282 15920 7288 15932
rect 7340 15920 7346 15972
rect 10244 15960 10272 16059
rect 11698 16056 11704 16108
rect 11756 16096 11762 16108
rect 12268 16105 12296 16136
rect 12621 16133 12633 16167
rect 12667 16164 12679 16167
rect 12710 16164 12716 16176
rect 12667 16136 12716 16164
rect 12667 16133 12679 16136
rect 12621 16127 12679 16133
rect 12710 16124 12716 16136
rect 12768 16124 12774 16176
rect 14568 16164 14596 16204
rect 14737 16201 14749 16204
rect 14783 16232 14795 16235
rect 15102 16232 15108 16244
rect 14783 16204 15108 16232
rect 14783 16201 14795 16204
rect 14737 16195 14795 16201
rect 15102 16192 15108 16204
rect 15160 16192 15166 16244
rect 17126 16192 17132 16244
rect 17184 16192 17190 16244
rect 17218 16192 17224 16244
rect 17276 16232 17282 16244
rect 17862 16232 17868 16244
rect 17276 16204 17868 16232
rect 17276 16192 17282 16204
rect 17862 16192 17868 16204
rect 17920 16192 17926 16244
rect 18046 16192 18052 16244
rect 18104 16192 18110 16244
rect 18874 16192 18880 16244
rect 18932 16232 18938 16244
rect 19610 16232 19616 16244
rect 18932 16204 19616 16232
rect 18932 16192 18938 16204
rect 19610 16192 19616 16204
rect 19668 16232 19674 16244
rect 20162 16232 20168 16244
rect 19668 16204 20168 16232
rect 19668 16192 19674 16204
rect 20162 16192 20168 16204
rect 20220 16192 20226 16244
rect 23198 16192 23204 16244
rect 23256 16192 23262 16244
rect 24026 16192 24032 16244
rect 24084 16192 24090 16244
rect 18064 16164 18092 16192
rect 19886 16164 19892 16176
rect 14108 16136 14596 16164
rect 14660 16136 18092 16164
rect 18156 16136 19012 16164
rect 12161 16099 12219 16105
rect 12161 16096 12173 16099
rect 11756 16068 12173 16096
rect 11756 16056 11762 16068
rect 12161 16065 12173 16068
rect 12207 16065 12219 16099
rect 12161 16059 12219 16065
rect 12253 16099 12311 16105
rect 12253 16065 12265 16099
rect 12299 16065 12311 16099
rect 12253 16059 12311 16065
rect 12529 16099 12587 16105
rect 12529 16065 12541 16099
rect 12575 16096 12587 16099
rect 13814 16096 13820 16108
rect 12575 16068 13820 16096
rect 12575 16065 12587 16068
rect 12529 16059 12587 16065
rect 13814 16056 13820 16068
rect 13872 16056 13878 16108
rect 10594 15988 10600 16040
rect 10652 16028 10658 16040
rect 14108 16028 14136 16136
rect 14458 16056 14464 16108
rect 14516 16096 14522 16108
rect 14660 16105 14688 16136
rect 14553 16099 14611 16105
rect 14553 16096 14565 16099
rect 14516 16068 14565 16096
rect 14516 16056 14522 16068
rect 14553 16065 14565 16068
rect 14599 16065 14611 16099
rect 14553 16059 14611 16065
rect 14645 16099 14703 16105
rect 14645 16065 14657 16099
rect 14691 16065 14703 16099
rect 14645 16059 14703 16065
rect 14921 16099 14979 16105
rect 14921 16065 14933 16099
rect 14967 16096 14979 16099
rect 15010 16096 15016 16108
rect 14967 16068 15016 16096
rect 14967 16065 14979 16068
rect 14921 16059 14979 16065
rect 15010 16056 15016 16068
rect 15068 16056 15074 16108
rect 15381 16099 15439 16105
rect 15381 16065 15393 16099
rect 15427 16096 15439 16099
rect 16669 16099 16727 16105
rect 16669 16096 16681 16099
rect 15427 16068 16681 16096
rect 15427 16065 15439 16068
rect 15381 16059 15439 16065
rect 16669 16065 16681 16068
rect 16715 16065 16727 16099
rect 16669 16059 16727 16065
rect 16945 16099 17003 16105
rect 16945 16065 16957 16099
rect 16991 16096 17003 16099
rect 17218 16096 17224 16108
rect 16991 16068 17224 16096
rect 16991 16065 17003 16068
rect 16945 16059 17003 16065
rect 17218 16056 17224 16068
rect 17276 16056 17282 16108
rect 17402 16056 17408 16108
rect 17460 16056 17466 16108
rect 17865 16099 17923 16105
rect 17865 16065 17877 16099
rect 17911 16065 17923 16099
rect 17865 16059 17923 16065
rect 10652 16000 14136 16028
rect 14185 16031 14243 16037
rect 10652 15988 10658 16000
rect 14185 15997 14197 16031
rect 14231 16028 14243 16031
rect 15194 16028 15200 16040
rect 14231 16000 15200 16028
rect 14231 15997 14243 16000
rect 14185 15991 14243 15997
rect 15194 15988 15200 16000
rect 15252 15988 15258 16040
rect 16853 16031 16911 16037
rect 16853 15997 16865 16031
rect 16899 16028 16911 16031
rect 17770 16028 17776 16040
rect 16899 16000 17776 16028
rect 16899 15997 16911 16000
rect 16853 15991 16911 15997
rect 17770 15988 17776 16000
rect 17828 15988 17834 16040
rect 9324 15932 10272 15960
rect 9324 15904 9352 15932
rect 13998 15920 14004 15972
rect 14056 15960 14062 15972
rect 15013 15963 15071 15969
rect 15013 15960 15025 15963
rect 14056 15932 15025 15960
rect 14056 15920 14062 15932
rect 15013 15929 15025 15932
rect 15059 15929 15071 15963
rect 15013 15923 15071 15929
rect 16942 15920 16948 15972
rect 17000 15960 17006 15972
rect 17126 15960 17132 15972
rect 17000 15932 17132 15960
rect 17000 15920 17006 15932
rect 17126 15920 17132 15932
rect 17184 15960 17190 15972
rect 17681 15963 17739 15969
rect 17681 15960 17693 15963
rect 17184 15932 17693 15960
rect 17184 15920 17190 15932
rect 17681 15929 17693 15932
rect 17727 15929 17739 15963
rect 17880 15960 17908 16059
rect 18046 16056 18052 16108
rect 18104 16056 18110 16108
rect 18156 16105 18184 16136
rect 18141 16099 18199 16105
rect 18141 16065 18153 16099
rect 18187 16065 18199 16099
rect 18141 16059 18199 16065
rect 18874 16056 18880 16108
rect 18932 16056 18938 16108
rect 18984 16096 19012 16136
rect 19306 16136 19892 16164
rect 19306 16096 19334 16136
rect 19886 16124 19892 16136
rect 19944 16124 19950 16176
rect 22278 16124 22284 16176
rect 22336 16164 22342 16176
rect 23661 16167 23719 16173
rect 23661 16164 23673 16167
rect 22336 16136 23673 16164
rect 22336 16124 22342 16136
rect 23661 16133 23673 16136
rect 23707 16133 23719 16167
rect 24044 16164 24072 16192
rect 24044 16136 24150 16164
rect 23661 16127 23719 16133
rect 18984 16068 19334 16096
rect 19521 16099 19579 16105
rect 19521 16065 19533 16099
rect 19567 16065 19579 16099
rect 19521 16059 19579 16065
rect 19797 16099 19855 16105
rect 19797 16065 19809 16099
rect 19843 16096 19855 16099
rect 20898 16096 20904 16108
rect 19843 16068 20904 16096
rect 19843 16065 19855 16068
rect 19797 16059 19855 16065
rect 18064 16028 18092 16056
rect 18785 16031 18843 16037
rect 18785 16028 18797 16031
rect 18064 16000 18797 16028
rect 18785 15997 18797 16000
rect 18831 15997 18843 16031
rect 18785 15991 18843 15997
rect 19536 16028 19564 16059
rect 20898 16056 20904 16068
rect 20956 16056 20962 16108
rect 23293 16099 23351 16105
rect 23293 16065 23305 16099
rect 23339 16065 23351 16099
rect 23293 16059 23351 16065
rect 20438 16028 20444 16040
rect 19536 16000 20444 16028
rect 19334 15960 19340 15972
rect 17880 15932 19340 15960
rect 17681 15923 17739 15929
rect 19334 15920 19340 15932
rect 19392 15920 19398 15972
rect 3786 15852 3792 15904
rect 3844 15852 3850 15904
rect 4614 15852 4620 15904
rect 4672 15852 4678 15904
rect 5718 15852 5724 15904
rect 5776 15852 5782 15904
rect 7009 15895 7067 15901
rect 7009 15861 7021 15895
rect 7055 15892 7067 15895
rect 8110 15892 8116 15904
rect 7055 15864 8116 15892
rect 7055 15861 7067 15864
rect 7009 15855 7067 15861
rect 8110 15852 8116 15864
rect 8168 15852 8174 15904
rect 9306 15852 9312 15904
rect 9364 15852 9370 15904
rect 9674 15852 9680 15904
rect 9732 15852 9738 15904
rect 13814 15852 13820 15904
rect 13872 15852 13878 15904
rect 14090 15852 14096 15904
rect 14148 15852 14154 15904
rect 14274 15852 14280 15904
rect 14332 15852 14338 15904
rect 15102 15852 15108 15904
rect 15160 15852 15166 15904
rect 16666 15852 16672 15904
rect 16724 15852 16730 15904
rect 17218 15852 17224 15904
rect 17276 15892 17282 15904
rect 17313 15895 17371 15901
rect 17313 15892 17325 15895
rect 17276 15864 17325 15892
rect 17276 15852 17282 15864
rect 17313 15861 17325 15864
rect 17359 15861 17371 15895
rect 17313 15855 17371 15861
rect 17402 15852 17408 15904
rect 17460 15892 17466 15904
rect 19536 15892 19564 16000
rect 20438 15988 20444 16000
rect 20496 16028 20502 16040
rect 21082 16028 21088 16040
rect 20496 16000 21088 16028
rect 20496 15988 20502 16000
rect 21082 15988 21088 16000
rect 21140 15988 21146 16040
rect 21634 15988 21640 16040
rect 21692 16028 21698 16040
rect 23308 16028 23336 16059
rect 23382 16056 23388 16108
rect 23440 16056 23446 16108
rect 23750 16028 23756 16040
rect 21692 16000 23756 16028
rect 21692 15988 21698 16000
rect 23750 15988 23756 16000
rect 23808 16028 23814 16040
rect 25133 16031 25191 16037
rect 25133 16028 25145 16031
rect 23808 16000 25145 16028
rect 23808 15988 23814 16000
rect 25133 15997 25145 16000
rect 25179 15997 25191 16031
rect 25133 15991 25191 15997
rect 17460 15864 19564 15892
rect 19981 15895 20039 15901
rect 17460 15852 17466 15864
rect 19981 15861 19993 15895
rect 20027 15892 20039 15895
rect 20254 15892 20260 15904
rect 20027 15864 20260 15892
rect 20027 15861 20039 15864
rect 19981 15855 20039 15861
rect 20254 15852 20260 15864
rect 20312 15852 20318 15904
rect 1104 15802 28152 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 28152 15802
rect 1104 15728 28152 15750
rect 12158 15648 12164 15700
rect 12216 15648 12222 15700
rect 13814 15648 13820 15700
rect 13872 15688 13878 15700
rect 16117 15691 16175 15697
rect 16117 15688 16129 15691
rect 13872 15660 16129 15688
rect 13872 15648 13878 15660
rect 16117 15657 16129 15660
rect 16163 15657 16175 15691
rect 16117 15651 16175 15657
rect 16577 15691 16635 15697
rect 16577 15657 16589 15691
rect 16623 15688 16635 15691
rect 16850 15688 16856 15700
rect 16623 15660 16856 15688
rect 16623 15657 16635 15660
rect 16577 15651 16635 15657
rect 16850 15648 16856 15660
rect 16908 15648 16914 15700
rect 18690 15648 18696 15700
rect 18748 15688 18754 15700
rect 22830 15688 22836 15700
rect 18748 15660 22836 15688
rect 18748 15648 18754 15660
rect 22830 15648 22836 15660
rect 22888 15648 22894 15700
rect 23566 15648 23572 15700
rect 23624 15688 23630 15700
rect 23937 15691 23995 15697
rect 23937 15688 23949 15691
rect 23624 15660 23949 15688
rect 23624 15648 23630 15660
rect 23937 15657 23949 15660
rect 23983 15657 23995 15691
rect 23937 15651 23995 15657
rect 24581 15691 24639 15697
rect 24581 15657 24593 15691
rect 24627 15688 24639 15691
rect 24762 15688 24768 15700
rect 24627 15660 24768 15688
rect 24627 15657 24639 15660
rect 24581 15651 24639 15657
rect 24762 15648 24768 15660
rect 24820 15648 24826 15700
rect 16942 15580 16948 15632
rect 17000 15580 17006 15632
rect 19610 15620 19616 15632
rect 19076 15592 19616 15620
rect 4433 15555 4491 15561
rect 4433 15521 4445 15555
rect 4479 15552 4491 15555
rect 4614 15552 4620 15564
rect 4479 15524 4620 15552
rect 4479 15521 4491 15524
rect 4433 15515 4491 15521
rect 4614 15512 4620 15524
rect 4672 15512 4678 15564
rect 13354 15512 13360 15564
rect 13412 15552 13418 15564
rect 16209 15555 16267 15561
rect 16209 15552 16221 15555
rect 13412 15524 16221 15552
rect 13412 15512 13418 15524
rect 16209 15521 16221 15524
rect 16255 15521 16267 15555
rect 16209 15515 16267 15521
rect 3786 15444 3792 15496
rect 3844 15484 3850 15496
rect 4341 15487 4399 15493
rect 4341 15484 4353 15487
rect 3844 15456 4353 15484
rect 3844 15444 3850 15456
rect 4341 15453 4353 15456
rect 4387 15453 4399 15487
rect 4341 15447 4399 15453
rect 7282 15444 7288 15496
rect 7340 15444 7346 15496
rect 8110 15444 8116 15496
rect 8168 15444 8174 15496
rect 9306 15444 9312 15496
rect 9364 15444 9370 15496
rect 9674 15444 9680 15496
rect 9732 15484 9738 15496
rect 9769 15487 9827 15493
rect 9769 15484 9781 15487
rect 9732 15456 9781 15484
rect 9732 15444 9738 15456
rect 9769 15453 9781 15456
rect 9815 15453 9827 15487
rect 9769 15447 9827 15453
rect 10502 15444 10508 15496
rect 10560 15484 10566 15496
rect 11609 15487 11667 15493
rect 10560 15456 11376 15484
rect 10560 15444 10566 15456
rect 8757 15419 8815 15425
rect 8757 15385 8769 15419
rect 8803 15416 8815 15419
rect 9858 15416 9864 15428
rect 8803 15388 9864 15416
rect 8803 15385 8815 15388
rect 8757 15379 8815 15385
rect 9858 15376 9864 15388
rect 9916 15376 9922 15428
rect 11348 15416 11376 15456
rect 11609 15453 11621 15487
rect 11655 15484 11667 15487
rect 11698 15484 11704 15496
rect 11655 15456 11704 15484
rect 11655 15453 11667 15456
rect 11609 15447 11667 15453
rect 11698 15444 11704 15456
rect 11756 15444 11762 15496
rect 11790 15444 11796 15496
rect 11848 15444 11854 15496
rect 11974 15444 11980 15496
rect 12032 15444 12038 15496
rect 16393 15487 16451 15493
rect 16393 15453 16405 15487
rect 16439 15484 16451 15487
rect 16574 15484 16580 15496
rect 16439 15456 16580 15484
rect 16439 15453 16451 15456
rect 16393 15447 16451 15453
rect 16574 15444 16580 15456
rect 16632 15444 16638 15496
rect 16758 15444 16764 15496
rect 16816 15444 16822 15496
rect 16960 15493 16988 15580
rect 17034 15512 17040 15564
rect 17092 15512 17098 15564
rect 19076 15561 19104 15592
rect 19610 15580 19616 15592
rect 19668 15580 19674 15632
rect 23198 15580 23204 15632
rect 23256 15620 23262 15632
rect 23385 15623 23443 15629
rect 23385 15620 23397 15623
rect 23256 15592 23397 15620
rect 23256 15580 23262 15592
rect 23385 15589 23397 15592
rect 23431 15589 23443 15623
rect 23385 15583 23443 15589
rect 23474 15580 23480 15632
rect 23532 15620 23538 15632
rect 24397 15623 24455 15629
rect 24397 15620 24409 15623
rect 23532 15592 24409 15620
rect 23532 15580 23538 15592
rect 24397 15589 24409 15592
rect 24443 15589 24455 15623
rect 24397 15583 24455 15589
rect 19061 15555 19119 15561
rect 19061 15521 19073 15555
rect 19107 15521 19119 15555
rect 19061 15515 19119 15521
rect 20254 15512 20260 15564
rect 20312 15512 20318 15564
rect 20714 15512 20720 15564
rect 20772 15552 20778 15564
rect 21450 15552 21456 15564
rect 20772 15524 21456 15552
rect 20772 15512 20778 15524
rect 16945 15487 17003 15493
rect 16945 15453 16957 15487
rect 16991 15453 17003 15487
rect 16945 15447 17003 15453
rect 19978 15444 19984 15496
rect 20036 15444 20042 15496
rect 20165 15487 20223 15493
rect 20165 15453 20177 15487
rect 20211 15484 20223 15487
rect 20806 15484 20812 15496
rect 20211 15456 20812 15484
rect 20211 15453 20223 15456
rect 20165 15447 20223 15453
rect 20806 15444 20812 15456
rect 20864 15444 20870 15496
rect 20916 15493 20944 15524
rect 21450 15512 21456 15524
rect 21508 15512 21514 15564
rect 24854 15552 24860 15564
rect 22066 15524 24860 15552
rect 20901 15487 20959 15493
rect 20901 15453 20913 15487
rect 20947 15453 20959 15487
rect 20901 15447 20959 15453
rect 21085 15487 21143 15493
rect 21085 15453 21097 15487
rect 21131 15484 21143 15487
rect 21634 15484 21640 15496
rect 21131 15456 21640 15484
rect 21131 15453 21143 15456
rect 21085 15447 21143 15453
rect 21634 15444 21640 15456
rect 21692 15444 21698 15496
rect 11885 15419 11943 15425
rect 11885 15416 11897 15419
rect 10718 15388 11284 15416
rect 11348 15388 11897 15416
rect 4706 15308 4712 15360
rect 4764 15308 4770 15360
rect 11256 15348 11284 15388
rect 11885 15385 11897 15388
rect 11931 15385 11943 15419
rect 16117 15419 16175 15425
rect 11885 15379 11943 15385
rect 11992 15388 12434 15416
rect 11992 15348 12020 15388
rect 11256 15320 12020 15348
rect 12406 15348 12434 15388
rect 16117 15385 16129 15419
rect 16163 15416 16175 15419
rect 16853 15419 16911 15425
rect 16163 15388 16804 15416
rect 16163 15385 16175 15388
rect 16117 15379 16175 15385
rect 16776 15360 16804 15388
rect 16853 15385 16865 15419
rect 16899 15416 16911 15419
rect 17313 15419 17371 15425
rect 17313 15416 17325 15419
rect 16899 15388 17325 15416
rect 16899 15385 16911 15388
rect 16853 15379 16911 15385
rect 17313 15385 17325 15388
rect 17359 15385 17371 15419
rect 19518 15416 19524 15428
rect 18538 15388 19524 15416
rect 17313 15379 17371 15385
rect 19518 15376 19524 15388
rect 19576 15416 19582 15428
rect 20346 15416 20352 15428
rect 19576 15388 20352 15416
rect 19576 15376 19582 15388
rect 20346 15376 20352 15388
rect 20404 15416 20410 15428
rect 22066 15416 22094 15524
rect 24854 15512 24860 15524
rect 24912 15512 24918 15564
rect 23106 15444 23112 15496
rect 23164 15484 23170 15496
rect 23201 15487 23259 15493
rect 23201 15484 23213 15487
rect 23164 15456 23213 15484
rect 23164 15444 23170 15456
rect 23201 15453 23213 15456
rect 23247 15453 23259 15487
rect 23201 15447 23259 15453
rect 23566 15444 23572 15496
rect 23624 15444 23630 15496
rect 23661 15487 23719 15493
rect 23661 15453 23673 15487
rect 23707 15484 23719 15487
rect 24210 15484 24216 15496
rect 23707 15456 24216 15484
rect 23707 15453 23719 15456
rect 23661 15447 23719 15453
rect 24210 15444 24216 15456
rect 24268 15444 24274 15496
rect 20404 15388 22094 15416
rect 20404 15376 20410 15388
rect 23750 15376 23756 15428
rect 23808 15416 23814 15428
rect 24765 15419 24823 15425
rect 24765 15416 24777 15419
rect 23808 15388 24777 15416
rect 23808 15376 23814 15388
rect 24765 15385 24777 15388
rect 24811 15385 24823 15419
rect 24765 15379 24823 15385
rect 16022 15348 16028 15360
rect 12406 15320 16028 15348
rect 16022 15308 16028 15320
rect 16080 15308 16086 15360
rect 16758 15308 16764 15360
rect 16816 15308 16822 15360
rect 19794 15308 19800 15360
rect 19852 15308 19858 15360
rect 21082 15308 21088 15360
rect 21140 15308 21146 15360
rect 24026 15308 24032 15360
rect 24084 15348 24090 15360
rect 24555 15351 24613 15357
rect 24555 15348 24567 15351
rect 24084 15320 24567 15348
rect 24084 15308 24090 15320
rect 24555 15317 24567 15320
rect 24601 15317 24613 15351
rect 24555 15311 24613 15317
rect 1104 15258 28152 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 28152 15258
rect 1104 15184 28152 15206
rect 7282 15104 7288 15156
rect 7340 15144 7346 15156
rect 8573 15147 8631 15153
rect 7340 15116 8432 15144
rect 7340 15104 7346 15116
rect 3436 15048 4384 15076
rect 2406 14968 2412 15020
rect 2464 15008 2470 15020
rect 2501 15011 2559 15017
rect 2501 15008 2513 15011
rect 2464 14980 2513 15008
rect 2464 14968 2470 14980
rect 2501 14977 2513 14980
rect 2547 14977 2559 15011
rect 2501 14971 2559 14977
rect 2682 14968 2688 15020
rect 2740 14968 2746 15020
rect 3326 14968 3332 15020
rect 3384 15008 3390 15020
rect 3436 15017 3464 15048
rect 3421 15011 3479 15017
rect 3421 15008 3433 15011
rect 3384 14980 3433 15008
rect 3384 14968 3390 14980
rect 3421 14977 3433 14980
rect 3467 14977 3479 15011
rect 3421 14971 3479 14977
rect 3510 14968 3516 15020
rect 3568 15008 3574 15020
rect 4356 15017 4384 15048
rect 8110 15036 8116 15088
rect 8168 15076 8174 15088
rect 8404 15085 8432 15116
rect 8573 15113 8585 15147
rect 8619 15144 8631 15147
rect 9582 15144 9588 15156
rect 8619 15116 9588 15144
rect 8619 15113 8631 15116
rect 8573 15107 8631 15113
rect 9582 15104 9588 15116
rect 9640 15104 9646 15156
rect 12066 15104 12072 15156
rect 12124 15104 12130 15156
rect 12342 15104 12348 15156
rect 12400 15104 12406 15156
rect 14185 15147 14243 15153
rect 14185 15113 14197 15147
rect 14231 15144 14243 15147
rect 14274 15144 14280 15156
rect 14231 15116 14280 15144
rect 14231 15113 14243 15116
rect 14185 15107 14243 15113
rect 14274 15104 14280 15116
rect 14332 15104 14338 15156
rect 16758 15104 16764 15156
rect 16816 15144 16822 15156
rect 16853 15147 16911 15153
rect 16853 15144 16865 15147
rect 16816 15116 16865 15144
rect 16816 15104 16822 15116
rect 16853 15113 16865 15116
rect 16899 15113 16911 15147
rect 16853 15107 16911 15113
rect 16942 15104 16948 15156
rect 17000 15144 17006 15156
rect 17405 15147 17463 15153
rect 17405 15144 17417 15147
rect 17000 15116 17417 15144
rect 17000 15104 17006 15116
rect 17405 15113 17417 15116
rect 17451 15113 17463 15147
rect 17405 15107 17463 15113
rect 20806 15104 20812 15156
rect 20864 15104 20870 15156
rect 23382 15104 23388 15156
rect 23440 15144 23446 15156
rect 23842 15144 23848 15156
rect 23440 15116 23848 15144
rect 23440 15104 23446 15116
rect 23842 15104 23848 15116
rect 23900 15104 23906 15156
rect 10692 15088 10744 15094
rect 8205 15079 8263 15085
rect 8205 15076 8217 15079
rect 8168 15048 8217 15076
rect 8168 15036 8174 15048
rect 8205 15045 8217 15048
rect 8251 15045 8263 15079
rect 8205 15039 8263 15045
rect 8389 15079 8447 15085
rect 8389 15045 8401 15079
rect 8435 15045 8447 15079
rect 8389 15039 8447 15045
rect 9033 15079 9091 15085
rect 9033 15045 9045 15079
rect 9079 15076 9091 15079
rect 9079 15048 10088 15076
rect 9079 15045 9091 15048
rect 9033 15039 9091 15045
rect 10060 15020 10088 15048
rect 12084 15076 12112 15104
rect 12084 15048 12756 15076
rect 10692 15030 10744 15036
rect 4157 15011 4215 15017
rect 4157 15008 4169 15011
rect 3568 14980 4169 15008
rect 3568 14968 3574 14980
rect 4157 14977 4169 14980
rect 4203 14977 4215 15011
rect 4157 14971 4215 14977
rect 4341 15011 4399 15017
rect 4341 14977 4353 15011
rect 4387 14977 4399 15011
rect 4341 14971 4399 14977
rect 4706 14968 4712 15020
rect 4764 15008 4770 15020
rect 5077 15011 5135 15017
rect 5077 15008 5089 15011
rect 4764 14980 5089 15008
rect 4764 14968 4770 14980
rect 5077 14977 5089 14980
rect 5123 14977 5135 15011
rect 5077 14971 5135 14977
rect 5258 14968 5264 15020
rect 5316 14968 5322 15020
rect 5718 14968 5724 15020
rect 5776 15008 5782 15020
rect 6365 15011 6423 15017
rect 6365 15008 6377 15011
rect 5776 14980 6377 15008
rect 5776 14968 5782 14980
rect 6365 14977 6377 14980
rect 6411 14977 6423 15011
rect 6365 14971 6423 14977
rect 7285 15011 7343 15017
rect 7285 14977 7297 15011
rect 7331 15008 7343 15011
rect 7374 15008 7380 15020
rect 7331 14980 7380 15008
rect 7331 14977 7343 14980
rect 7285 14971 7343 14977
rect 7374 14968 7380 14980
rect 7432 14968 7438 15020
rect 7466 14968 7472 15020
rect 7524 14968 7530 15020
rect 8662 14968 8668 15020
rect 8720 14968 8726 15020
rect 8849 15011 8907 15017
rect 8849 14977 8861 15011
rect 8895 14977 8907 15011
rect 8849 14971 8907 14977
rect 4062 14900 4068 14952
rect 4120 14900 4126 14952
rect 6089 14943 6147 14949
rect 6089 14909 6101 14943
rect 6135 14940 6147 14943
rect 6822 14940 6828 14952
rect 6135 14912 6828 14940
rect 6135 14909 6147 14912
rect 6089 14903 6147 14909
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 6733 14875 6791 14881
rect 6733 14841 6745 14875
rect 6779 14872 6791 14875
rect 7190 14872 7196 14884
rect 6779 14844 7196 14872
rect 6779 14841 6791 14844
rect 6733 14835 6791 14841
rect 7190 14832 7196 14844
rect 7248 14832 7254 14884
rect 7392 14872 7420 14968
rect 8570 14900 8576 14952
rect 8628 14940 8634 14952
rect 8864 14940 8892 14971
rect 9858 14968 9864 15020
rect 9916 14968 9922 15020
rect 10042 14968 10048 15020
rect 10100 15008 10106 15020
rect 10321 15011 10379 15017
rect 10321 15008 10333 15011
rect 10100 14980 10333 15008
rect 10100 14968 10106 14980
rect 10321 14977 10333 14980
rect 10367 14977 10379 15011
rect 10321 14971 10379 14977
rect 11790 14968 11796 15020
rect 11848 14968 11854 15020
rect 11977 15011 12035 15017
rect 11977 14977 11989 15011
rect 12023 14977 12035 15011
rect 11977 14971 12035 14977
rect 8628 14912 8892 14940
rect 8628 14900 8634 14912
rect 7926 14872 7932 14884
rect 7392 14844 7932 14872
rect 7926 14832 7932 14844
rect 7984 14872 7990 14884
rect 10502 14872 10508 14884
rect 7984 14844 10508 14872
rect 7984 14832 7990 14844
rect 10502 14832 10508 14844
rect 10560 14832 10566 14884
rect 11992 14872 12020 14971
rect 12066 14968 12072 15020
rect 12124 14968 12130 15020
rect 12161 15011 12219 15017
rect 12161 14977 12173 15011
rect 12207 14977 12219 15011
rect 12161 14971 12219 14977
rect 12066 14872 12072 14884
rect 11992 14844 12072 14872
rect 12066 14832 12072 14844
rect 12124 14832 12130 14884
rect 2685 14807 2743 14813
rect 2685 14773 2697 14807
rect 2731 14804 2743 14807
rect 2866 14804 2872 14816
rect 2731 14776 2872 14804
rect 2731 14773 2743 14776
rect 2685 14767 2743 14773
rect 2866 14764 2872 14776
rect 2924 14764 2930 14816
rect 3878 14764 3884 14816
rect 3936 14804 3942 14816
rect 4249 14807 4307 14813
rect 4249 14804 4261 14807
rect 3936 14776 4261 14804
rect 3936 14764 3942 14776
rect 4249 14773 4261 14776
rect 4295 14773 4307 14807
rect 4249 14767 4307 14773
rect 11330 14764 11336 14816
rect 11388 14804 11394 14816
rect 12176 14804 12204 14971
rect 12434 14968 12440 15020
rect 12492 15008 12498 15020
rect 12728 15017 12756 15048
rect 14366 15036 14372 15088
rect 14424 15076 14430 15088
rect 18046 15076 18052 15088
rect 14424 15048 14596 15076
rect 14424 15036 14430 15048
rect 12621 15011 12679 15017
rect 12621 15008 12633 15011
rect 12492 14980 12633 15008
rect 12492 14968 12498 14980
rect 12621 14977 12633 14980
rect 12667 14977 12679 15011
rect 12621 14971 12679 14977
rect 12713 15011 12771 15017
rect 12713 14977 12725 15011
rect 12759 14977 12771 15011
rect 12713 14971 12771 14977
rect 12894 14968 12900 15020
rect 12952 14968 12958 15020
rect 12989 15011 13047 15017
rect 12989 14977 13001 15011
rect 13035 15008 13047 15011
rect 13354 15008 13360 15020
rect 13035 14980 13360 15008
rect 13035 14977 13047 14980
rect 12989 14971 13047 14977
rect 13354 14968 13360 14980
rect 13412 14968 13418 15020
rect 14274 14968 14280 15020
rect 14332 14968 14338 15020
rect 14568 15017 14596 15048
rect 17604 15048 18052 15076
rect 14553 15011 14611 15017
rect 14553 14977 14565 15011
rect 14599 15008 14611 15011
rect 14826 15008 14832 15020
rect 14599 14980 14832 15008
rect 14599 14977 14611 14980
rect 14553 14971 14611 14977
rect 14826 14968 14832 14980
rect 14884 14968 14890 15020
rect 17034 14968 17040 15020
rect 17092 14968 17098 15020
rect 17604 15017 17632 15048
rect 18046 15036 18052 15048
rect 18104 15036 18110 15088
rect 20622 15076 20628 15088
rect 18156 15048 20628 15076
rect 18156 15020 18184 15048
rect 20622 15036 20628 15048
rect 20680 15036 20686 15088
rect 20717 15079 20775 15085
rect 20717 15045 20729 15079
rect 20763 15076 20775 15079
rect 22186 15076 22192 15088
rect 20763 15048 21128 15076
rect 20763 15045 20775 15048
rect 20717 15039 20775 15045
rect 21100 15020 21128 15048
rect 21468 15048 22192 15076
rect 21468 15020 21496 15048
rect 22186 15036 22192 15048
rect 22244 15036 22250 15088
rect 23750 15036 23756 15088
rect 23808 15036 23814 15088
rect 17313 15011 17371 15017
rect 17313 15008 17325 15011
rect 17144 14980 17325 15008
rect 14182 14900 14188 14952
rect 14240 14900 14246 14952
rect 14369 14943 14427 14949
rect 14369 14909 14381 14943
rect 14415 14940 14427 14943
rect 14458 14940 14464 14952
rect 14415 14912 14464 14940
rect 14415 14909 14427 14912
rect 14369 14903 14427 14909
rect 14458 14900 14464 14912
rect 14516 14900 14522 14952
rect 14645 14943 14703 14949
rect 14645 14909 14657 14943
rect 14691 14940 14703 14943
rect 14734 14940 14740 14952
rect 14691 14912 14740 14940
rect 14691 14909 14703 14912
rect 14645 14903 14703 14909
rect 14734 14900 14740 14912
rect 14792 14940 14798 14952
rect 15010 14940 15016 14952
rect 14792 14912 15016 14940
rect 14792 14900 14798 14912
rect 15010 14900 15016 14912
rect 15068 14900 15074 14952
rect 15286 14900 15292 14952
rect 15344 14940 15350 14952
rect 17144 14940 17172 14980
rect 17313 14977 17325 14980
rect 17359 14977 17371 15011
rect 17313 14971 17371 14977
rect 17589 15011 17647 15017
rect 17589 14977 17601 15011
rect 17635 14977 17647 15011
rect 17589 14971 17647 14977
rect 17957 15011 18015 15017
rect 17957 14977 17969 15011
rect 18003 14977 18015 15011
rect 17957 14971 18015 14977
rect 15344 14912 17172 14940
rect 17221 14943 17279 14949
rect 15344 14900 15350 14912
rect 17221 14909 17233 14943
rect 17267 14940 17279 14943
rect 17402 14940 17408 14952
rect 17267 14912 17408 14940
rect 17267 14909 17279 14912
rect 17221 14903 17279 14909
rect 17402 14900 17408 14912
rect 17460 14900 17466 14952
rect 17770 14900 17776 14952
rect 17828 14900 17834 14952
rect 17865 14943 17923 14949
rect 17865 14909 17877 14943
rect 17911 14909 17923 14943
rect 17972 14940 18000 14971
rect 18138 14968 18144 15020
rect 18196 14968 18202 15020
rect 19978 14968 19984 15020
rect 20036 14968 20042 15020
rect 20254 14968 20260 15020
rect 20312 14968 20318 15020
rect 20898 15008 20904 15020
rect 20364 14980 20904 15008
rect 20364 14940 20392 14980
rect 20898 14968 20904 14980
rect 20956 14968 20962 15020
rect 20990 14968 20996 15020
rect 21048 14968 21054 15020
rect 21082 14968 21088 15020
rect 21140 15008 21146 15020
rect 21269 15011 21327 15017
rect 21269 15008 21281 15011
rect 21140 14980 21281 15008
rect 21140 14968 21146 14980
rect 21269 14977 21281 14980
rect 21315 14977 21327 15011
rect 21269 14971 21327 14977
rect 21450 14968 21456 15020
rect 21508 14968 21514 15020
rect 21634 14968 21640 15020
rect 21692 14968 21698 15020
rect 22370 14968 22376 15020
rect 22428 15008 22434 15020
rect 23109 15011 23167 15017
rect 23109 15008 23121 15011
rect 22428 14980 23121 15008
rect 22428 14968 22434 14980
rect 23109 14977 23121 14980
rect 23155 14977 23167 15011
rect 23109 14971 23167 14977
rect 23934 14968 23940 15020
rect 23992 14968 23998 15020
rect 24026 14968 24032 15020
rect 24084 14968 24090 15020
rect 17972 14912 20392 14940
rect 20441 14943 20499 14949
rect 17865 14903 17923 14909
rect 20441 14909 20453 14943
rect 20487 14940 20499 14943
rect 20622 14940 20628 14952
rect 20487 14912 20628 14940
rect 20487 14909 20499 14912
rect 20441 14903 20499 14909
rect 17586 14832 17592 14884
rect 17644 14872 17650 14884
rect 17880 14872 17908 14903
rect 20622 14900 20628 14912
rect 20680 14900 20686 14952
rect 20714 14900 20720 14952
rect 20772 14940 20778 14952
rect 24210 14940 24216 14952
rect 20772 14912 24216 14940
rect 20772 14900 20778 14912
rect 24210 14900 24216 14912
rect 24268 14900 24274 14952
rect 18782 14872 18788 14884
rect 17644 14844 18788 14872
rect 17644 14832 17650 14844
rect 18782 14832 18788 14844
rect 18840 14832 18846 14884
rect 21085 14875 21143 14881
rect 21085 14872 21097 14875
rect 20640 14844 21097 14872
rect 11388 14776 12204 14804
rect 11388 14764 11394 14776
rect 12250 14764 12256 14816
rect 12308 14804 12314 14816
rect 12437 14807 12495 14813
rect 12437 14804 12449 14807
rect 12308 14776 12449 14804
rect 12308 14764 12314 14776
rect 12437 14773 12449 14776
rect 12483 14773 12495 14807
rect 12437 14767 12495 14773
rect 14918 14764 14924 14816
rect 14976 14804 14982 14816
rect 16942 14804 16948 14816
rect 14976 14776 16948 14804
rect 14976 14764 14982 14776
rect 16942 14764 16948 14776
rect 17000 14764 17006 14816
rect 17310 14764 17316 14816
rect 17368 14764 17374 14816
rect 18693 14807 18751 14813
rect 18693 14773 18705 14807
rect 18739 14804 18751 14807
rect 19702 14804 19708 14816
rect 18739 14776 19708 14804
rect 18739 14773 18751 14776
rect 18693 14767 18751 14773
rect 19702 14764 19708 14776
rect 19760 14764 19766 14816
rect 20070 14764 20076 14816
rect 20128 14764 20134 14816
rect 20640 14813 20668 14844
rect 21085 14841 21097 14844
rect 21131 14841 21143 14875
rect 21085 14835 21143 14841
rect 20625 14807 20683 14813
rect 20625 14773 20637 14807
rect 20671 14773 20683 14807
rect 21100 14804 21128 14835
rect 21174 14832 21180 14884
rect 21232 14832 21238 14884
rect 21818 14832 21824 14884
rect 21876 14872 21882 14884
rect 23290 14872 23296 14884
rect 21876 14844 23296 14872
rect 21876 14832 21882 14844
rect 23290 14832 23296 14844
rect 23348 14832 23354 14884
rect 23566 14832 23572 14884
rect 23624 14872 23630 14884
rect 23753 14875 23811 14881
rect 23753 14872 23765 14875
rect 23624 14844 23765 14872
rect 23624 14832 23630 14844
rect 23753 14841 23765 14844
rect 23799 14841 23811 14875
rect 23753 14835 23811 14841
rect 21453 14807 21511 14813
rect 21453 14804 21465 14807
rect 21100 14776 21465 14804
rect 20625 14767 20683 14773
rect 21453 14773 21465 14776
rect 21499 14773 21511 14807
rect 21453 14767 21511 14773
rect 22002 14764 22008 14816
rect 22060 14804 22066 14816
rect 23382 14804 23388 14816
rect 22060 14776 23388 14804
rect 22060 14764 22066 14776
rect 23382 14764 23388 14776
rect 23440 14764 23446 14816
rect 1104 14714 28152 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 28152 14714
rect 1104 14640 28152 14662
rect 3326 14560 3332 14612
rect 3384 14560 3390 14612
rect 3786 14560 3792 14612
rect 3844 14600 3850 14612
rect 3844 14572 4108 14600
rect 3844 14560 3850 14572
rect 2593 14535 2651 14541
rect 2593 14501 2605 14535
rect 2639 14532 2651 14535
rect 2774 14532 2780 14544
rect 2639 14504 2780 14532
rect 2639 14501 2651 14504
rect 2593 14495 2651 14501
rect 2774 14492 2780 14504
rect 2832 14532 2838 14544
rect 2832 14504 3188 14532
rect 2832 14492 2838 14504
rect 2317 14467 2375 14473
rect 2317 14433 2329 14467
rect 2363 14464 2375 14467
rect 2682 14464 2688 14476
rect 2363 14436 2688 14464
rect 2363 14433 2375 14436
rect 2317 14427 2375 14433
rect 2682 14424 2688 14436
rect 2740 14424 2746 14476
rect 2866 14424 2872 14476
rect 2924 14424 2930 14476
rect 3160 14473 3188 14504
rect 3970 14492 3976 14544
rect 4028 14492 4034 14544
rect 4080 14541 4108 14572
rect 12066 14560 12072 14612
rect 12124 14600 12130 14612
rect 14918 14600 14924 14612
rect 12124 14572 14924 14600
rect 12124 14560 12130 14572
rect 14918 14560 14924 14572
rect 14976 14560 14982 14612
rect 15105 14603 15163 14609
rect 15105 14569 15117 14603
rect 15151 14600 15163 14603
rect 15286 14600 15292 14612
rect 15151 14572 15292 14600
rect 15151 14569 15163 14572
rect 15105 14563 15163 14569
rect 15286 14560 15292 14572
rect 15344 14560 15350 14612
rect 17034 14560 17040 14612
rect 17092 14600 17098 14612
rect 17589 14603 17647 14609
rect 17589 14600 17601 14603
rect 17092 14572 17601 14600
rect 17092 14560 17098 14572
rect 17589 14569 17601 14572
rect 17635 14569 17647 14603
rect 17589 14563 17647 14569
rect 18417 14603 18475 14609
rect 18417 14569 18429 14603
rect 18463 14569 18475 14603
rect 18417 14563 18475 14569
rect 4065 14535 4123 14541
rect 4065 14501 4077 14535
rect 4111 14501 4123 14535
rect 4065 14495 4123 14501
rect 4706 14492 4712 14544
rect 4764 14532 4770 14544
rect 5537 14535 5595 14541
rect 5537 14532 5549 14535
rect 4764 14504 5549 14532
rect 4764 14492 4770 14504
rect 5537 14501 5549 14504
rect 5583 14501 5595 14535
rect 5537 14495 5595 14501
rect 6365 14535 6423 14541
rect 6365 14501 6377 14535
rect 6411 14532 6423 14535
rect 7282 14532 7288 14544
rect 6411 14504 7288 14532
rect 6411 14501 6423 14504
rect 6365 14495 6423 14501
rect 7282 14492 7288 14504
rect 7340 14492 7346 14544
rect 16850 14492 16856 14544
rect 16908 14532 16914 14544
rect 17359 14535 17417 14541
rect 17359 14532 17371 14535
rect 16908 14504 17371 14532
rect 16908 14492 16914 14504
rect 17359 14501 17371 14504
rect 17405 14501 17417 14535
rect 18432 14532 18460 14563
rect 18598 14560 18604 14612
rect 18656 14560 18662 14612
rect 21358 14560 21364 14612
rect 21416 14600 21422 14612
rect 22097 14603 22155 14609
rect 22097 14600 22109 14603
rect 21416 14572 22109 14600
rect 21416 14560 21422 14572
rect 22097 14569 22109 14572
rect 22143 14600 22155 14603
rect 22554 14600 22560 14612
rect 22143 14572 22560 14600
rect 22143 14569 22155 14572
rect 22097 14563 22155 14569
rect 22554 14560 22560 14572
rect 22612 14560 22618 14612
rect 23106 14560 23112 14612
rect 23164 14600 23170 14612
rect 23750 14600 23756 14612
rect 23164 14572 23756 14600
rect 23164 14560 23170 14572
rect 23750 14560 23756 14572
rect 23808 14560 23814 14612
rect 19242 14532 19248 14544
rect 18432 14504 19248 14532
rect 17359 14495 17417 14501
rect 19242 14492 19248 14504
rect 19300 14492 19306 14544
rect 19426 14492 19432 14544
rect 19484 14492 19490 14544
rect 20622 14492 20628 14544
rect 20680 14492 20686 14544
rect 23290 14532 23296 14544
rect 22020 14504 23296 14532
rect 3145 14467 3203 14473
rect 3145 14433 3157 14467
rect 3191 14433 3203 14467
rect 3988 14464 4016 14492
rect 4341 14467 4399 14473
rect 3145 14427 3203 14433
rect 3620 14436 4200 14464
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 2406 14396 2412 14408
rect 2271 14368 2412 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 2406 14356 2412 14368
rect 2464 14356 2470 14408
rect 2961 14399 3019 14405
rect 2961 14365 2973 14399
rect 3007 14365 3019 14399
rect 2961 14359 3019 14365
rect 3053 14399 3111 14405
rect 3053 14365 3065 14399
rect 3099 14396 3111 14399
rect 3326 14396 3332 14408
rect 3099 14368 3332 14396
rect 3099 14365 3111 14368
rect 3053 14359 3111 14365
rect 2976 14328 3004 14359
rect 3326 14356 3332 14368
rect 3384 14356 3390 14408
rect 3620 14340 3648 14436
rect 3878 14356 3884 14408
rect 3936 14356 3942 14408
rect 4172 14405 4200 14436
rect 4341 14433 4353 14467
rect 4387 14464 4399 14467
rect 5258 14464 5264 14476
rect 4387 14436 5264 14464
rect 4387 14433 4399 14436
rect 4341 14427 4399 14433
rect 5258 14424 5264 14436
rect 5316 14424 5322 14476
rect 5721 14467 5779 14473
rect 5721 14433 5733 14467
rect 5767 14464 5779 14467
rect 5767 14436 6132 14464
rect 5767 14433 5779 14436
rect 5721 14427 5779 14433
rect 6104 14405 6132 14436
rect 6822 14424 6828 14476
rect 6880 14464 6886 14476
rect 6917 14467 6975 14473
rect 6917 14464 6929 14467
rect 6880 14436 6929 14464
rect 6880 14424 6886 14436
rect 6917 14433 6929 14436
rect 6963 14433 6975 14467
rect 6917 14427 6975 14433
rect 11057 14467 11115 14473
rect 11057 14433 11069 14467
rect 11103 14464 11115 14467
rect 13998 14464 14004 14476
rect 11103 14436 14004 14464
rect 11103 14433 11115 14436
rect 11057 14427 11115 14433
rect 13998 14424 14004 14436
rect 14056 14424 14062 14476
rect 14642 14424 14648 14476
rect 14700 14464 14706 14476
rect 14875 14467 14933 14473
rect 14875 14464 14887 14467
rect 14700 14436 14887 14464
rect 14700 14424 14706 14436
rect 14875 14433 14887 14436
rect 14921 14433 14933 14467
rect 14875 14427 14933 14433
rect 15013 14467 15071 14473
rect 15013 14433 15025 14467
rect 15059 14464 15071 14467
rect 15378 14464 15384 14476
rect 15059 14436 15384 14464
rect 15059 14433 15071 14436
rect 15013 14427 15071 14433
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 16945 14467 17003 14473
rect 16945 14433 16957 14467
rect 16991 14464 17003 14467
rect 17034 14464 17040 14476
rect 16991 14436 17040 14464
rect 16991 14433 17003 14436
rect 16945 14427 17003 14433
rect 17034 14424 17040 14436
rect 17092 14424 17098 14476
rect 17129 14467 17187 14473
rect 17129 14433 17141 14467
rect 17175 14464 17187 14467
rect 17175 14436 17264 14464
rect 17175 14433 17187 14436
rect 17129 14427 17187 14433
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 4157 14399 4215 14405
rect 4157 14365 4169 14399
rect 4203 14365 4215 14399
rect 4157 14359 4215 14365
rect 6089 14399 6147 14405
rect 6089 14365 6101 14399
rect 6135 14365 6147 14399
rect 6089 14359 6147 14365
rect 3142 14328 3148 14340
rect 2976 14300 3148 14328
rect 3142 14288 3148 14300
rect 3200 14328 3206 14340
rect 3602 14328 3608 14340
rect 3200 14300 3608 14328
rect 3200 14288 3206 14300
rect 3602 14288 3608 14300
rect 3660 14288 3666 14340
rect 3988 14328 4016 14359
rect 6730 14356 6736 14408
rect 6788 14356 6794 14408
rect 13173 14399 13231 14405
rect 13173 14365 13185 14399
rect 13219 14396 13231 14399
rect 13262 14396 13268 14408
rect 13219 14368 13268 14396
rect 13219 14365 13231 14368
rect 13173 14359 13231 14365
rect 13262 14356 13268 14368
rect 13320 14356 13326 14408
rect 13446 14356 13452 14408
rect 13504 14356 13510 14408
rect 14737 14399 14795 14405
rect 14737 14365 14749 14399
rect 14783 14365 14795 14399
rect 14737 14359 14795 14365
rect 3988 14300 4200 14328
rect 4172 14272 4200 14300
rect 11330 14288 11336 14340
rect 11388 14288 11394 14340
rect 14550 14328 14556 14340
rect 12558 14300 14556 14328
rect 14550 14288 14556 14300
rect 14608 14288 14614 14340
rect 14752 14328 14780 14359
rect 15194 14356 15200 14408
rect 15252 14356 15258 14408
rect 16850 14356 16856 14408
rect 16908 14356 16914 14408
rect 17052 14328 17080 14424
rect 17236 14408 17264 14436
rect 17954 14424 17960 14476
rect 18012 14464 18018 14476
rect 18233 14467 18291 14473
rect 18233 14464 18245 14467
rect 18012 14436 18245 14464
rect 18012 14424 18018 14436
rect 18233 14433 18245 14436
rect 18279 14433 18291 14467
rect 19613 14467 19671 14473
rect 19613 14464 19625 14467
rect 18233 14427 18291 14433
rect 18432 14436 19625 14464
rect 17218 14356 17224 14408
rect 17276 14356 17282 14408
rect 17497 14399 17555 14405
rect 17497 14365 17509 14399
rect 17543 14365 17555 14399
rect 17497 14359 17555 14365
rect 17512 14328 17540 14359
rect 17678 14356 17684 14408
rect 17736 14356 17742 14408
rect 18432 14405 18460 14436
rect 19613 14433 19625 14436
rect 19659 14464 19671 14467
rect 20070 14464 20076 14476
rect 19659 14436 20076 14464
rect 19659 14433 19671 14436
rect 19613 14427 19671 14433
rect 20070 14424 20076 14436
rect 20128 14424 20134 14476
rect 20898 14424 20904 14476
rect 20956 14464 20962 14476
rect 21174 14464 21180 14476
rect 20956 14436 21180 14464
rect 20956 14424 20962 14436
rect 21174 14424 21180 14436
rect 21232 14424 21238 14476
rect 18417 14399 18475 14405
rect 18417 14365 18429 14399
rect 18463 14365 18475 14399
rect 18417 14359 18475 14365
rect 19426 14356 19432 14408
rect 19484 14356 19490 14408
rect 19794 14356 19800 14408
rect 19852 14356 19858 14408
rect 20990 14356 20996 14408
rect 21048 14396 21054 14408
rect 22020 14396 22048 14504
rect 23290 14492 23296 14504
rect 23348 14532 23354 14544
rect 23385 14535 23443 14541
rect 23385 14532 23397 14535
rect 23348 14504 23397 14532
rect 23348 14492 23354 14504
rect 23385 14501 23397 14504
rect 23431 14501 23443 14535
rect 23934 14532 23940 14544
rect 23385 14495 23443 14501
rect 23584 14504 23940 14532
rect 22094 14424 22100 14476
rect 22152 14464 22158 14476
rect 22152 14436 22876 14464
rect 22152 14424 22158 14436
rect 22465 14399 22523 14405
rect 22465 14396 22477 14399
rect 21048 14368 22477 14396
rect 21048 14356 21054 14368
rect 22465 14365 22477 14368
rect 22511 14365 22523 14399
rect 22465 14359 22523 14365
rect 22557 14399 22615 14405
rect 22557 14365 22569 14399
rect 22603 14396 22615 14399
rect 22646 14396 22652 14408
rect 22603 14368 22652 14396
rect 22603 14365 22615 14368
rect 22557 14359 22615 14365
rect 22646 14356 22652 14368
rect 22704 14356 22710 14408
rect 22848 14405 22876 14436
rect 22741 14399 22799 14405
rect 22741 14365 22753 14399
rect 22787 14365 22799 14399
rect 22741 14359 22799 14365
rect 22833 14399 22891 14405
rect 22833 14365 22845 14399
rect 22879 14365 22891 14399
rect 22833 14359 22891 14365
rect 23477 14399 23535 14405
rect 23477 14365 23489 14399
rect 23523 14396 23535 14399
rect 23584 14396 23612 14504
rect 23934 14492 23940 14504
rect 23992 14532 23998 14544
rect 24762 14532 24768 14544
rect 23992 14504 24768 14532
rect 23992 14492 23998 14504
rect 24762 14492 24768 14504
rect 24820 14492 24826 14544
rect 23658 14424 23664 14476
rect 23716 14464 23722 14476
rect 23845 14467 23903 14473
rect 23845 14464 23857 14467
rect 23716 14436 23857 14464
rect 23716 14424 23722 14436
rect 23845 14433 23857 14436
rect 23891 14433 23903 14467
rect 23845 14427 23903 14433
rect 23523 14368 23612 14396
rect 23523 14365 23535 14368
rect 23477 14359 23535 14365
rect 14752 14300 14964 14328
rect 17052 14300 17540 14328
rect 14936 14272 14964 14300
rect 18138 14288 18144 14340
rect 18196 14288 18202 14340
rect 19334 14288 19340 14340
rect 19392 14328 19398 14340
rect 21818 14328 21824 14340
rect 19392 14300 21824 14328
rect 19392 14288 19398 14300
rect 21818 14288 21824 14300
rect 21876 14328 21882 14340
rect 22002 14328 22008 14340
rect 21876 14300 22008 14328
rect 21876 14288 21882 14300
rect 22002 14288 22008 14300
rect 22060 14288 22066 14340
rect 22756 14328 22784 14359
rect 23750 14356 23756 14408
rect 23808 14356 23814 14408
rect 23934 14356 23940 14408
rect 23992 14356 23998 14408
rect 24029 14399 24087 14405
rect 24029 14365 24041 14399
rect 24075 14396 24087 14399
rect 24210 14396 24216 14408
rect 24075 14368 24216 14396
rect 24075 14365 24087 14368
rect 24029 14359 24087 14365
rect 24210 14356 24216 14368
rect 24268 14356 24274 14408
rect 22572 14300 22784 14328
rect 4154 14220 4160 14272
rect 4212 14220 4218 14272
rect 12802 14220 12808 14272
rect 12860 14220 12866 14272
rect 12986 14220 12992 14272
rect 13044 14220 13050 14272
rect 13354 14220 13360 14272
rect 13412 14220 13418 14272
rect 14918 14220 14924 14272
rect 14976 14220 14982 14272
rect 17126 14220 17132 14272
rect 17184 14220 17190 14272
rect 19058 14220 19064 14272
rect 19116 14260 19122 14272
rect 22572 14260 22600 14300
rect 23382 14288 23388 14340
rect 23440 14328 23446 14340
rect 23440 14300 23704 14328
rect 23440 14288 23446 14300
rect 19116 14232 22600 14260
rect 19116 14220 19122 14232
rect 22922 14220 22928 14272
rect 22980 14260 22986 14272
rect 23017 14263 23075 14269
rect 23017 14260 23029 14263
rect 22980 14232 23029 14260
rect 22980 14220 22986 14232
rect 23017 14229 23029 14232
rect 23063 14229 23075 14263
rect 23017 14223 23075 14229
rect 23566 14220 23572 14272
rect 23624 14220 23630 14272
rect 23676 14260 23704 14300
rect 24486 14288 24492 14340
rect 24544 14288 24550 14340
rect 24581 14263 24639 14269
rect 24581 14260 24593 14263
rect 23676 14232 24593 14260
rect 24581 14229 24593 14232
rect 24627 14229 24639 14263
rect 24581 14223 24639 14229
rect 1104 14170 28152 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 28152 14170
rect 1104 14096 28152 14118
rect 3326 14056 3332 14068
rect 2148 14028 3332 14056
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 1946 13812 1952 13864
rect 2004 13852 2010 13864
rect 2148 13861 2176 14028
rect 3326 14016 3332 14028
rect 3384 14016 3390 14068
rect 3786 14016 3792 14068
rect 3844 14056 3850 14068
rect 4062 14056 4068 14068
rect 3844 14028 4068 14056
rect 3844 14016 3850 14028
rect 4062 14016 4068 14028
rect 4120 14056 4126 14068
rect 4120 14028 10732 14056
rect 4120 14016 4126 14028
rect 3237 13991 3295 13997
rect 3237 13988 3249 13991
rect 2700 13960 3249 13988
rect 2700 13929 2728 13960
rect 3237 13957 3249 13960
rect 3283 13957 3295 13991
rect 3237 13951 3295 13957
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13889 2743 13923
rect 2685 13883 2743 13889
rect 3142 13880 3148 13932
rect 3200 13880 3206 13932
rect 3344 13929 3372 14016
rect 3602 13948 3608 14000
rect 3660 13988 3666 14000
rect 3881 13991 3939 13997
rect 3660 13960 3832 13988
rect 3660 13948 3666 13960
rect 3804 13929 3832 13960
rect 3881 13957 3893 13991
rect 3927 13988 3939 13991
rect 7926 13988 7932 14000
rect 3927 13960 4384 13988
rect 3927 13957 3939 13960
rect 3881 13951 3939 13957
rect 3329 13923 3387 13929
rect 3329 13889 3341 13923
rect 3375 13889 3387 13923
rect 3329 13883 3387 13889
rect 3795 13923 3853 13929
rect 3795 13889 3807 13923
rect 3841 13889 3853 13923
rect 3795 13883 3853 13889
rect 3973 13923 4031 13929
rect 3973 13889 3985 13923
rect 4019 13920 4031 13923
rect 4062 13920 4068 13932
rect 4019 13892 4068 13920
rect 4019 13889 4031 13892
rect 3973 13883 4031 13889
rect 2133 13855 2191 13861
rect 2133 13852 2145 13855
rect 2004 13824 2145 13852
rect 2004 13812 2010 13824
rect 2133 13821 2145 13824
rect 2179 13821 2191 13855
rect 2133 13815 2191 13821
rect 2774 13812 2780 13864
rect 2832 13812 2838 13864
rect 3344 13852 3372 13883
rect 4062 13880 4068 13892
rect 4120 13880 4126 13932
rect 4154 13880 4160 13932
rect 4212 13880 4218 13932
rect 4356 13929 4384 13960
rect 6472 13960 7932 13988
rect 4341 13923 4399 13929
rect 4341 13889 4353 13923
rect 4387 13889 4399 13923
rect 6472 13920 6500 13960
rect 7926 13948 7932 13960
rect 7984 13948 7990 14000
rect 4341 13883 4399 13889
rect 4448 13892 6500 13920
rect 6549 13923 6607 13929
rect 4448 13852 4476 13892
rect 6549 13889 6561 13923
rect 6595 13920 6607 13923
rect 6730 13920 6736 13932
rect 6595 13892 6736 13920
rect 6595 13889 6607 13892
rect 6549 13883 6607 13889
rect 6730 13880 6736 13892
rect 6788 13880 6794 13932
rect 10502 13880 10508 13932
rect 10560 13920 10566 13932
rect 10597 13923 10655 13929
rect 10597 13920 10609 13923
rect 10560 13892 10609 13920
rect 10560 13880 10566 13892
rect 10597 13889 10609 13892
rect 10643 13889 10655 13923
rect 10597 13883 10655 13889
rect 3344 13824 4476 13852
rect 5169 13855 5227 13861
rect 5169 13821 5181 13855
rect 5215 13852 5227 13855
rect 5534 13852 5540 13864
rect 5215 13824 5540 13852
rect 5215 13821 5227 13824
rect 5169 13815 5227 13821
rect 5534 13812 5540 13824
rect 5592 13812 5598 13864
rect 6641 13855 6699 13861
rect 6641 13821 6653 13855
rect 6687 13852 6699 13855
rect 6822 13852 6828 13864
rect 6687 13824 6828 13852
rect 6687 13821 6699 13824
rect 6641 13815 6699 13821
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 8294 13812 8300 13864
rect 8352 13852 8358 13864
rect 10704 13861 10732 14028
rect 11330 14016 11336 14068
rect 11388 14056 11394 14068
rect 11609 14059 11667 14065
rect 11609 14056 11621 14059
rect 11388 14028 11621 14056
rect 11388 14016 11394 14028
rect 11609 14025 11621 14028
rect 11655 14025 11667 14059
rect 11609 14019 11667 14025
rect 11885 14059 11943 14065
rect 11885 14025 11897 14059
rect 11931 14056 11943 14059
rect 11974 14056 11980 14068
rect 11931 14028 11980 14056
rect 11931 14025 11943 14028
rect 11885 14019 11943 14025
rect 11701 13923 11759 13929
rect 11701 13889 11713 13923
rect 11747 13920 11759 13923
rect 11900 13920 11928 14019
rect 11974 14016 11980 14028
rect 12032 14016 12038 14068
rect 12250 14056 12256 14068
rect 12176 14028 12256 14056
rect 12176 13929 12204 14028
rect 12250 14016 12256 14028
rect 12308 14016 12314 14068
rect 15654 14016 15660 14068
rect 15712 14056 15718 14068
rect 15841 14059 15899 14065
rect 15841 14056 15853 14059
rect 15712 14028 15853 14056
rect 15712 14016 15718 14028
rect 15841 14025 15853 14028
rect 15887 14025 15899 14059
rect 15841 14019 15899 14025
rect 20806 14016 20812 14068
rect 20864 14056 20870 14068
rect 20864 14028 22048 14056
rect 20864 14016 20870 14028
rect 12986 13988 12992 14000
rect 12360 13960 12992 13988
rect 12360 13929 12388 13960
rect 12986 13948 12992 13960
rect 13044 13948 13050 14000
rect 14384 13960 14780 13988
rect 11747 13892 11928 13920
rect 12161 13923 12219 13929
rect 11747 13889 11759 13892
rect 11701 13883 11759 13889
rect 12161 13889 12173 13923
rect 12207 13889 12219 13923
rect 12161 13883 12219 13889
rect 12345 13923 12403 13929
rect 12345 13889 12357 13923
rect 12391 13889 12403 13923
rect 12345 13883 12403 13889
rect 12529 13923 12587 13929
rect 12529 13889 12541 13923
rect 12575 13920 12587 13923
rect 12802 13920 12808 13932
rect 12575 13892 12808 13920
rect 12575 13889 12587 13892
rect 12529 13883 12587 13889
rect 8481 13855 8539 13861
rect 8481 13852 8493 13855
rect 8352 13824 8493 13852
rect 8352 13812 8358 13824
rect 8481 13821 8493 13824
rect 8527 13821 8539 13855
rect 8481 13815 8539 13821
rect 10689 13855 10747 13861
rect 10689 13821 10701 13855
rect 10735 13852 10747 13855
rect 11054 13852 11060 13864
rect 10735 13824 11060 13852
rect 10735 13821 10747 13824
rect 10689 13815 10747 13821
rect 11054 13812 11060 13824
rect 11112 13852 11118 13864
rect 11974 13852 11980 13864
rect 11112 13824 11980 13852
rect 11112 13812 11118 13824
rect 11974 13812 11980 13824
rect 12032 13812 12038 13864
rect 12066 13812 12072 13864
rect 12124 13812 12130 13864
rect 12253 13855 12311 13861
rect 12253 13821 12265 13855
rect 12299 13852 12311 13855
rect 12434 13852 12440 13864
rect 12299 13824 12440 13852
rect 12299 13821 12311 13824
rect 12253 13815 12311 13821
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 3050 13744 3056 13796
rect 3108 13744 3114 13796
rect 8570 13744 8576 13796
rect 8628 13784 8634 13796
rect 8757 13787 8815 13793
rect 8757 13784 8769 13787
rect 8628 13756 8769 13784
rect 8628 13744 8634 13756
rect 8757 13753 8769 13756
rect 8803 13753 8815 13787
rect 8757 13747 8815 13753
rect 12342 13744 12348 13796
rect 12400 13784 12406 13796
rect 12544 13784 12572 13883
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 14384 13929 14412 13960
rect 14369 13923 14427 13929
rect 14369 13889 14381 13923
rect 14415 13889 14427 13923
rect 14369 13883 14427 13889
rect 14553 13923 14611 13929
rect 14553 13889 14565 13923
rect 14599 13920 14611 13923
rect 14599 13892 14688 13920
rect 14599 13889 14611 13892
rect 14553 13883 14611 13889
rect 14660 13864 14688 13892
rect 14642 13812 14648 13864
rect 14700 13812 14706 13864
rect 14752 13861 14780 13960
rect 14826 13948 14832 14000
rect 14884 13988 14890 14000
rect 15473 13991 15531 13997
rect 15473 13988 15485 13991
rect 14884 13960 15485 13988
rect 14884 13948 14890 13960
rect 15473 13957 15485 13960
rect 15519 13957 15531 13991
rect 15473 13951 15531 13957
rect 15565 13991 15623 13997
rect 15565 13957 15577 13991
rect 15611 13988 15623 13991
rect 18601 13991 18659 13997
rect 15611 13960 18092 13988
rect 15611 13957 15623 13960
rect 15565 13951 15623 13957
rect 14918 13880 14924 13932
rect 14976 13880 14982 13932
rect 15010 13880 15016 13932
rect 15068 13920 15074 13932
rect 18064 13929 18092 13960
rect 18601 13957 18613 13991
rect 18647 13988 18659 13991
rect 18647 13960 21588 13988
rect 18647 13957 18659 13960
rect 18601 13951 18659 13957
rect 15289 13923 15347 13929
rect 15289 13920 15301 13923
rect 15068 13892 15301 13920
rect 15068 13880 15074 13892
rect 15289 13889 15301 13892
rect 15335 13889 15347 13923
rect 15289 13883 15347 13889
rect 15657 13923 15715 13929
rect 15657 13889 15669 13923
rect 15703 13920 15715 13923
rect 18049 13923 18107 13929
rect 15703 13892 17816 13920
rect 15703 13889 15715 13892
rect 15657 13883 15715 13889
rect 14737 13855 14795 13861
rect 14737 13821 14749 13855
rect 14783 13852 14795 13855
rect 15378 13852 15384 13864
rect 14783 13824 15384 13852
rect 14783 13821 14795 13824
rect 14737 13815 14795 13821
rect 15378 13812 15384 13824
rect 15436 13852 15442 13864
rect 15930 13852 15936 13864
rect 15436 13824 15936 13852
rect 15436 13812 15442 13824
rect 15930 13812 15936 13824
rect 15988 13812 15994 13864
rect 17788 13852 17816 13892
rect 18049 13889 18061 13923
rect 18095 13920 18107 13923
rect 18230 13920 18236 13932
rect 18095 13892 18236 13920
rect 18095 13889 18107 13892
rect 18049 13883 18107 13889
rect 18230 13880 18236 13892
rect 18288 13880 18294 13932
rect 18322 13880 18328 13932
rect 18380 13880 18386 13932
rect 18417 13923 18475 13929
rect 18417 13889 18429 13923
rect 18463 13920 18475 13923
rect 18506 13920 18512 13932
rect 18463 13892 18512 13920
rect 18463 13889 18475 13892
rect 18417 13883 18475 13889
rect 18506 13880 18512 13892
rect 18564 13880 18570 13932
rect 19610 13920 19616 13932
rect 18616 13892 19616 13920
rect 18141 13855 18199 13861
rect 18141 13852 18153 13855
rect 17788 13824 18153 13852
rect 18141 13821 18153 13824
rect 18187 13852 18199 13855
rect 18616 13852 18644 13892
rect 19610 13880 19616 13892
rect 19668 13880 19674 13932
rect 18187 13824 18644 13852
rect 18187 13821 18199 13824
rect 18141 13815 18199 13821
rect 12400 13756 12572 13784
rect 12400 13744 12406 13756
rect 15102 13744 15108 13796
rect 15160 13744 15166 13796
rect 16114 13744 16120 13796
rect 16172 13784 16178 13796
rect 18874 13784 18880 13796
rect 16172 13756 18880 13784
rect 16172 13744 16178 13756
rect 18874 13744 18880 13756
rect 18932 13784 18938 13796
rect 20898 13784 20904 13796
rect 18932 13756 20904 13784
rect 18932 13744 18938 13756
rect 20898 13744 20904 13756
rect 20956 13784 20962 13796
rect 21450 13784 21456 13796
rect 20956 13756 21456 13784
rect 20956 13744 20962 13756
rect 21450 13744 21456 13756
rect 21508 13744 21514 13796
rect 21560 13784 21588 13960
rect 22020 13929 22048 14028
rect 22370 14016 22376 14068
rect 22428 14016 22434 14068
rect 22557 14059 22615 14065
rect 22557 14025 22569 14059
rect 22603 14056 22615 14059
rect 23474 14056 23480 14068
rect 22603 14028 23480 14056
rect 22603 14025 22615 14028
rect 22557 14019 22615 14025
rect 23474 14016 23480 14028
rect 23532 14056 23538 14068
rect 23532 14028 23888 14056
rect 23532 14016 23538 14028
rect 23566 13988 23572 14000
rect 23032 13960 23572 13988
rect 22005 13923 22063 13929
rect 22005 13889 22017 13923
rect 22051 13889 22063 13923
rect 22005 13883 22063 13889
rect 22094 13880 22100 13932
rect 22152 13880 22158 13932
rect 22922 13880 22928 13932
rect 22980 13880 22986 13932
rect 21913 13855 21971 13861
rect 21913 13821 21925 13855
rect 21959 13852 21971 13855
rect 22189 13855 22247 13861
rect 21959 13824 22140 13852
rect 21959 13821 21971 13824
rect 21913 13815 21971 13821
rect 22002 13784 22008 13796
rect 21560 13756 22008 13784
rect 22002 13744 22008 13756
rect 22060 13744 22066 13796
rect 22112 13784 22140 13824
rect 22189 13821 22201 13855
rect 22235 13852 22247 13855
rect 22278 13852 22284 13864
rect 22235 13824 22284 13852
rect 22235 13821 22247 13824
rect 22189 13815 22247 13821
rect 22278 13812 22284 13824
rect 22336 13812 22342 13864
rect 22465 13855 22523 13861
rect 22465 13821 22477 13855
rect 22511 13852 22523 13855
rect 22554 13852 22560 13864
rect 22511 13824 22560 13852
rect 22511 13821 22523 13824
rect 22465 13815 22523 13821
rect 22554 13812 22560 13824
rect 22612 13812 22618 13864
rect 23032 13861 23060 13960
rect 23566 13948 23572 13960
rect 23624 13948 23630 14000
rect 23860 13997 23888 14028
rect 24762 14016 24768 14068
rect 24820 14056 24826 14068
rect 25317 14059 25375 14065
rect 25317 14056 25329 14059
rect 24820 14028 25329 14056
rect 24820 14016 24826 14028
rect 25317 14025 25329 14028
rect 25363 14025 25375 14059
rect 25317 14019 25375 14025
rect 25774 14016 25780 14068
rect 25832 14056 25838 14068
rect 27617 14059 27675 14065
rect 27617 14056 27629 14059
rect 25832 14028 27629 14056
rect 25832 14016 25838 14028
rect 27617 14025 27629 14028
rect 27663 14025 27675 14059
rect 27617 14019 27675 14025
rect 23845 13991 23903 13997
rect 23845 13957 23857 13991
rect 23891 13957 23903 13991
rect 23845 13951 23903 13957
rect 25130 13948 25136 14000
rect 25188 13988 25194 14000
rect 25501 13991 25559 13997
rect 25501 13988 25513 13991
rect 25188 13960 25513 13988
rect 25188 13948 25194 13960
rect 25501 13957 25513 13960
rect 25547 13957 25559 13991
rect 25501 13951 25559 13957
rect 23290 13880 23296 13932
rect 23348 13880 23354 13932
rect 23382 13880 23388 13932
rect 23440 13880 23446 13932
rect 24946 13880 24952 13932
rect 25004 13880 25010 13932
rect 27522 13880 27528 13932
rect 27580 13920 27586 13932
rect 27801 13923 27859 13929
rect 27801 13920 27813 13923
rect 27580 13892 27813 13920
rect 27580 13880 27586 13892
rect 27801 13889 27813 13892
rect 27847 13889 27859 13923
rect 27801 13883 27859 13889
rect 23017 13855 23075 13861
rect 23017 13821 23029 13855
rect 23063 13821 23075 13855
rect 23017 13815 23075 13821
rect 23106 13812 23112 13864
rect 23164 13852 23170 13864
rect 23164 13824 23428 13852
rect 23164 13812 23170 13824
rect 23400 13796 23428 13824
rect 23566 13812 23572 13864
rect 23624 13812 23630 13864
rect 24210 13812 24216 13864
rect 24268 13852 24274 13864
rect 25777 13855 25835 13861
rect 25777 13852 25789 13855
rect 24268 13824 25789 13852
rect 24268 13812 24274 13824
rect 25777 13821 25789 13824
rect 25823 13821 25835 13855
rect 25777 13815 25835 13821
rect 22370 13784 22376 13796
rect 22112 13756 22376 13784
rect 22370 13744 22376 13756
rect 22428 13744 22434 13796
rect 23382 13744 23388 13796
rect 23440 13744 23446 13796
rect 6822 13676 6828 13728
rect 6880 13676 6886 13728
rect 8938 13676 8944 13728
rect 8996 13676 9002 13728
rect 12158 13676 12164 13728
rect 12216 13716 12222 13728
rect 12621 13719 12679 13725
rect 12621 13716 12633 13719
rect 12216 13688 12633 13716
rect 12216 13676 12222 13688
rect 12621 13685 12633 13688
rect 12667 13716 12679 13719
rect 13354 13716 13360 13728
rect 12667 13688 13360 13716
rect 12667 13685 12679 13688
rect 12621 13679 12679 13685
rect 13354 13676 13360 13688
rect 13412 13676 13418 13728
rect 14366 13676 14372 13728
rect 14424 13676 14430 13728
rect 15286 13676 15292 13728
rect 15344 13716 15350 13728
rect 17770 13716 17776 13728
rect 15344 13688 17776 13716
rect 15344 13676 15350 13688
rect 17770 13676 17776 13688
rect 17828 13676 17834 13728
rect 1104 13626 28152 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 28152 13626
rect 1104 13552 28152 13574
rect 2406 13472 2412 13524
rect 2464 13472 2470 13524
rect 7377 13515 7435 13521
rect 7377 13481 7389 13515
rect 7423 13512 7435 13515
rect 8570 13512 8576 13524
rect 7423 13484 8576 13512
rect 7423 13481 7435 13484
rect 7377 13475 7435 13481
rect 8570 13472 8576 13484
rect 8628 13472 8634 13524
rect 8662 13472 8668 13524
rect 8720 13472 8726 13524
rect 12066 13472 12072 13524
rect 12124 13512 12130 13524
rect 12161 13515 12219 13521
rect 12161 13512 12173 13515
rect 12124 13484 12173 13512
rect 12124 13472 12130 13484
rect 12161 13481 12173 13484
rect 12207 13481 12219 13515
rect 12161 13475 12219 13481
rect 12434 13472 12440 13524
rect 12492 13472 12498 13524
rect 22738 13512 22744 13524
rect 14200 13484 22744 13512
rect 7837 13447 7895 13453
rect 7837 13413 7849 13447
rect 7883 13413 7895 13447
rect 7837 13407 7895 13413
rect 1946 13336 1952 13388
rect 2004 13336 2010 13388
rect 2222 13336 2228 13388
rect 2280 13336 2286 13388
rect 7852 13376 7880 13407
rect 11882 13404 11888 13456
rect 11940 13444 11946 13456
rect 14200 13444 14228 13484
rect 22738 13472 22744 13484
rect 22796 13472 22802 13524
rect 22925 13515 22983 13521
rect 22925 13481 22937 13515
rect 22971 13512 22983 13515
rect 23201 13515 23259 13521
rect 23201 13512 23213 13515
rect 22971 13484 23213 13512
rect 22971 13481 22983 13484
rect 22925 13475 22983 13481
rect 23201 13481 23213 13484
rect 23247 13481 23259 13515
rect 23201 13475 23259 13481
rect 11940 13416 14228 13444
rect 11940 13404 11946 13416
rect 15930 13404 15936 13456
rect 15988 13404 15994 13456
rect 17402 13404 17408 13456
rect 17460 13404 17466 13456
rect 17862 13404 17868 13456
rect 17920 13444 17926 13456
rect 17920 13416 21404 13444
rect 17920 13404 17926 13416
rect 8294 13376 8300 13388
rect 7116 13348 7604 13376
rect 7852 13348 8300 13376
rect 1854 13268 1860 13320
rect 1912 13268 1918 13320
rect 2240 13308 2268 13336
rect 7116 13320 7144 13348
rect 2317 13311 2375 13317
rect 2317 13308 2329 13311
rect 2240 13280 2329 13308
rect 2317 13277 2329 13280
rect 2363 13277 2375 13311
rect 2317 13271 2375 13277
rect 2501 13311 2559 13317
rect 2501 13277 2513 13311
rect 2547 13308 2559 13311
rect 2958 13308 2964 13320
rect 2547 13280 2964 13308
rect 2547 13277 2559 13280
rect 2501 13271 2559 13277
rect 2958 13268 2964 13280
rect 3016 13268 3022 13320
rect 6822 13268 6828 13320
rect 6880 13268 6886 13320
rect 7098 13268 7104 13320
rect 7156 13268 7162 13320
rect 7466 13268 7472 13320
rect 7524 13268 7530 13320
rect 7576 13317 7604 13348
rect 7561 13311 7619 13317
rect 7561 13277 7573 13311
rect 7607 13277 7619 13311
rect 7561 13271 7619 13277
rect 8110 13268 8116 13320
rect 8168 13268 8174 13320
rect 8220 13317 8248 13348
rect 8294 13336 8300 13348
rect 8352 13336 8358 13388
rect 12802 13376 12808 13388
rect 12360 13348 12808 13376
rect 8205 13311 8263 13317
rect 8205 13277 8217 13311
rect 8251 13277 8263 13311
rect 8205 13271 8263 13277
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 8481 13311 8539 13317
rect 8481 13277 8493 13311
rect 8527 13277 8539 13311
rect 8481 13271 8539 13277
rect 6840 13172 6868 13268
rect 7484 13240 7512 13268
rect 7653 13243 7711 13249
rect 7653 13240 7665 13243
rect 7484 13212 7665 13240
rect 7653 13209 7665 13212
rect 7699 13209 7711 13243
rect 7653 13203 7711 13209
rect 7837 13243 7895 13249
rect 7837 13209 7849 13243
rect 7883 13209 7895 13243
rect 7837 13203 7895 13209
rect 7852 13172 7880 13203
rect 8294 13200 8300 13252
rect 8352 13240 8358 13252
rect 8404 13240 8432 13271
rect 8352 13212 8432 13240
rect 8352 13200 8358 13212
rect 6840 13144 7880 13172
rect 8018 13132 8024 13184
rect 8076 13172 8082 13184
rect 8496 13172 8524 13271
rect 8938 13268 8944 13320
rect 8996 13308 9002 13320
rect 9033 13311 9091 13317
rect 9033 13308 9045 13311
rect 8996 13280 9045 13308
rect 8996 13268 9002 13280
rect 9033 13277 9045 13280
rect 9079 13277 9091 13311
rect 9033 13271 9091 13277
rect 9214 13268 9220 13320
rect 9272 13268 9278 13320
rect 12250 13268 12256 13320
rect 12308 13268 12314 13320
rect 12360 13317 12388 13348
rect 12802 13336 12808 13348
rect 12860 13336 12866 13388
rect 13998 13336 14004 13388
rect 14056 13376 14062 13388
rect 14093 13379 14151 13385
rect 14093 13376 14105 13379
rect 14056 13348 14105 13376
rect 14056 13336 14062 13348
rect 14093 13345 14105 13348
rect 14139 13376 14151 13379
rect 16666 13376 16672 13388
rect 14139 13348 16672 13376
rect 14139 13345 14151 13348
rect 14093 13339 14151 13345
rect 16666 13336 16672 13348
rect 16724 13336 16730 13388
rect 17681 13379 17739 13385
rect 17681 13345 17693 13379
rect 17727 13376 17739 13379
rect 18046 13376 18052 13388
rect 17727 13348 18052 13376
rect 17727 13345 17739 13348
rect 17681 13339 17739 13345
rect 18046 13336 18052 13348
rect 18104 13336 18110 13388
rect 19334 13336 19340 13388
rect 19392 13376 19398 13388
rect 19978 13376 19984 13388
rect 19392 13348 19984 13376
rect 19392 13336 19398 13348
rect 19978 13336 19984 13348
rect 20036 13376 20042 13388
rect 20036 13348 20208 13376
rect 20036 13336 20042 13348
rect 12345 13311 12403 13317
rect 12345 13277 12357 13311
rect 12391 13277 12403 13311
rect 12345 13271 12403 13277
rect 12437 13311 12495 13317
rect 12437 13277 12449 13311
rect 12483 13277 12495 13311
rect 12437 13271 12495 13277
rect 12989 13311 13047 13317
rect 12989 13277 13001 13311
rect 13035 13308 13047 13311
rect 13906 13308 13912 13320
rect 13035 13280 13912 13308
rect 13035 13277 13047 13280
rect 12989 13271 13047 13277
rect 10045 13243 10103 13249
rect 10045 13209 10057 13243
rect 10091 13209 10103 13243
rect 12268 13240 12296 13268
rect 12452 13240 12480 13271
rect 13906 13268 13912 13280
rect 13964 13268 13970 13320
rect 16117 13311 16175 13317
rect 16117 13277 16129 13311
rect 16163 13308 16175 13311
rect 16206 13308 16212 13320
rect 16163 13280 16212 13308
rect 16163 13277 16175 13280
rect 16117 13271 16175 13277
rect 16206 13268 16212 13280
rect 16264 13268 16270 13320
rect 16393 13311 16451 13317
rect 16393 13277 16405 13311
rect 16439 13277 16451 13311
rect 16393 13271 16451 13277
rect 12268 13212 12480 13240
rect 10045 13203 10103 13209
rect 8076 13144 8524 13172
rect 10060 13172 10088 13203
rect 12618 13200 12624 13252
rect 12676 13200 12682 13252
rect 14366 13200 14372 13252
rect 14424 13200 14430 13252
rect 14826 13240 14832 13252
rect 14568 13212 14832 13240
rect 14568 13184 14596 13212
rect 14826 13200 14832 13212
rect 14884 13200 14890 13252
rect 16408 13240 16436 13271
rect 16942 13268 16948 13320
rect 17000 13308 17006 13320
rect 17494 13308 17500 13320
rect 17000 13280 17500 13308
rect 17000 13268 17006 13280
rect 17494 13268 17500 13280
rect 17552 13268 17558 13320
rect 17589 13311 17647 13317
rect 17589 13277 17601 13311
rect 17635 13277 17647 13311
rect 17589 13271 17647 13277
rect 16132 13212 16436 13240
rect 16132 13184 16160 13212
rect 17034 13200 17040 13252
rect 17092 13240 17098 13252
rect 17313 13243 17371 13249
rect 17313 13240 17325 13243
rect 17092 13212 17325 13240
rect 17092 13200 17098 13212
rect 17313 13209 17325 13212
rect 17359 13209 17371 13243
rect 17604 13240 17632 13271
rect 17862 13268 17868 13320
rect 17920 13268 17926 13320
rect 20180 13317 20208 13348
rect 20165 13311 20223 13317
rect 20165 13277 20177 13311
rect 20211 13277 20223 13311
rect 20165 13271 20223 13277
rect 20533 13311 20591 13317
rect 20533 13277 20545 13311
rect 20579 13308 20591 13311
rect 21266 13308 21272 13320
rect 20579 13280 21272 13308
rect 20579 13277 20591 13280
rect 20533 13271 20591 13277
rect 21266 13268 21272 13280
rect 21324 13268 21330 13320
rect 19334 13240 19340 13252
rect 17604 13212 19340 13240
rect 17313 13203 17371 13209
rect 19334 13200 19340 13212
rect 19392 13200 19398 13252
rect 12710 13172 12716 13184
rect 10060 13144 12716 13172
rect 8076 13132 8082 13144
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 12802 13132 12808 13184
rect 12860 13132 12866 13184
rect 14550 13132 14556 13184
rect 14608 13132 14614 13184
rect 15746 13132 15752 13184
rect 15804 13172 15810 13184
rect 15841 13175 15899 13181
rect 15841 13172 15853 13175
rect 15804 13144 15853 13172
rect 15804 13132 15810 13144
rect 15841 13141 15853 13144
rect 15887 13141 15899 13175
rect 15841 13135 15899 13141
rect 16114 13132 16120 13184
rect 16172 13132 16178 13184
rect 16298 13132 16304 13184
rect 16356 13132 16362 13184
rect 20070 13132 20076 13184
rect 20128 13132 20134 13184
rect 20254 13132 20260 13184
rect 20312 13172 20318 13184
rect 20441 13175 20499 13181
rect 20441 13172 20453 13175
rect 20312 13144 20453 13172
rect 20312 13132 20318 13144
rect 20441 13141 20453 13144
rect 20487 13141 20499 13175
rect 21376 13172 21404 13416
rect 22002 13404 22008 13456
rect 22060 13444 22066 13456
rect 22060 13416 23888 13444
rect 22060 13404 22066 13416
rect 21450 13336 21456 13388
rect 21508 13376 21514 13388
rect 21508 13348 23060 13376
rect 21508 13336 21514 13348
rect 21542 13268 21548 13320
rect 21600 13308 21606 13320
rect 21913 13311 21971 13317
rect 21913 13308 21925 13311
rect 21600 13280 21925 13308
rect 21600 13268 21606 13280
rect 21913 13277 21925 13280
rect 21959 13277 21971 13311
rect 21913 13271 21971 13277
rect 22094 13268 22100 13320
rect 22152 13268 22158 13320
rect 22278 13268 22284 13320
rect 22336 13308 22342 13320
rect 22465 13311 22523 13317
rect 22465 13308 22477 13311
rect 22336 13280 22477 13308
rect 22336 13268 22342 13280
rect 22465 13277 22477 13280
rect 22511 13277 22523 13311
rect 22465 13271 22523 13277
rect 22830 13268 22836 13320
rect 22888 13268 22894 13320
rect 22922 13268 22928 13320
rect 22980 13268 22986 13320
rect 23032 13308 23060 13348
rect 23474 13336 23480 13388
rect 23532 13336 23538 13388
rect 23860 13376 23888 13416
rect 23934 13404 23940 13456
rect 23992 13444 23998 13456
rect 24397 13447 24455 13453
rect 24397 13444 24409 13447
rect 23992 13416 24409 13444
rect 23992 13404 23998 13416
rect 24397 13413 24409 13416
rect 24443 13413 24455 13447
rect 24397 13407 24455 13413
rect 24026 13376 24032 13388
rect 23860 13348 24032 13376
rect 24026 13336 24032 13348
rect 24084 13376 24090 13388
rect 24673 13379 24731 13385
rect 24673 13376 24685 13379
rect 24084 13348 24685 13376
rect 24084 13336 24090 13348
rect 24673 13345 24685 13348
rect 24719 13345 24731 13379
rect 24673 13339 24731 13345
rect 23569 13311 23627 13317
rect 23569 13308 23581 13311
rect 23032 13280 23581 13308
rect 23569 13277 23581 13280
rect 23615 13277 23627 13311
rect 23569 13271 23627 13277
rect 24762 13268 24768 13320
rect 24820 13268 24826 13320
rect 22066 13212 22416 13240
rect 22066 13172 22094 13212
rect 21376 13144 22094 13172
rect 20441 13135 20499 13141
rect 22278 13132 22284 13184
rect 22336 13132 22342 13184
rect 22388 13172 22416 13212
rect 23109 13175 23167 13181
rect 23109 13172 23121 13175
rect 22388 13144 23121 13172
rect 23109 13141 23121 13144
rect 23155 13141 23167 13175
rect 23109 13135 23167 13141
rect 1104 13082 28152 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 28152 13082
rect 1104 13008 28152 13030
rect 6641 12971 6699 12977
rect 6641 12937 6653 12971
rect 6687 12968 6699 12971
rect 7098 12968 7104 12980
rect 6687 12940 7104 12968
rect 6687 12937 6699 12940
rect 6641 12931 6699 12937
rect 7098 12928 7104 12940
rect 7156 12928 7162 12980
rect 8113 12971 8171 12977
rect 8113 12937 8125 12971
rect 8159 12968 8171 12971
rect 8294 12968 8300 12980
rect 8159 12940 8300 12968
rect 8159 12937 8171 12940
rect 8113 12931 8171 12937
rect 8294 12928 8300 12940
rect 8352 12928 8358 12980
rect 8481 12971 8539 12977
rect 8481 12937 8493 12971
rect 8527 12968 8539 12971
rect 9214 12968 9220 12980
rect 8527 12940 9220 12968
rect 8527 12937 8539 12940
rect 8481 12931 8539 12937
rect 9214 12928 9220 12940
rect 9272 12928 9278 12980
rect 12250 12928 12256 12980
rect 12308 12928 12314 12980
rect 12437 12971 12495 12977
rect 12437 12937 12449 12971
rect 12483 12968 12495 12971
rect 12618 12968 12624 12980
rect 12483 12940 12624 12968
rect 12483 12937 12495 12940
rect 12437 12931 12495 12937
rect 12618 12928 12624 12940
rect 12676 12928 12682 12980
rect 14642 12928 14648 12980
rect 14700 12968 14706 12980
rect 14921 12971 14979 12977
rect 14921 12968 14933 12971
rect 14700 12940 14933 12968
rect 14700 12928 14706 12940
rect 14921 12937 14933 12940
rect 14967 12937 14979 12971
rect 14921 12931 14979 12937
rect 15028 12940 18184 12968
rect 8312 12900 8340 12928
rect 11885 12903 11943 12909
rect 8312 12872 8892 12900
rect 1949 12835 2007 12841
rect 1949 12801 1961 12835
rect 1995 12832 2007 12835
rect 2958 12832 2964 12844
rect 1995 12804 2964 12832
rect 1995 12801 2007 12804
rect 1949 12795 2007 12801
rect 2958 12792 2964 12804
rect 3016 12792 3022 12844
rect 5534 12792 5540 12844
rect 5592 12792 5598 12844
rect 6178 12792 6184 12844
rect 6236 12832 6242 12844
rect 6457 12835 6515 12841
rect 6457 12832 6469 12835
rect 6236 12804 6469 12832
rect 6236 12792 6242 12804
rect 6457 12801 6469 12804
rect 6503 12801 6515 12835
rect 6457 12795 6515 12801
rect 6638 12792 6644 12844
rect 6696 12792 6702 12844
rect 8018 12792 8024 12844
rect 8076 12792 8082 12844
rect 8202 12792 8208 12844
rect 8260 12832 8266 12844
rect 8864 12841 8892 12872
rect 11885 12869 11897 12903
rect 11931 12869 11943 12903
rect 11885 12863 11943 12869
rect 8297 12835 8355 12841
rect 8297 12832 8309 12835
rect 8260 12804 8309 12832
rect 8260 12792 8266 12804
rect 8297 12801 8309 12804
rect 8343 12801 8355 12835
rect 8297 12795 8355 12801
rect 8849 12835 8907 12841
rect 8849 12801 8861 12835
rect 8895 12801 8907 12835
rect 8849 12795 8907 12801
rect 11422 12792 11428 12844
rect 11480 12832 11486 12844
rect 11900 12832 11928 12863
rect 12066 12860 12072 12912
rect 12124 12909 12130 12912
rect 12124 12903 12143 12909
rect 12131 12869 12143 12903
rect 12124 12863 12143 12869
rect 12124 12860 12130 12863
rect 12710 12860 12716 12912
rect 12768 12900 12774 12912
rect 15028 12900 15056 12940
rect 15841 12903 15899 12909
rect 15841 12900 15853 12903
rect 12768 12872 15056 12900
rect 15120 12872 15853 12900
rect 12768 12860 12774 12872
rect 12342 12832 12348 12844
rect 11480 12804 12348 12832
rect 11480 12792 11486 12804
rect 12342 12792 12348 12804
rect 12400 12792 12406 12844
rect 12529 12835 12587 12841
rect 12529 12801 12541 12835
rect 12575 12832 12587 12835
rect 12618 12832 12624 12844
rect 12575 12804 12624 12832
rect 12575 12801 12587 12804
rect 12529 12795 12587 12801
rect 12618 12792 12624 12804
rect 12676 12792 12682 12844
rect 14550 12792 14556 12844
rect 14608 12832 14614 12844
rect 15120 12841 15148 12872
rect 15841 12869 15853 12872
rect 15887 12900 15899 12903
rect 16298 12900 16304 12912
rect 15887 12872 16304 12900
rect 15887 12869 15899 12872
rect 15841 12863 15899 12869
rect 16298 12860 16304 12872
rect 16356 12860 16362 12912
rect 15105 12835 15163 12841
rect 15105 12832 15117 12835
rect 14608 12804 15117 12832
rect 14608 12792 14614 12804
rect 15105 12801 15117 12804
rect 15151 12801 15163 12835
rect 15105 12795 15163 12801
rect 15286 12792 15292 12844
rect 15344 12792 15350 12844
rect 15470 12792 15476 12844
rect 15528 12792 15534 12844
rect 15562 12792 15568 12844
rect 15620 12832 15626 12844
rect 15657 12835 15715 12841
rect 15657 12832 15669 12835
rect 15620 12804 15669 12832
rect 15620 12792 15626 12804
rect 15657 12801 15669 12804
rect 15703 12801 15715 12835
rect 15657 12795 15715 12801
rect 15746 12792 15752 12844
rect 15804 12792 15810 12844
rect 18046 12792 18052 12844
rect 18104 12792 18110 12844
rect 18156 12832 18184 12940
rect 20622 12928 20628 12980
rect 20680 12968 20686 12980
rect 20680 12940 21128 12968
rect 20680 12928 20686 12940
rect 18230 12860 18236 12912
rect 18288 12900 18294 12912
rect 19245 12903 19303 12909
rect 19245 12900 19257 12903
rect 18288 12872 19257 12900
rect 18288 12860 18294 12872
rect 19245 12869 19257 12872
rect 19291 12869 19303 12903
rect 20070 12900 20076 12912
rect 19245 12863 19303 12869
rect 19352 12872 20076 12900
rect 18414 12832 18420 12844
rect 18156 12804 18420 12832
rect 18414 12792 18420 12804
rect 18472 12792 18478 12844
rect 18506 12792 18512 12844
rect 18564 12832 18570 12844
rect 19352 12832 19380 12872
rect 20070 12860 20076 12872
rect 20128 12860 20134 12912
rect 21100 12900 21128 12940
rect 21266 12928 21272 12980
rect 21324 12928 21330 12980
rect 22738 12928 22744 12980
rect 22796 12968 22802 12980
rect 23290 12968 23296 12980
rect 22796 12940 23296 12968
rect 22796 12928 22802 12940
rect 23290 12928 23296 12940
rect 23348 12968 23354 12980
rect 23385 12971 23443 12977
rect 23385 12968 23397 12971
rect 23348 12940 23397 12968
rect 23348 12928 23354 12940
rect 23385 12937 23397 12940
rect 23431 12937 23443 12971
rect 23385 12931 23443 12937
rect 22189 12903 22247 12909
rect 22189 12900 22201 12903
rect 21100 12872 22201 12900
rect 22189 12869 22201 12872
rect 22235 12869 22247 12903
rect 22189 12863 22247 12869
rect 22370 12860 22376 12912
rect 22428 12900 22434 12912
rect 22428 12872 23796 12900
rect 22428 12860 22434 12872
rect 18564 12804 19380 12832
rect 18564 12792 18570 12804
rect 20898 12792 20904 12844
rect 20956 12792 20962 12844
rect 21818 12792 21824 12844
rect 21876 12792 21882 12844
rect 22002 12792 22008 12844
rect 22060 12792 22066 12844
rect 23768 12841 23796 12872
rect 23385 12835 23443 12841
rect 23385 12832 23397 12835
rect 22112 12804 23397 12832
rect 2041 12767 2099 12773
rect 2041 12733 2053 12767
rect 2087 12764 2099 12767
rect 2222 12764 2228 12776
rect 2087 12736 2228 12764
rect 2087 12733 2099 12736
rect 2041 12727 2099 12733
rect 2222 12724 2228 12736
rect 2280 12724 2286 12776
rect 5350 12724 5356 12776
rect 5408 12724 5414 12776
rect 8036 12764 8064 12792
rect 8757 12767 8815 12773
rect 8757 12764 8769 12767
rect 8036 12736 8769 12764
rect 8757 12733 8769 12736
rect 8803 12733 8815 12767
rect 8757 12727 8815 12733
rect 9677 12767 9735 12773
rect 9677 12733 9689 12767
rect 9723 12764 9735 12767
rect 9766 12764 9772 12776
rect 9723 12736 9772 12764
rect 9723 12733 9735 12736
rect 9677 12727 9735 12733
rect 9766 12724 9772 12736
rect 9824 12724 9830 12776
rect 15194 12724 15200 12776
rect 15252 12764 15258 12776
rect 15381 12767 15439 12773
rect 15381 12764 15393 12767
rect 15252 12736 15393 12764
rect 15252 12724 15258 12736
rect 15381 12733 15393 12736
rect 15427 12733 15439 12767
rect 15381 12727 15439 12733
rect 17773 12767 17831 12773
rect 17773 12733 17785 12767
rect 17819 12764 17831 12767
rect 17862 12764 17868 12776
rect 17819 12736 17868 12764
rect 17819 12733 17831 12736
rect 17773 12727 17831 12733
rect 17862 12724 17868 12736
rect 17920 12764 17926 12776
rect 18325 12767 18383 12773
rect 18325 12764 18337 12767
rect 17920 12736 18337 12764
rect 17920 12724 17926 12736
rect 18325 12733 18337 12736
rect 18371 12733 18383 12767
rect 18432 12764 18460 12792
rect 19150 12764 19156 12776
rect 18432 12736 19156 12764
rect 18325 12727 18383 12733
rect 19150 12724 19156 12736
rect 19208 12724 19214 12776
rect 19518 12724 19524 12776
rect 19576 12724 19582 12776
rect 19794 12724 19800 12776
rect 19852 12724 19858 12776
rect 20806 12724 20812 12776
rect 20864 12764 20870 12776
rect 22112 12764 22140 12804
rect 23385 12801 23397 12804
rect 23431 12801 23443 12835
rect 23385 12795 23443 12801
rect 23753 12835 23811 12841
rect 23753 12801 23765 12835
rect 23799 12832 23811 12835
rect 25774 12832 25780 12844
rect 23799 12804 25780 12832
rect 23799 12801 23811 12804
rect 23753 12795 23811 12801
rect 25774 12792 25780 12804
rect 25832 12792 25838 12844
rect 20864 12736 22140 12764
rect 23201 12767 23259 12773
rect 20864 12724 20870 12736
rect 23201 12733 23213 12767
rect 23247 12733 23259 12767
rect 23201 12727 23259 12733
rect 11790 12656 11796 12708
rect 11848 12696 11854 12708
rect 17034 12696 17040 12708
rect 11848 12668 12204 12696
rect 11848 12656 11854 12668
rect 2222 12588 2228 12640
rect 2280 12588 2286 12640
rect 12066 12588 12072 12640
rect 12124 12588 12130 12640
rect 12176 12628 12204 12668
rect 16776 12668 17040 12696
rect 16776 12628 16804 12668
rect 17034 12656 17040 12668
rect 17092 12656 17098 12708
rect 18874 12656 18880 12708
rect 18932 12656 18938 12708
rect 19334 12696 19340 12708
rect 18984 12668 19340 12696
rect 12176 12600 16804 12628
rect 16850 12588 16856 12640
rect 16908 12628 16914 12640
rect 17865 12631 17923 12637
rect 17865 12628 17877 12631
rect 16908 12600 17877 12628
rect 16908 12588 16914 12600
rect 17865 12597 17877 12600
rect 17911 12597 17923 12631
rect 17865 12591 17923 12597
rect 17957 12631 18015 12637
rect 17957 12597 17969 12631
rect 18003 12628 18015 12631
rect 18984 12628 19012 12668
rect 19334 12656 19340 12668
rect 19392 12656 19398 12708
rect 22278 12656 22284 12708
rect 22336 12696 22342 12708
rect 23216 12696 23244 12727
rect 23474 12696 23480 12708
rect 22336 12668 23480 12696
rect 22336 12656 22342 12668
rect 23474 12656 23480 12668
rect 23532 12656 23538 12708
rect 18003 12600 19012 12628
rect 18003 12597 18015 12600
rect 17957 12591 18015 12597
rect 19150 12588 19156 12640
rect 19208 12628 19214 12640
rect 19245 12631 19303 12637
rect 19245 12628 19257 12631
rect 19208 12600 19257 12628
rect 19208 12588 19214 12600
rect 19245 12597 19257 12600
rect 19291 12597 19303 12631
rect 19245 12591 19303 12597
rect 19429 12631 19487 12637
rect 19429 12597 19441 12631
rect 19475 12628 19487 12631
rect 22094 12628 22100 12640
rect 19475 12600 22100 12628
rect 19475 12597 19487 12600
rect 19429 12591 19487 12597
rect 22094 12588 22100 12600
rect 22152 12588 22158 12640
rect 1104 12538 28152 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 28152 12538
rect 1104 12464 28152 12486
rect 16206 12384 16212 12436
rect 16264 12424 16270 12436
rect 16264 12396 16988 12424
rect 16264 12384 16270 12396
rect 3234 12316 3240 12368
rect 3292 12356 3298 12368
rect 4617 12359 4675 12365
rect 3292 12328 4016 12356
rect 3292 12316 3298 12328
rect 3050 12248 3056 12300
rect 3108 12288 3114 12300
rect 3145 12291 3203 12297
rect 3145 12288 3157 12291
rect 3108 12260 3157 12288
rect 3108 12248 3114 12260
rect 3145 12257 3157 12260
rect 3191 12288 3203 12291
rect 3191 12260 3740 12288
rect 3191 12257 3203 12260
rect 3145 12251 3203 12257
rect 3234 12180 3240 12232
rect 3292 12180 3298 12232
rect 3712 12222 3740 12260
rect 3988 12229 4016 12328
rect 4617 12325 4629 12359
rect 4663 12325 4675 12359
rect 4617 12319 4675 12325
rect 5537 12359 5595 12365
rect 5537 12325 5549 12359
rect 5583 12356 5595 12359
rect 7374 12356 7380 12368
rect 5583 12328 7380 12356
rect 5583 12325 5595 12328
rect 5537 12319 5595 12325
rect 4632 12288 4660 12319
rect 7374 12316 7380 12328
rect 7432 12316 7438 12368
rect 15562 12356 15568 12368
rect 12176 12328 15568 12356
rect 5350 12288 5356 12300
rect 4632 12260 5356 12288
rect 5350 12248 5356 12260
rect 5408 12288 5414 12300
rect 5408 12260 5488 12288
rect 5408 12248 5414 12260
rect 3789 12223 3847 12229
rect 3789 12222 3801 12223
rect 3712 12194 3801 12222
rect 3789 12189 3801 12194
rect 3835 12189 3847 12223
rect 3789 12183 3847 12189
rect 3973 12223 4031 12229
rect 3973 12189 3985 12223
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 4525 12223 4583 12229
rect 4525 12189 4537 12223
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 3881 12155 3939 12161
rect 3881 12121 3893 12155
rect 3927 12152 3939 12155
rect 4249 12155 4307 12161
rect 4249 12152 4261 12155
rect 3927 12124 4261 12152
rect 3927 12121 3939 12124
rect 3881 12115 3939 12121
rect 4249 12121 4261 12124
rect 4295 12121 4307 12155
rect 4249 12115 4307 12121
rect 4540 12096 4568 12183
rect 4706 12180 4712 12232
rect 4764 12180 4770 12232
rect 4798 12180 4804 12232
rect 4856 12220 4862 12232
rect 5460 12229 5488 12260
rect 8294 12248 8300 12300
rect 8352 12248 8358 12300
rect 4893 12223 4951 12229
rect 4893 12220 4905 12223
rect 4856 12192 4905 12220
rect 4856 12180 4862 12192
rect 4893 12189 4905 12192
rect 4939 12189 4951 12223
rect 4893 12183 4951 12189
rect 5445 12223 5503 12229
rect 5445 12189 5457 12223
rect 5491 12189 5503 12223
rect 5445 12183 5503 12189
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 5629 12223 5687 12229
rect 5629 12220 5641 12223
rect 5592 12192 5641 12220
rect 5592 12180 5598 12192
rect 5629 12189 5641 12192
rect 5675 12189 5687 12223
rect 5629 12183 5687 12189
rect 6178 12180 6184 12232
rect 6236 12180 6242 12232
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12220 6607 12223
rect 6638 12220 6644 12232
rect 6595 12192 6644 12220
rect 6595 12189 6607 12192
rect 6549 12183 6607 12189
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 7098 12180 7104 12232
rect 7156 12220 7162 12232
rect 7377 12223 7435 12229
rect 7377 12220 7389 12223
rect 7156 12192 7389 12220
rect 7156 12180 7162 12192
rect 7377 12189 7389 12192
rect 7423 12189 7435 12223
rect 7377 12183 7435 12189
rect 7193 12155 7251 12161
rect 7193 12121 7205 12155
rect 7239 12152 7251 12155
rect 7484 12152 7512 12206
rect 11330 12180 11336 12232
rect 11388 12180 11394 12232
rect 12176 12229 12204 12328
rect 15562 12316 15568 12328
rect 15620 12356 15626 12368
rect 16482 12356 16488 12368
rect 15620 12328 16488 12356
rect 15620 12316 15626 12328
rect 16482 12316 16488 12328
rect 16540 12316 16546 12368
rect 16574 12316 16580 12368
rect 16632 12316 16638 12368
rect 12250 12248 12256 12300
rect 12308 12248 12314 12300
rect 12434 12248 12440 12300
rect 12492 12248 12498 12300
rect 12526 12248 12532 12300
rect 12584 12288 12590 12300
rect 12713 12291 12771 12297
rect 12713 12288 12725 12291
rect 12584 12260 12725 12288
rect 12584 12248 12590 12260
rect 12713 12257 12725 12260
rect 12759 12257 12771 12291
rect 12713 12251 12771 12257
rect 12802 12248 12808 12300
rect 12860 12288 12866 12300
rect 16393 12291 16451 12297
rect 12860 12260 12940 12288
rect 12860 12248 12866 12260
rect 12912 12229 12940 12260
rect 16393 12257 16405 12291
rect 16439 12288 16451 12291
rect 16850 12288 16856 12300
rect 16439 12260 16856 12288
rect 16439 12257 16451 12260
rect 16393 12251 16451 12257
rect 16850 12248 16856 12260
rect 16908 12248 16914 12300
rect 16960 12288 16988 12396
rect 18782 12384 18788 12436
rect 18840 12424 18846 12436
rect 18840 12396 19288 12424
rect 18840 12384 18846 12396
rect 18046 12316 18052 12368
rect 18104 12356 18110 12368
rect 19150 12356 19156 12368
rect 18104 12328 19156 12356
rect 18104 12316 18110 12328
rect 19150 12316 19156 12328
rect 19208 12316 19214 12368
rect 19260 12356 19288 12396
rect 19334 12384 19340 12436
rect 19392 12424 19398 12436
rect 19521 12427 19579 12433
rect 19521 12424 19533 12427
rect 19392 12396 19533 12424
rect 19392 12384 19398 12396
rect 19260 12328 19380 12356
rect 19352 12300 19380 12328
rect 18506 12288 18512 12300
rect 16960 12260 18512 12288
rect 11609 12223 11667 12229
rect 11609 12189 11621 12223
rect 11655 12220 11667 12223
rect 11885 12223 11943 12229
rect 11885 12220 11897 12223
rect 11655 12192 11897 12220
rect 11655 12189 11667 12192
rect 11609 12183 11667 12189
rect 11885 12189 11897 12192
rect 11931 12189 11943 12223
rect 11885 12183 11943 12189
rect 12161 12223 12219 12229
rect 12161 12189 12173 12223
rect 12207 12189 12219 12223
rect 12161 12183 12219 12189
rect 12345 12223 12403 12229
rect 12345 12189 12357 12223
rect 12391 12220 12403 12223
rect 12621 12223 12679 12229
rect 12391 12192 12572 12220
rect 12391 12189 12403 12192
rect 12345 12183 12403 12189
rect 7742 12152 7748 12164
rect 7239 12124 7748 12152
rect 7239 12121 7251 12124
rect 7193 12115 7251 12121
rect 7742 12112 7748 12124
rect 7800 12112 7806 12164
rect 3605 12087 3663 12093
rect 3605 12053 3617 12087
rect 3651 12084 3663 12087
rect 4522 12084 4528 12096
rect 3651 12056 4528 12084
rect 3651 12053 3663 12056
rect 3605 12047 3663 12053
rect 4522 12044 4528 12056
rect 4580 12044 4586 12096
rect 11146 12044 11152 12096
rect 11204 12044 11210 12096
rect 11514 12044 11520 12096
rect 11572 12044 11578 12096
rect 12544 12084 12572 12192
rect 12621 12189 12633 12223
rect 12667 12189 12679 12223
rect 12621 12183 12679 12189
rect 12897 12223 12955 12229
rect 12897 12189 12909 12223
rect 12943 12189 12955 12223
rect 12897 12183 12955 12189
rect 12636 12152 12664 12183
rect 16022 12180 16028 12232
rect 16080 12220 16086 12232
rect 16117 12223 16175 12229
rect 16117 12220 16129 12223
rect 16080 12192 16129 12220
rect 16080 12180 16086 12192
rect 16117 12189 16129 12192
rect 16163 12189 16175 12223
rect 16117 12183 16175 12189
rect 16298 12180 16304 12232
rect 16356 12180 16362 12232
rect 16960 12229 16988 12260
rect 18506 12248 18512 12260
rect 18564 12248 18570 12300
rect 19334 12248 19340 12300
rect 19392 12248 19398 12300
rect 16577 12223 16635 12229
rect 16577 12189 16589 12223
rect 16623 12189 16635 12223
rect 16577 12183 16635 12189
rect 16945 12223 17003 12229
rect 16945 12189 16957 12223
rect 16991 12189 17003 12223
rect 16945 12183 17003 12189
rect 12802 12152 12808 12164
rect 12636 12124 12808 12152
rect 12802 12112 12808 12124
rect 12860 12152 12866 12164
rect 13262 12152 13268 12164
rect 12860 12124 13268 12152
rect 12860 12112 12866 12124
rect 13262 12112 13268 12124
rect 13320 12112 13326 12164
rect 16592 12152 16620 12183
rect 17126 12180 17132 12232
rect 17184 12180 17190 12232
rect 17218 12180 17224 12232
rect 17276 12180 17282 12232
rect 18046 12180 18052 12232
rect 18104 12220 18110 12232
rect 18141 12223 18199 12229
rect 18141 12220 18153 12223
rect 18104 12192 18153 12220
rect 18104 12180 18110 12192
rect 18141 12189 18153 12192
rect 18187 12189 18199 12223
rect 18141 12183 18199 12189
rect 18414 12180 18420 12232
rect 18472 12220 18478 12232
rect 18601 12223 18659 12229
rect 18601 12220 18613 12223
rect 18472 12192 18613 12220
rect 18472 12180 18478 12192
rect 18601 12189 18613 12192
rect 18647 12189 18659 12223
rect 18601 12183 18659 12189
rect 17144 12152 17172 12180
rect 16592 12124 17172 12152
rect 18616 12152 18644 12183
rect 18782 12180 18788 12232
rect 18840 12220 18846 12232
rect 18877 12223 18935 12229
rect 18877 12220 18889 12223
rect 18840 12192 18889 12220
rect 18840 12180 18846 12192
rect 18877 12189 18889 12192
rect 18923 12189 18935 12223
rect 18877 12183 18935 12189
rect 19061 12223 19119 12229
rect 19061 12189 19073 12223
rect 19107 12189 19119 12223
rect 19061 12183 19119 12189
rect 19076 12152 19104 12183
rect 19150 12180 19156 12232
rect 19208 12220 19214 12232
rect 19444 12229 19472 12396
rect 19521 12393 19533 12396
rect 19567 12393 19579 12427
rect 19521 12387 19579 12393
rect 19886 12384 19892 12436
rect 19944 12424 19950 12436
rect 21082 12424 21088 12436
rect 19944 12396 21088 12424
rect 19944 12384 19950 12396
rect 21082 12384 21088 12396
rect 21140 12384 21146 12436
rect 21637 12427 21695 12433
rect 21637 12393 21649 12427
rect 21683 12424 21695 12427
rect 22002 12424 22008 12436
rect 21683 12396 22008 12424
rect 21683 12393 21695 12396
rect 21637 12387 21695 12393
rect 22002 12384 22008 12396
rect 22060 12384 22066 12436
rect 19904 12356 19932 12384
rect 21177 12359 21235 12365
rect 19904 12328 20024 12356
rect 19886 12288 19892 12300
rect 19720 12260 19892 12288
rect 19720 12229 19748 12260
rect 19886 12248 19892 12260
rect 19944 12248 19950 12300
rect 19996 12229 20024 12328
rect 21177 12325 21189 12359
rect 21223 12356 21235 12359
rect 21818 12356 21824 12368
rect 21223 12328 21824 12356
rect 21223 12325 21235 12328
rect 21177 12319 21235 12325
rect 21818 12316 21824 12328
rect 21876 12316 21882 12368
rect 20530 12248 20536 12300
rect 20588 12248 20594 12300
rect 20714 12248 20720 12300
rect 20772 12288 20778 12300
rect 21266 12288 21272 12300
rect 20772 12260 21272 12288
rect 20772 12248 20778 12260
rect 19245 12223 19303 12229
rect 19245 12220 19257 12223
rect 19208 12192 19257 12220
rect 19208 12180 19214 12192
rect 19245 12189 19257 12192
rect 19291 12189 19303 12223
rect 19245 12183 19303 12189
rect 19429 12223 19487 12229
rect 19429 12189 19441 12223
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 19705 12223 19763 12229
rect 19705 12189 19717 12223
rect 19751 12189 19763 12223
rect 19705 12183 19763 12189
rect 19981 12223 20039 12229
rect 19981 12189 19993 12223
rect 20027 12189 20039 12223
rect 19981 12183 20039 12189
rect 18616 12124 19104 12152
rect 12618 12084 12624 12096
rect 12544 12056 12624 12084
rect 12618 12044 12624 12056
rect 12676 12084 12682 12096
rect 12894 12084 12900 12096
rect 12676 12056 12900 12084
rect 12676 12044 12682 12056
rect 12894 12044 12900 12056
rect 12952 12084 12958 12096
rect 13081 12087 13139 12093
rect 13081 12084 13093 12087
rect 12952 12056 13093 12084
rect 12952 12044 12958 12056
rect 13081 12053 13093 12056
rect 13127 12053 13139 12087
rect 13081 12047 13139 12053
rect 13170 12044 13176 12096
rect 13228 12084 13234 12096
rect 16485 12087 16543 12093
rect 16485 12084 16497 12087
rect 13228 12056 16497 12084
rect 13228 12044 13234 12056
rect 16485 12053 16497 12056
rect 16531 12053 16543 12087
rect 16485 12047 16543 12053
rect 16574 12044 16580 12096
rect 16632 12084 16638 12096
rect 16761 12087 16819 12093
rect 16761 12084 16773 12087
rect 16632 12056 16773 12084
rect 16632 12044 16638 12056
rect 16761 12053 16773 12056
rect 16807 12053 16819 12087
rect 16761 12047 16819 12053
rect 17034 12044 17040 12096
rect 17092 12084 17098 12096
rect 17129 12087 17187 12093
rect 17129 12084 17141 12087
rect 17092 12056 17141 12084
rect 17092 12044 17098 12056
rect 17129 12053 17141 12056
rect 17175 12053 17187 12087
rect 17129 12047 17187 12053
rect 18230 12044 18236 12096
rect 18288 12044 18294 12096
rect 18690 12044 18696 12096
rect 18748 12044 18754 12096
rect 18969 12087 19027 12093
rect 18969 12053 18981 12087
rect 19015 12084 19027 12087
rect 19058 12084 19064 12096
rect 19015 12056 19064 12084
rect 19015 12053 19027 12056
rect 18969 12047 19027 12053
rect 19058 12044 19064 12056
rect 19116 12044 19122 12096
rect 19260 12084 19288 12183
rect 20254 12180 20260 12232
rect 20312 12180 20318 12232
rect 20441 12223 20499 12229
rect 20441 12189 20453 12223
rect 20487 12189 20499 12223
rect 20441 12183 20499 12189
rect 19337 12155 19395 12161
rect 19337 12121 19349 12155
rect 19383 12152 19395 12155
rect 19794 12152 19800 12164
rect 19383 12124 19800 12152
rect 19383 12121 19395 12124
rect 19337 12115 19395 12121
rect 19794 12112 19800 12124
rect 19852 12112 19858 12164
rect 19889 12155 19947 12161
rect 19889 12121 19901 12155
rect 19935 12152 19947 12155
rect 20272 12152 20300 12180
rect 19935 12124 20300 12152
rect 19935 12121 19947 12124
rect 19889 12115 19947 12121
rect 20073 12087 20131 12093
rect 20073 12084 20085 12087
rect 19260 12056 20085 12084
rect 20073 12053 20085 12056
rect 20119 12053 20131 12087
rect 20456 12084 20484 12183
rect 20622 12180 20628 12232
rect 20680 12180 20686 12232
rect 20806 12180 20812 12232
rect 20864 12180 20870 12232
rect 21008 12229 21036 12260
rect 21266 12248 21272 12260
rect 21324 12248 21330 12300
rect 20993 12223 21051 12229
rect 20993 12189 21005 12223
rect 21039 12189 21051 12223
rect 20993 12183 21051 12189
rect 21082 12180 21088 12232
rect 21140 12220 21146 12232
rect 21177 12223 21235 12229
rect 21177 12220 21189 12223
rect 21140 12192 21189 12220
rect 21140 12180 21146 12192
rect 21177 12189 21189 12192
rect 21223 12189 21235 12223
rect 21177 12183 21235 12189
rect 21453 12223 21511 12229
rect 21453 12189 21465 12223
rect 21499 12189 21511 12223
rect 21453 12183 21511 12189
rect 21192 12152 21220 12183
rect 21468 12152 21496 12183
rect 21192 12124 21496 12152
rect 21542 12112 21548 12164
rect 21600 12152 21606 12164
rect 23198 12152 23204 12164
rect 21600 12124 23204 12152
rect 21600 12112 21606 12124
rect 23198 12112 23204 12124
rect 23256 12112 23262 12164
rect 22462 12084 22468 12096
rect 20456 12056 22468 12084
rect 20073 12047 20131 12053
rect 22462 12044 22468 12056
rect 22520 12084 22526 12096
rect 23106 12084 23112 12096
rect 22520 12056 23112 12084
rect 22520 12044 22526 12056
rect 23106 12044 23112 12056
rect 23164 12044 23170 12096
rect 1104 11994 28152 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 28152 11994
rect 1104 11920 28152 11942
rect 3234 11840 3240 11892
rect 3292 11880 3298 11892
rect 3697 11883 3755 11889
rect 3697 11880 3709 11883
rect 3292 11852 3709 11880
rect 3292 11840 3298 11852
rect 3697 11849 3709 11852
rect 3743 11849 3755 11883
rect 3697 11843 3755 11849
rect 7653 11883 7711 11889
rect 7653 11849 7665 11883
rect 7699 11880 7711 11883
rect 8202 11880 8208 11892
rect 7699 11852 8208 11880
rect 7699 11849 7711 11852
rect 7653 11843 7711 11849
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 11330 11840 11336 11892
rect 11388 11840 11394 11892
rect 11514 11840 11520 11892
rect 11572 11840 11578 11892
rect 11808 11852 13768 11880
rect 2222 11772 2228 11824
rect 2280 11812 2286 11824
rect 4798 11812 4804 11824
rect 2280 11784 3096 11812
rect 2280 11772 2286 11784
rect 842 11704 848 11756
rect 900 11744 906 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 900 11716 1409 11744
rect 900 11704 906 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 2314 11704 2320 11756
rect 2372 11744 2378 11756
rect 3068 11753 3096 11784
rect 4080 11784 4804 11812
rect 4080 11756 4108 11784
rect 4798 11772 4804 11784
rect 4856 11812 4862 11824
rect 4856 11784 5304 11812
rect 4856 11772 4862 11784
rect 2869 11747 2927 11753
rect 2869 11744 2881 11747
rect 2372 11716 2881 11744
rect 2372 11704 2378 11716
rect 2869 11713 2881 11716
rect 2915 11713 2927 11747
rect 2869 11707 2927 11713
rect 3053 11747 3111 11753
rect 3053 11713 3065 11747
rect 3099 11713 3111 11747
rect 4062 11744 4068 11756
rect 3053 11707 3111 11713
rect 3344 11716 4068 11744
rect 3344 11688 3372 11716
rect 4062 11704 4068 11716
rect 4120 11704 4126 11756
rect 4617 11747 4675 11753
rect 4617 11713 4629 11747
rect 4663 11713 4675 11747
rect 4617 11707 4675 11713
rect 1673 11679 1731 11685
rect 1673 11645 1685 11679
rect 1719 11645 1731 11679
rect 1673 11639 1731 11645
rect 2961 11679 3019 11685
rect 2961 11645 2973 11679
rect 3007 11676 3019 11679
rect 3237 11679 3295 11685
rect 3237 11676 3249 11679
rect 3007 11648 3249 11676
rect 3007 11645 3019 11648
rect 2961 11639 3019 11645
rect 3237 11645 3249 11648
rect 3283 11645 3295 11679
rect 3237 11639 3295 11645
rect 1688 11608 1716 11639
rect 3326 11636 3332 11688
rect 3384 11636 3390 11688
rect 3421 11679 3479 11685
rect 3421 11645 3433 11679
rect 3467 11645 3479 11679
rect 3421 11639 3479 11645
rect 2774 11608 2780 11620
rect 1688 11580 2780 11608
rect 2774 11568 2780 11580
rect 2832 11608 2838 11620
rect 3436 11608 3464 11639
rect 3510 11636 3516 11688
rect 3568 11636 3574 11688
rect 4522 11636 4528 11688
rect 4580 11636 4586 11688
rect 4632 11676 4660 11707
rect 4706 11704 4712 11756
rect 4764 11744 4770 11756
rect 5074 11744 5080 11756
rect 4764 11716 5080 11744
rect 4764 11704 4770 11716
rect 5074 11704 5080 11716
rect 5132 11704 5138 11756
rect 5276 11753 5304 11784
rect 10502 11772 10508 11824
rect 10560 11812 10566 11824
rect 10965 11815 11023 11821
rect 10965 11812 10977 11815
rect 10560 11784 10977 11812
rect 10560 11772 10566 11784
rect 10965 11781 10977 11784
rect 11011 11812 11023 11815
rect 11011 11784 11560 11812
rect 11011 11781 11023 11784
rect 10965 11775 11023 11781
rect 5261 11747 5319 11753
rect 5261 11713 5273 11747
rect 5307 11713 5319 11747
rect 5261 11707 5319 11713
rect 7098 11704 7104 11756
rect 7156 11744 7162 11756
rect 7561 11747 7619 11753
rect 7561 11744 7573 11747
rect 7156 11716 7573 11744
rect 7156 11704 7162 11716
rect 7561 11713 7573 11716
rect 7607 11713 7619 11747
rect 7561 11707 7619 11713
rect 7742 11704 7748 11756
rect 7800 11704 7806 11756
rect 10870 11704 10876 11756
rect 10928 11704 10934 11756
rect 11149 11747 11207 11753
rect 11149 11713 11161 11747
rect 11195 11713 11207 11747
rect 11149 11707 11207 11713
rect 5169 11679 5227 11685
rect 5169 11676 5181 11679
rect 4632 11648 5181 11676
rect 5169 11645 5181 11648
rect 5215 11645 5227 11679
rect 5169 11639 5227 11645
rect 2832 11580 3464 11608
rect 2832 11568 2838 11580
rect 3436 11540 3464 11580
rect 4985 11611 5043 11617
rect 4985 11577 4997 11611
rect 5031 11608 5043 11611
rect 5534 11608 5540 11620
rect 5031 11580 5540 11608
rect 5031 11577 5043 11580
rect 4985 11571 5043 11577
rect 5534 11568 5540 11580
rect 5592 11568 5598 11620
rect 6730 11540 6736 11552
rect 3436 11512 6736 11540
rect 6730 11500 6736 11512
rect 6788 11500 6794 11552
rect 11164 11540 11192 11707
rect 11532 11608 11560 11784
rect 11698 11704 11704 11756
rect 11756 11704 11762 11756
rect 11808 11753 11836 11852
rect 12526 11812 12532 11824
rect 12084 11784 12532 11812
rect 11793 11747 11851 11753
rect 11793 11713 11805 11747
rect 11839 11713 11851 11747
rect 11793 11707 11851 11713
rect 11974 11704 11980 11756
rect 12032 11704 12038 11756
rect 12084 11753 12112 11784
rect 12526 11772 12532 11784
rect 12584 11772 12590 11824
rect 12069 11747 12127 11753
rect 12069 11713 12081 11747
rect 12115 11713 12127 11747
rect 12069 11707 12127 11713
rect 12084 11608 12112 11707
rect 12158 11704 12164 11756
rect 12216 11704 12222 11756
rect 12250 11704 12256 11756
rect 12308 11704 12314 11756
rect 12345 11747 12403 11753
rect 12345 11713 12357 11747
rect 12391 11744 12403 11747
rect 12434 11744 12440 11756
rect 12391 11716 12440 11744
rect 12391 11713 12403 11716
rect 12345 11707 12403 11713
rect 12434 11704 12440 11716
rect 12492 11744 12498 11756
rect 12621 11747 12679 11753
rect 12621 11744 12633 11747
rect 12492 11716 12633 11744
rect 12492 11704 12498 11716
rect 12621 11713 12633 11716
rect 12667 11713 12679 11747
rect 12621 11707 12679 11713
rect 13740 11676 13768 11852
rect 13814 11840 13820 11892
rect 13872 11880 13878 11892
rect 16206 11880 16212 11892
rect 13872 11852 16212 11880
rect 13872 11840 13878 11852
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 16298 11840 16304 11892
rect 16356 11880 16362 11892
rect 16393 11883 16451 11889
rect 16393 11880 16405 11883
rect 16356 11852 16405 11880
rect 16356 11840 16362 11852
rect 16393 11849 16405 11852
rect 16439 11849 16451 11883
rect 16393 11843 16451 11849
rect 19337 11883 19395 11889
rect 19337 11849 19349 11883
rect 19383 11880 19395 11883
rect 19426 11880 19432 11892
rect 19383 11852 19432 11880
rect 19383 11849 19395 11852
rect 19337 11843 19395 11849
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 19518 11840 19524 11892
rect 19576 11880 19582 11892
rect 20162 11880 20168 11892
rect 19576 11852 20168 11880
rect 19576 11840 19582 11852
rect 20162 11840 20168 11852
rect 20220 11880 20226 11892
rect 21085 11883 21143 11889
rect 21085 11880 21097 11883
rect 20220 11852 21097 11880
rect 20220 11840 20226 11852
rect 21085 11849 21097 11852
rect 21131 11849 21143 11883
rect 21085 11843 21143 11849
rect 22830 11840 22836 11892
rect 22888 11880 22894 11892
rect 23017 11883 23075 11889
rect 23017 11880 23029 11883
rect 22888 11852 23029 11880
rect 22888 11840 22894 11852
rect 23017 11849 23029 11852
rect 23063 11849 23075 11883
rect 23017 11843 23075 11849
rect 23290 11840 23296 11892
rect 23348 11840 23354 11892
rect 23474 11840 23480 11892
rect 23532 11880 23538 11892
rect 23532 11852 23704 11880
rect 23532 11840 23538 11852
rect 17034 11812 17040 11824
rect 15488 11784 17040 11812
rect 14734 11704 14740 11756
rect 14792 11744 14798 11756
rect 15488 11753 15516 11784
rect 17034 11772 17040 11784
rect 17092 11772 17098 11824
rect 17770 11772 17776 11824
rect 17828 11812 17834 11824
rect 23308 11812 23336 11840
rect 23385 11815 23443 11821
rect 23385 11812 23397 11815
rect 17828 11784 19932 11812
rect 17828 11772 17834 11784
rect 15473 11747 15531 11753
rect 15473 11744 15485 11747
rect 14792 11716 15485 11744
rect 14792 11704 14798 11716
rect 15473 11713 15485 11716
rect 15519 11713 15531 11747
rect 15473 11707 15531 11713
rect 15562 11704 15568 11756
rect 15620 11704 15626 11756
rect 15749 11747 15807 11753
rect 15749 11713 15761 11747
rect 15795 11713 15807 11747
rect 15749 11707 15807 11713
rect 15764 11676 15792 11707
rect 15838 11704 15844 11756
rect 15896 11704 15902 11756
rect 15930 11704 15936 11756
rect 15988 11744 15994 11756
rect 16117 11747 16175 11753
rect 16117 11744 16129 11747
rect 15988 11716 16129 11744
rect 15988 11704 15994 11716
rect 16117 11713 16129 11716
rect 16163 11713 16175 11747
rect 16117 11707 16175 11713
rect 16209 11747 16267 11753
rect 16209 11713 16221 11747
rect 16255 11713 16267 11747
rect 16209 11707 16267 11713
rect 16485 11747 16543 11753
rect 16485 11713 16497 11747
rect 16531 11744 16543 11747
rect 16574 11744 16580 11756
rect 16531 11716 16580 11744
rect 16531 11713 16543 11716
rect 16485 11707 16543 11713
rect 13740 11648 15792 11676
rect 11532 11580 12112 11608
rect 12158 11568 12164 11620
rect 12216 11608 12222 11620
rect 12710 11608 12716 11620
rect 12216 11580 12716 11608
rect 12216 11568 12222 11580
rect 12710 11568 12716 11580
rect 12768 11568 12774 11620
rect 15764 11608 15792 11648
rect 16025 11611 16083 11617
rect 15764 11580 15976 11608
rect 13814 11540 13820 11552
rect 11164 11512 13820 11540
rect 13814 11500 13820 11512
rect 13872 11500 13878 11552
rect 15948 11540 15976 11580
rect 16025 11577 16037 11611
rect 16071 11608 16083 11611
rect 16114 11608 16120 11620
rect 16071 11580 16120 11608
rect 16071 11577 16083 11580
rect 16025 11571 16083 11577
rect 16114 11568 16120 11580
rect 16172 11608 16178 11620
rect 16224 11608 16252 11707
rect 16574 11704 16580 11716
rect 16632 11704 16638 11756
rect 16666 11704 16672 11756
rect 16724 11704 16730 11756
rect 18690 11704 18696 11756
rect 18748 11704 18754 11756
rect 18874 11704 18880 11756
rect 18932 11704 18938 11756
rect 19058 11704 19064 11756
rect 19116 11704 19122 11756
rect 19153 11747 19211 11753
rect 19153 11713 19165 11747
rect 19199 11713 19211 11747
rect 19153 11707 19211 11713
rect 16301 11679 16359 11685
rect 16301 11645 16313 11679
rect 16347 11676 16359 11679
rect 16347 11648 16528 11676
rect 16347 11645 16359 11648
rect 16301 11639 16359 11645
rect 16500 11620 16528 11648
rect 18230 11636 18236 11688
rect 18288 11676 18294 11688
rect 18969 11679 19027 11685
rect 18969 11676 18981 11679
rect 18288 11648 18981 11676
rect 18288 11636 18294 11648
rect 18969 11645 18981 11648
rect 19015 11645 19027 11679
rect 19168 11676 19196 11707
rect 19518 11704 19524 11756
rect 19576 11704 19582 11756
rect 19702 11704 19708 11756
rect 19760 11744 19766 11756
rect 19797 11747 19855 11753
rect 19797 11744 19809 11747
rect 19760 11716 19809 11744
rect 19760 11704 19766 11716
rect 19797 11713 19809 11716
rect 19843 11713 19855 11747
rect 19904 11744 19932 11784
rect 22848 11784 23397 11812
rect 22848 11756 22876 11784
rect 23385 11781 23397 11784
rect 23431 11781 23443 11815
rect 23385 11775 23443 11781
rect 19904 11716 22094 11744
rect 19797 11707 19855 11713
rect 20990 11676 20996 11688
rect 19168 11648 20996 11676
rect 18969 11639 19027 11645
rect 20990 11636 20996 11648
rect 21048 11636 21054 11688
rect 22066 11676 22094 11716
rect 22830 11704 22836 11756
rect 22888 11704 22894 11756
rect 23198 11704 23204 11756
rect 23256 11704 23262 11756
rect 23290 11704 23296 11756
rect 23348 11704 23354 11756
rect 23474 11704 23480 11756
rect 23532 11744 23538 11756
rect 23676 11753 23704 11852
rect 23569 11747 23627 11753
rect 23569 11744 23581 11747
rect 23532 11716 23581 11744
rect 23532 11704 23538 11716
rect 23569 11713 23581 11716
rect 23615 11713 23627 11747
rect 23569 11707 23627 11713
rect 23661 11747 23719 11753
rect 23661 11713 23673 11747
rect 23707 11713 23719 11747
rect 23661 11707 23719 11713
rect 24026 11676 24032 11688
rect 22066 11648 24032 11676
rect 24026 11636 24032 11648
rect 24084 11636 24090 11688
rect 16172 11580 16252 11608
rect 16172 11568 16178 11580
rect 16482 11568 16488 11620
rect 16540 11568 16546 11620
rect 18322 11568 18328 11620
rect 18380 11608 18386 11620
rect 22738 11608 22744 11620
rect 18380 11580 22744 11608
rect 18380 11568 18386 11580
rect 22738 11568 22744 11580
rect 22796 11608 22802 11620
rect 23658 11608 23664 11620
rect 22796 11580 23664 11608
rect 22796 11568 22802 11580
rect 23658 11568 23664 11580
rect 23716 11568 23722 11620
rect 17310 11540 17316 11552
rect 15948 11512 17316 11540
rect 17310 11500 17316 11512
rect 17368 11500 17374 11552
rect 18782 11500 18788 11552
rect 18840 11540 18846 11552
rect 20714 11540 20720 11552
rect 18840 11512 20720 11540
rect 18840 11500 18846 11512
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 21266 11500 21272 11552
rect 21324 11540 21330 11552
rect 23014 11540 23020 11552
rect 21324 11512 23020 11540
rect 21324 11500 21330 11512
rect 23014 11500 23020 11512
rect 23072 11500 23078 11552
rect 1104 11450 28152 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 28152 11450
rect 1104 11376 28152 11398
rect 2685 11339 2743 11345
rect 2685 11305 2697 11339
rect 2731 11336 2743 11339
rect 2958 11336 2964 11348
rect 2731 11308 2964 11336
rect 2731 11305 2743 11308
rect 2685 11299 2743 11305
rect 2958 11296 2964 11308
rect 3016 11336 3022 11348
rect 3510 11336 3516 11348
rect 3016 11308 3516 11336
rect 3016 11296 3022 11308
rect 3510 11296 3516 11308
rect 3568 11296 3574 11348
rect 10042 11296 10048 11348
rect 10100 11296 10106 11348
rect 10226 11296 10232 11348
rect 10284 11296 10290 11348
rect 10778 11296 10784 11348
rect 10836 11336 10842 11348
rect 11701 11339 11759 11345
rect 11701 11336 11713 11339
rect 10836 11308 11713 11336
rect 10836 11296 10842 11308
rect 11701 11305 11713 11308
rect 11747 11305 11759 11339
rect 11701 11299 11759 11305
rect 12066 11296 12072 11348
rect 12124 11336 12130 11348
rect 12434 11336 12440 11348
rect 12124 11308 12440 11336
rect 12124 11296 12130 11308
rect 12434 11296 12440 11308
rect 12492 11296 12498 11348
rect 12526 11296 12532 11348
rect 12584 11296 12590 11348
rect 12989 11339 13047 11345
rect 12989 11305 13001 11339
rect 13035 11336 13047 11339
rect 13170 11336 13176 11348
rect 13035 11308 13176 11336
rect 13035 11305 13047 11308
rect 12989 11299 13047 11305
rect 13170 11296 13176 11308
rect 13228 11296 13234 11348
rect 14458 11296 14464 11348
rect 14516 11336 14522 11348
rect 15105 11339 15163 11345
rect 15105 11336 15117 11339
rect 14516 11308 15117 11336
rect 14516 11296 14522 11308
rect 15105 11305 15117 11308
rect 15151 11305 15163 11339
rect 16574 11336 16580 11348
rect 15105 11299 15163 11305
rect 15764 11308 16580 11336
rect 6730 11228 6736 11280
rect 6788 11268 6794 11280
rect 11514 11268 11520 11280
rect 6788 11240 9674 11268
rect 6788 11228 6794 11240
rect 2222 11160 2228 11212
rect 2280 11160 2286 11212
rect 7190 11160 7196 11212
rect 7248 11160 7254 11212
rect 9646 11200 9674 11240
rect 10980 11240 11520 11268
rect 10134 11200 10140 11212
rect 9646 11172 10140 11200
rect 10134 11160 10140 11172
rect 10192 11200 10198 11212
rect 10980 11209 11008 11240
rect 11514 11228 11520 11240
rect 11572 11228 11578 11280
rect 11606 11228 11612 11280
rect 11664 11228 11670 11280
rect 15013 11271 15071 11277
rect 11808 11240 12434 11268
rect 10965 11203 11023 11209
rect 10965 11200 10977 11203
rect 10192 11172 10977 11200
rect 10192 11160 10198 11172
rect 2314 11092 2320 11144
rect 2372 11092 2378 11144
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11132 7159 11135
rect 7374 11132 7380 11144
rect 7147 11104 7380 11132
rect 7147 11101 7159 11104
rect 7101 11095 7159 11101
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 10502 11092 10508 11144
rect 10560 11092 10566 11144
rect 10612 11141 10640 11172
rect 10965 11169 10977 11172
rect 11011 11169 11023 11203
rect 10965 11163 11023 11169
rect 11057 11203 11115 11209
rect 11057 11169 11069 11203
rect 11103 11200 11115 11203
rect 11146 11200 11152 11212
rect 11103 11172 11152 11200
rect 11103 11169 11115 11172
rect 11057 11163 11115 11169
rect 11146 11160 11152 11172
rect 11204 11160 11210 11212
rect 11425 11203 11483 11209
rect 11425 11169 11437 11203
rect 11471 11200 11483 11203
rect 11808 11200 11836 11240
rect 11471 11172 11836 11200
rect 11471 11169 11483 11172
rect 11425 11163 11483 11169
rect 11974 11160 11980 11212
rect 12032 11160 12038 11212
rect 12406 11200 12434 11240
rect 15013 11237 15025 11271
rect 15059 11237 15071 11271
rect 15013 11231 15071 11237
rect 14918 11200 14924 11212
rect 12406 11172 12940 11200
rect 10597 11135 10655 11141
rect 10597 11101 10609 11135
rect 10643 11101 10655 11135
rect 10597 11095 10655 11101
rect 10778 11092 10784 11144
rect 10836 11092 10842 11144
rect 10870 11092 10876 11144
rect 10928 11092 10934 11144
rect 11330 11092 11336 11144
rect 11388 11092 11394 11144
rect 11839 11135 11897 11141
rect 11839 11101 11851 11135
rect 11885 11132 11897 11135
rect 11992 11132 12020 11160
rect 11885 11104 12020 11132
rect 11885 11103 11928 11104
rect 11885 11101 11897 11103
rect 11839 11095 11897 11101
rect 12250 11092 12256 11144
rect 12308 11092 12314 11144
rect 12912 11141 12940 11172
rect 14660 11172 14924 11200
rect 12345 11135 12403 11141
rect 12345 11101 12357 11135
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 12437 11135 12495 11141
rect 12437 11101 12449 11135
rect 12483 11101 12495 11135
rect 12437 11095 12495 11101
rect 12897 11135 12955 11141
rect 12897 11101 12909 11135
rect 12943 11101 12955 11135
rect 12897 11095 12955 11101
rect 6546 11024 6552 11076
rect 6604 11024 6610 11076
rect 9766 11024 9772 11076
rect 9824 11064 9830 11076
rect 9861 11067 9919 11073
rect 9861 11064 9873 11067
rect 9824 11036 9873 11064
rect 9824 11024 9830 11036
rect 9861 11033 9873 11036
rect 9907 11033 9919 11067
rect 9861 11027 9919 11033
rect 10321 11067 10379 11073
rect 10321 11033 10333 11067
rect 10367 11064 10379 11067
rect 10367 11036 10916 11064
rect 10367 11033 10379 11036
rect 10321 11027 10379 11033
rect 7098 10956 7104 11008
rect 7156 10956 7162 11008
rect 9950 10956 9956 11008
rect 10008 10996 10014 11008
rect 10061 10999 10119 11005
rect 10061 10996 10073 10999
rect 10008 10968 10073 10996
rect 10008 10956 10014 10968
rect 10061 10965 10073 10968
rect 10107 10965 10119 10999
rect 10888 10996 10916 11036
rect 11054 11024 11060 11076
rect 11112 11064 11118 11076
rect 11977 11067 12035 11073
rect 11977 11064 11989 11067
rect 11112 11036 11989 11064
rect 11112 11024 11118 11036
rect 11977 11033 11989 11036
rect 12023 11033 12035 11067
rect 11977 11027 12035 11033
rect 12066 11024 12072 11076
rect 12124 11024 12130 11076
rect 12158 11024 12164 11076
rect 12216 11064 12222 11076
rect 12360 11064 12388 11095
rect 12216 11036 12388 11064
rect 12216 11024 12222 11036
rect 11790 10996 11796 11008
rect 10888 10968 11796 10996
rect 10061 10959 10119 10965
rect 11790 10956 11796 10968
rect 11848 10956 11854 11008
rect 11882 10956 11888 11008
rect 11940 10996 11946 11008
rect 12452 10996 12480 11095
rect 12912 11064 12940 11095
rect 13078 11092 13084 11144
rect 13136 11092 13142 11144
rect 14461 11135 14519 11141
rect 14461 11101 14473 11135
rect 14507 11132 14519 11135
rect 14550 11132 14556 11144
rect 14507 11104 14556 11132
rect 14507 11101 14519 11104
rect 14461 11095 14519 11101
rect 14550 11092 14556 11104
rect 14608 11092 14614 11144
rect 14660 11141 14688 11172
rect 14918 11160 14924 11172
rect 14976 11160 14982 11212
rect 15028 11200 15056 11231
rect 15378 11200 15384 11212
rect 15028 11172 15384 11200
rect 15378 11160 15384 11172
rect 15436 11160 15442 11212
rect 15764 11200 15792 11308
rect 16574 11296 16580 11308
rect 16632 11296 16638 11348
rect 16758 11296 16764 11348
rect 16816 11336 16822 11348
rect 18233 11339 18291 11345
rect 18233 11336 18245 11339
rect 16816 11308 18245 11336
rect 16816 11296 16822 11308
rect 18233 11305 18245 11308
rect 18279 11336 18291 11339
rect 18322 11336 18328 11348
rect 18279 11308 18328 11336
rect 18279 11305 18291 11308
rect 18233 11299 18291 11305
rect 18322 11296 18328 11308
rect 18380 11296 18386 11348
rect 19242 11296 19248 11348
rect 19300 11336 19306 11348
rect 19429 11339 19487 11345
rect 19429 11336 19441 11339
rect 19300 11308 19441 11336
rect 19300 11296 19306 11308
rect 19429 11305 19441 11308
rect 19475 11305 19487 11339
rect 19429 11299 19487 11305
rect 19889 11339 19947 11345
rect 19889 11305 19901 11339
rect 19935 11336 19947 11339
rect 20165 11339 20223 11345
rect 20165 11336 20177 11339
rect 19935 11308 20177 11336
rect 19935 11305 19947 11308
rect 19889 11299 19947 11305
rect 20165 11305 20177 11308
rect 20211 11305 20223 11339
rect 20165 11299 20223 11305
rect 20254 11296 20260 11348
rect 20312 11336 20318 11348
rect 20312 11308 20944 11336
rect 20312 11296 20318 11308
rect 18046 11228 18052 11280
rect 18104 11268 18110 11280
rect 18104 11240 20392 11268
rect 18104 11228 18110 11240
rect 15672 11172 15792 11200
rect 16117 11203 16175 11209
rect 14645 11135 14703 11141
rect 14645 11101 14657 11135
rect 14691 11101 14703 11135
rect 14645 11095 14703 11101
rect 14734 11092 14740 11144
rect 14792 11092 14798 11144
rect 14829 11135 14887 11141
rect 14829 11101 14841 11135
rect 14875 11101 14887 11135
rect 14829 11095 14887 11101
rect 13170 11064 13176 11076
rect 12912 11036 13176 11064
rect 13170 11024 13176 11036
rect 13228 11024 13234 11076
rect 14844 11064 14872 11095
rect 15286 11092 15292 11144
rect 15344 11092 15350 11144
rect 15562 11132 15568 11144
rect 15396 11104 15568 11132
rect 15396 11073 15424 11104
rect 15562 11092 15568 11104
rect 15620 11092 15626 11144
rect 15672 11141 15700 11172
rect 16117 11169 16129 11203
rect 16163 11200 16175 11203
rect 16850 11200 16856 11212
rect 16163 11172 16856 11200
rect 16163 11169 16175 11172
rect 16117 11163 16175 11169
rect 16850 11160 16856 11172
rect 16908 11160 16914 11212
rect 19058 11160 19064 11212
rect 19116 11200 19122 11212
rect 20364 11209 20392 11240
rect 19705 11203 19763 11209
rect 19705 11200 19717 11203
rect 19116 11172 19717 11200
rect 19116 11160 19122 11172
rect 19705 11169 19717 11172
rect 19751 11169 19763 11203
rect 19705 11163 19763 11169
rect 20349 11203 20407 11209
rect 20349 11169 20361 11203
rect 20395 11169 20407 11203
rect 20349 11163 20407 11169
rect 20916 11200 20944 11308
rect 22572 11308 23336 11336
rect 22002 11200 22008 11212
rect 20916 11172 22008 11200
rect 15657 11135 15715 11141
rect 15657 11101 15669 11135
rect 15703 11101 15715 11135
rect 15657 11095 15715 11101
rect 15749 11135 15807 11141
rect 15749 11101 15761 11135
rect 15795 11101 15807 11135
rect 15749 11095 15807 11101
rect 15381 11067 15439 11073
rect 14844 11036 15332 11064
rect 11940 10968 12480 10996
rect 11940 10956 11946 10968
rect 12526 10956 12532 11008
rect 12584 10996 12590 11008
rect 12713 10999 12771 11005
rect 12713 10996 12725 10999
rect 12584 10968 12725 10996
rect 12584 10956 12590 10968
rect 12713 10965 12725 10968
rect 12759 10965 12771 10999
rect 12713 10959 12771 10965
rect 13262 10956 13268 11008
rect 13320 10996 13326 11008
rect 15010 10996 15016 11008
rect 13320 10968 15016 10996
rect 13320 10956 13326 10968
rect 15010 10956 15016 10968
rect 15068 10956 15074 11008
rect 15304 10996 15332 11036
rect 15381 11033 15393 11067
rect 15427 11033 15439 11067
rect 15381 11027 15439 11033
rect 15470 11024 15476 11076
rect 15528 11024 15534 11076
rect 15764 10996 15792 11095
rect 16022 11092 16028 11144
rect 16080 11092 16086 11144
rect 18046 11092 18052 11144
rect 18104 11092 18110 11144
rect 18690 11092 18696 11144
rect 18748 11132 18754 11144
rect 20916 11141 20944 11172
rect 22002 11160 22008 11172
rect 22060 11160 22066 11212
rect 19981 11135 20039 11141
rect 19981 11132 19993 11135
rect 18748 11104 19993 11132
rect 18748 11092 18754 11104
rect 19981 11101 19993 11104
rect 20027 11101 20039 11135
rect 19981 11095 20039 11101
rect 20441 11135 20499 11141
rect 20441 11101 20453 11135
rect 20487 11101 20499 11135
rect 20441 11095 20499 11101
rect 20901 11135 20959 11141
rect 20901 11101 20913 11135
rect 20947 11101 20959 11135
rect 20901 11095 20959 11101
rect 16298 11024 16304 11076
rect 16356 11064 16362 11076
rect 16393 11067 16451 11073
rect 16393 11064 16405 11067
rect 16356 11036 16405 11064
rect 16356 11024 16362 11036
rect 16393 11033 16405 11036
rect 16439 11033 16451 11067
rect 16393 11027 16451 11033
rect 16850 11024 16856 11076
rect 16908 11024 16914 11076
rect 20456 11064 20484 11095
rect 20990 11092 20996 11144
rect 21048 11132 21054 11144
rect 21085 11135 21143 11141
rect 21085 11132 21097 11135
rect 21048 11104 21097 11132
rect 21048 11092 21054 11104
rect 21085 11101 21097 11104
rect 21131 11101 21143 11135
rect 21085 11095 21143 11101
rect 21174 11092 21180 11144
rect 21232 11132 21238 11144
rect 21726 11132 21732 11144
rect 21232 11104 21732 11132
rect 21232 11092 21238 11104
rect 21726 11092 21732 11104
rect 21784 11132 21790 11144
rect 22572 11141 22600 11308
rect 22833 11271 22891 11277
rect 22833 11237 22845 11271
rect 22879 11268 22891 11271
rect 23014 11268 23020 11280
rect 22879 11240 23020 11268
rect 22879 11237 22891 11240
rect 22833 11231 22891 11237
rect 23014 11228 23020 11240
rect 23072 11228 23078 11280
rect 23106 11228 23112 11280
rect 23164 11268 23170 11280
rect 23308 11277 23336 11308
rect 23474 11296 23480 11348
rect 23532 11336 23538 11348
rect 23569 11339 23627 11345
rect 23569 11336 23581 11339
rect 23532 11308 23581 11336
rect 23532 11296 23538 11308
rect 23569 11305 23581 11308
rect 23615 11336 23627 11339
rect 23658 11336 23664 11348
rect 23615 11308 23664 11336
rect 23615 11305 23627 11308
rect 23569 11299 23627 11305
rect 23658 11296 23664 11308
rect 23716 11296 23722 11348
rect 23201 11271 23259 11277
rect 23201 11268 23213 11271
rect 23164 11240 23213 11268
rect 23164 11228 23170 11240
rect 23201 11237 23213 11240
rect 23247 11237 23259 11271
rect 23201 11231 23259 11237
rect 23293 11271 23351 11277
rect 23293 11237 23305 11271
rect 23339 11268 23351 11271
rect 24486 11268 24492 11280
rect 23339 11240 24492 11268
rect 23339 11237 23351 11240
rect 23293 11231 23351 11237
rect 24486 11228 24492 11240
rect 24544 11228 24550 11280
rect 23934 11200 23940 11212
rect 23308 11172 23940 11200
rect 22557 11135 22615 11141
rect 22557 11132 22569 11135
rect 21784 11104 22569 11132
rect 21784 11092 21790 11104
rect 22557 11101 22569 11104
rect 22603 11101 22615 11135
rect 22557 11095 22615 11101
rect 22925 11135 22983 11141
rect 22925 11101 22937 11135
rect 22971 11101 22983 11135
rect 22925 11095 22983 11101
rect 21450 11064 21456 11076
rect 20456 11036 21456 11064
rect 21450 11024 21456 11036
rect 21508 11024 21514 11076
rect 22186 11024 22192 11076
rect 22244 11064 22250 11076
rect 22833 11067 22891 11073
rect 22833 11064 22845 11067
rect 22244 11036 22845 11064
rect 22244 11024 22250 11036
rect 22833 11033 22845 11036
rect 22879 11033 22891 11067
rect 22940 11064 22968 11095
rect 23014 11092 23020 11144
rect 23072 11126 23078 11144
rect 23110 11135 23168 11141
rect 23110 11126 23122 11135
rect 23072 11101 23122 11126
rect 23156 11101 23168 11135
rect 23072 11098 23168 11101
rect 23072 11092 23078 11098
rect 23110 11095 23168 11098
rect 23308 11064 23336 11172
rect 23934 11160 23940 11172
rect 23992 11160 23998 11212
rect 24026 11160 24032 11212
rect 24084 11200 24090 11212
rect 24581 11203 24639 11209
rect 24581 11200 24593 11203
rect 24084 11172 24593 11200
rect 24084 11160 24090 11172
rect 24581 11169 24593 11172
rect 24627 11169 24639 11203
rect 24581 11163 24639 11169
rect 23385 11135 23443 11141
rect 23385 11101 23397 11135
rect 23431 11101 23443 11135
rect 23385 11095 23443 11101
rect 22940 11036 23336 11064
rect 23400 11064 23428 11095
rect 23750 11064 23756 11076
rect 23400 11036 23756 11064
rect 22833 11027 22891 11033
rect 23750 11024 23756 11036
rect 23808 11024 23814 11076
rect 23842 11024 23848 11076
rect 23900 11024 23906 11076
rect 23934 11024 23940 11076
rect 23992 11064 23998 11076
rect 24029 11067 24087 11073
rect 24029 11064 24041 11067
rect 23992 11036 24041 11064
rect 23992 11024 23998 11036
rect 24029 11033 24041 11036
rect 24075 11033 24087 11067
rect 24029 11027 24087 11033
rect 24857 11067 24915 11073
rect 24857 11033 24869 11067
rect 24903 11064 24915 11067
rect 25222 11064 25228 11076
rect 24903 11036 25228 11064
rect 24903 11033 24915 11036
rect 24857 11027 24915 11033
rect 15933 10999 15991 11005
rect 15933 10996 15945 10999
rect 15304 10968 15945 10996
rect 15933 10965 15945 10968
rect 15979 10996 15991 10999
rect 16114 10996 16120 11008
rect 15979 10968 16120 10996
rect 15979 10965 15991 10968
rect 15933 10959 15991 10965
rect 16114 10956 16120 10968
rect 16172 10956 16178 11008
rect 17865 10999 17923 11005
rect 17865 10965 17877 10999
rect 17911 10996 17923 10999
rect 18414 10996 18420 11008
rect 17911 10968 18420 10996
rect 17911 10965 17923 10968
rect 17865 10959 17923 10965
rect 18414 10956 18420 10968
rect 18472 10956 18478 11008
rect 20714 10956 20720 11008
rect 20772 10956 20778 11008
rect 22462 10956 22468 11008
rect 22520 10996 22526 11008
rect 22649 10999 22707 11005
rect 22649 10996 22661 10999
rect 22520 10968 22661 10996
rect 22520 10956 22526 10968
rect 22649 10965 22661 10968
rect 22695 10965 22707 10999
rect 22649 10959 22707 10965
rect 23014 10956 23020 11008
rect 23072 10996 23078 11008
rect 23290 10996 23296 11008
rect 23072 10968 23296 10996
rect 23072 10956 23078 10968
rect 23290 10956 23296 10968
rect 23348 10996 23354 11008
rect 23661 10999 23719 11005
rect 23661 10996 23673 10999
rect 23348 10968 23673 10996
rect 23348 10956 23354 10968
rect 23661 10965 23673 10968
rect 23707 10965 23719 10999
rect 24044 10996 24072 11027
rect 25222 11024 25228 11036
rect 25280 11024 25286 11076
rect 25314 10996 25320 11008
rect 24044 10968 25320 10996
rect 23661 10959 23719 10965
rect 25314 10956 25320 10968
rect 25372 10956 25378 11008
rect 1104 10906 28152 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 28152 10906
rect 1104 10832 28152 10854
rect 2314 10752 2320 10804
rect 2372 10792 2378 10804
rect 2409 10795 2467 10801
rect 2409 10792 2421 10795
rect 2372 10764 2421 10792
rect 2372 10752 2378 10764
rect 2409 10761 2421 10764
rect 2455 10761 2467 10795
rect 2682 10792 2688 10804
rect 2409 10755 2467 10761
rect 2516 10764 2688 10792
rect 1946 10724 1952 10736
rect 1872 10696 1952 10724
rect 1872 10665 1900 10696
rect 1946 10684 1952 10696
rect 2004 10684 2010 10736
rect 2516 10724 2544 10764
rect 2682 10752 2688 10764
rect 2740 10792 2746 10804
rect 2774 10792 2780 10804
rect 2740 10764 2780 10792
rect 2740 10752 2746 10764
rect 2774 10752 2780 10764
rect 2832 10752 2838 10804
rect 6546 10752 6552 10804
rect 6604 10792 6610 10804
rect 6733 10795 6791 10801
rect 6733 10792 6745 10795
rect 6604 10764 6745 10792
rect 6604 10752 6610 10764
rect 6733 10761 6745 10764
rect 6779 10761 6791 10795
rect 6733 10755 6791 10761
rect 8110 10752 8116 10804
rect 8168 10792 8174 10804
rect 8168 10764 9168 10792
rect 8168 10752 8174 10764
rect 2148 10696 2544 10724
rect 2792 10724 2820 10752
rect 2792 10696 3740 10724
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10625 1915 10659
rect 1857 10619 1915 10625
rect 1949 10591 2007 10597
rect 1949 10557 1961 10591
rect 1995 10588 2007 10591
rect 2148 10588 2176 10696
rect 2317 10659 2375 10665
rect 2317 10656 2329 10659
rect 1995 10560 2176 10588
rect 2240 10628 2329 10656
rect 1995 10557 2007 10560
rect 1949 10551 2007 10557
rect 2130 10412 2136 10464
rect 2188 10452 2194 10464
rect 2240 10461 2268 10628
rect 2317 10625 2329 10628
rect 2363 10625 2375 10659
rect 2317 10619 2375 10625
rect 2501 10659 2559 10665
rect 2501 10625 2513 10659
rect 2547 10656 2559 10659
rect 2590 10656 2596 10668
rect 2547 10628 2596 10656
rect 2547 10625 2559 10628
rect 2501 10619 2559 10625
rect 2590 10616 2596 10628
rect 2648 10616 2654 10668
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10625 3111 10659
rect 3053 10619 3111 10625
rect 2958 10548 2964 10600
rect 3016 10548 3022 10600
rect 3068 10588 3096 10619
rect 3326 10616 3332 10668
rect 3384 10656 3390 10668
rect 3712 10665 3740 10696
rect 7650 10684 7656 10736
rect 7708 10724 7714 10736
rect 9140 10733 9168 10764
rect 10870 10752 10876 10804
rect 10928 10792 10934 10804
rect 11241 10795 11299 10801
rect 11241 10792 11253 10795
rect 10928 10764 11253 10792
rect 10928 10752 10934 10764
rect 11241 10761 11253 10764
rect 11287 10792 11299 10795
rect 12158 10792 12164 10804
rect 11287 10764 12164 10792
rect 11287 10761 11299 10764
rect 11241 10755 11299 10761
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 12342 10792 12348 10804
rect 12268 10764 12348 10792
rect 7745 10727 7803 10733
rect 7745 10724 7757 10727
rect 7708 10696 7757 10724
rect 7708 10684 7714 10696
rect 7745 10693 7757 10696
rect 7791 10693 7803 10727
rect 7745 10687 7803 10693
rect 7929 10727 7987 10733
rect 7929 10693 7941 10727
rect 7975 10724 7987 10727
rect 9125 10727 9183 10733
rect 7975 10696 8708 10724
rect 7975 10693 7987 10696
rect 7929 10687 7987 10693
rect 3513 10659 3571 10665
rect 3513 10656 3525 10659
rect 3384 10628 3525 10656
rect 3384 10616 3390 10628
rect 3513 10625 3525 10628
rect 3559 10625 3571 10659
rect 3513 10619 3571 10625
rect 3697 10659 3755 10665
rect 3697 10625 3709 10659
rect 3743 10625 3755 10659
rect 3697 10619 3755 10625
rect 5626 10616 5632 10668
rect 5684 10656 5690 10668
rect 6365 10659 6423 10665
rect 6365 10656 6377 10659
rect 5684 10628 6377 10656
rect 5684 10616 5690 10628
rect 6365 10625 6377 10628
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 6458 10659 6516 10665
rect 6458 10625 6470 10659
rect 6504 10625 6516 10659
rect 6458 10619 6516 10625
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10656 7067 10659
rect 7374 10656 7380 10668
rect 7055 10628 7380 10656
rect 7055 10625 7067 10628
rect 7009 10619 7067 10625
rect 3605 10591 3663 10597
rect 3605 10588 3617 10591
rect 3068 10560 3617 10588
rect 3605 10557 3617 10560
rect 3651 10557 3663 10591
rect 3605 10551 3663 10557
rect 5534 10548 5540 10600
rect 5592 10588 5598 10600
rect 6472 10588 6500 10619
rect 7374 10616 7380 10628
rect 7432 10656 7438 10668
rect 7561 10659 7619 10665
rect 7561 10656 7573 10659
rect 7432 10628 7573 10656
rect 7432 10616 7438 10628
rect 7561 10625 7573 10628
rect 7607 10625 7619 10659
rect 7561 10619 7619 10625
rect 8386 10616 8392 10668
rect 8444 10616 8450 10668
rect 8680 10665 8708 10696
rect 9125 10693 9137 10727
rect 9171 10693 9183 10727
rect 12268 10724 12296 10764
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 12434 10752 12440 10804
rect 12492 10792 12498 10804
rect 12894 10792 12900 10804
rect 12952 10801 12958 10804
rect 12952 10795 12976 10801
rect 12492 10764 12900 10792
rect 12492 10752 12498 10764
rect 12894 10752 12900 10764
rect 12964 10761 12976 10795
rect 12952 10755 12976 10761
rect 12952 10752 12958 10755
rect 13998 10752 14004 10804
rect 14056 10792 14062 10804
rect 14277 10795 14335 10801
rect 14056 10764 14228 10792
rect 14056 10752 14062 10764
rect 9125 10687 9183 10693
rect 12100 10696 12296 10724
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 8846 10616 8852 10668
rect 8904 10616 8910 10668
rect 8941 10659 8999 10665
rect 8941 10625 8953 10659
rect 8987 10656 8999 10659
rect 8987 10628 9260 10656
rect 8987 10625 8999 10628
rect 8941 10619 8999 10625
rect 5592 10560 6500 10588
rect 6917 10591 6975 10597
rect 5592 10548 5598 10560
rect 6917 10557 6929 10591
rect 6963 10588 6975 10591
rect 7190 10588 7196 10600
rect 6963 10560 7196 10588
rect 6963 10557 6975 10560
rect 6917 10551 6975 10557
rect 3421 10523 3479 10529
rect 3421 10489 3433 10523
rect 3467 10520 3479 10523
rect 3970 10520 3976 10532
rect 3467 10492 3976 10520
rect 3467 10489 3479 10492
rect 3421 10483 3479 10489
rect 3970 10480 3976 10492
rect 4028 10480 4034 10532
rect 5997 10523 6055 10529
rect 5997 10489 6009 10523
rect 6043 10520 6055 10523
rect 6932 10520 6960 10551
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 8021 10591 8079 10597
rect 8021 10588 8033 10591
rect 7392 10560 8033 10588
rect 7392 10529 7420 10560
rect 8021 10557 8033 10560
rect 8067 10588 8079 10591
rect 8294 10588 8300 10600
rect 8067 10560 8300 10588
rect 8067 10557 8079 10560
rect 8021 10551 8079 10557
rect 8294 10548 8300 10560
rect 8352 10548 8358 10600
rect 8573 10591 8631 10597
rect 8573 10557 8585 10591
rect 8619 10588 8631 10591
rect 9122 10588 9128 10600
rect 8619 10560 9128 10588
rect 8619 10557 8631 10560
rect 8573 10551 8631 10557
rect 9122 10548 9128 10560
rect 9180 10548 9186 10600
rect 9232 10588 9260 10628
rect 9306 10616 9312 10668
rect 9364 10616 9370 10668
rect 11054 10616 11060 10668
rect 11112 10656 11118 10668
rect 11149 10659 11207 10665
rect 11149 10656 11161 10659
rect 11112 10628 11161 10656
rect 11112 10616 11118 10628
rect 11149 10625 11161 10628
rect 11195 10625 11207 10659
rect 11149 10619 11207 10625
rect 11333 10659 11391 10665
rect 11333 10625 11345 10659
rect 11379 10656 11391 10659
rect 11422 10656 11428 10668
rect 11379 10628 11428 10656
rect 11379 10625 11391 10628
rect 11333 10619 11391 10625
rect 11422 10616 11428 10628
rect 11480 10616 11486 10668
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 10042 10588 10048 10600
rect 9232 10560 10048 10588
rect 10042 10548 10048 10560
rect 10100 10588 10106 10600
rect 11606 10588 11612 10600
rect 10100 10560 11612 10588
rect 10100 10548 10106 10560
rect 11606 10548 11612 10560
rect 11664 10548 11670 10600
rect 6043 10492 6960 10520
rect 7377 10523 7435 10529
rect 6043 10489 6055 10492
rect 5997 10483 6055 10489
rect 7377 10489 7389 10523
rect 7423 10489 7435 10523
rect 7377 10483 7435 10489
rect 8757 10523 8815 10529
rect 8757 10489 8769 10523
rect 8803 10520 8815 10523
rect 11330 10520 11336 10532
rect 8803 10492 11336 10520
rect 8803 10489 8815 10492
rect 8757 10483 8815 10489
rect 11330 10480 11336 10492
rect 11388 10480 11394 10532
rect 11716 10520 11744 10619
rect 11882 10616 11888 10668
rect 11940 10616 11946 10668
rect 12100 10665 12128 10696
rect 12526 10684 12532 10736
rect 12584 10684 12590 10736
rect 12618 10684 12624 10736
rect 12676 10724 12682 10736
rect 12713 10727 12771 10733
rect 12713 10724 12725 10727
rect 12676 10696 12725 10724
rect 12676 10684 12682 10696
rect 12713 10693 12725 10696
rect 12759 10724 12771 10727
rect 14090 10724 14096 10736
rect 12759 10696 14096 10724
rect 12759 10693 12771 10696
rect 12713 10687 12771 10693
rect 14090 10684 14096 10696
rect 14148 10684 14154 10736
rect 14200 10724 14228 10764
rect 14277 10761 14289 10795
rect 14323 10792 14335 10795
rect 14918 10792 14924 10804
rect 14323 10764 14924 10792
rect 14323 10761 14335 10764
rect 14277 10755 14335 10761
rect 14918 10752 14924 10764
rect 14976 10752 14982 10804
rect 15102 10752 15108 10804
rect 15160 10752 15166 10804
rect 15286 10752 15292 10804
rect 15344 10792 15350 10804
rect 15657 10795 15715 10801
rect 15657 10792 15669 10795
rect 15344 10764 15669 10792
rect 15344 10752 15350 10764
rect 15657 10761 15669 10764
rect 15703 10792 15715 10795
rect 15930 10792 15936 10804
rect 15703 10764 15936 10792
rect 15703 10761 15715 10764
rect 15657 10755 15715 10761
rect 15930 10752 15936 10764
rect 15988 10752 15994 10804
rect 18509 10795 18567 10801
rect 18509 10761 18521 10795
rect 18555 10792 18567 10795
rect 18874 10792 18880 10804
rect 18555 10764 18880 10792
rect 18555 10761 18567 10764
rect 18509 10755 18567 10761
rect 18874 10752 18880 10764
rect 18932 10752 18938 10804
rect 20714 10792 20720 10804
rect 20364 10764 20720 10792
rect 14553 10727 14611 10733
rect 14200 10696 14504 10724
rect 12069 10659 12128 10665
rect 12069 10625 12081 10659
rect 12115 10628 12128 10659
rect 12115 10625 12127 10628
rect 12069 10619 12127 10625
rect 12250 10616 12256 10668
rect 12308 10616 12314 10668
rect 12544 10656 12572 10684
rect 12360 10628 12572 10656
rect 14185 10659 14243 10665
rect 11790 10548 11796 10600
rect 11848 10588 11854 10600
rect 11977 10591 12035 10597
rect 11977 10588 11989 10591
rect 11848 10560 11989 10588
rect 11848 10548 11854 10560
rect 11977 10557 11989 10560
rect 12023 10557 12035 10591
rect 12360 10588 12388 10628
rect 14185 10625 14197 10659
rect 14231 10656 14243 10659
rect 14366 10656 14372 10668
rect 14231 10628 14372 10656
rect 14231 10625 14243 10628
rect 14185 10619 14243 10625
rect 14366 10616 14372 10628
rect 14424 10616 14430 10668
rect 14476 10665 14504 10696
rect 14553 10693 14565 10727
rect 14599 10724 14611 10727
rect 14737 10727 14795 10733
rect 14737 10724 14749 10727
rect 14599 10696 14749 10724
rect 14599 10693 14611 10696
rect 14553 10687 14611 10693
rect 14737 10693 14749 10696
rect 14783 10693 14795 10727
rect 14737 10687 14795 10693
rect 14826 10684 14832 10736
rect 14884 10724 14890 10736
rect 15197 10727 15255 10733
rect 15197 10724 15209 10727
rect 14884 10696 15209 10724
rect 14884 10684 14890 10696
rect 15197 10693 15209 10696
rect 15243 10693 15255 10727
rect 15197 10687 15255 10693
rect 15378 10684 15384 10736
rect 15436 10724 15442 10736
rect 15562 10724 15568 10736
rect 15436 10696 15568 10724
rect 15436 10684 15442 10696
rect 15562 10684 15568 10696
rect 15620 10724 15626 10736
rect 15620 10696 15976 10724
rect 15620 10684 15626 10696
rect 14461 10659 14519 10665
rect 14461 10625 14473 10659
rect 14507 10625 14519 10659
rect 14645 10659 14703 10665
rect 14645 10658 14657 10659
rect 14461 10619 14519 10625
rect 14568 10630 14657 10658
rect 11977 10551 12035 10557
rect 12084 10560 12388 10588
rect 12084 10520 12112 10560
rect 12526 10548 12532 10600
rect 12584 10588 12590 10600
rect 12710 10588 12716 10600
rect 12584 10560 12716 10588
rect 12584 10548 12590 10560
rect 12710 10548 12716 10560
rect 12768 10548 12774 10600
rect 14568 10588 14596 10630
rect 14645 10625 14657 10630
rect 14691 10625 14703 10659
rect 14645 10619 14703 10625
rect 14918 10616 14924 10668
rect 14976 10616 14982 10668
rect 15010 10616 15016 10668
rect 15068 10656 15074 10668
rect 15473 10659 15531 10665
rect 15473 10656 15485 10659
rect 15068 10628 15485 10656
rect 15068 10616 15074 10628
rect 15473 10625 15485 10628
rect 15519 10625 15531 10659
rect 15473 10619 15531 10625
rect 15749 10659 15807 10665
rect 15749 10625 15761 10659
rect 15795 10656 15807 10659
rect 15838 10656 15844 10668
rect 15795 10628 15844 10656
rect 15795 10625 15807 10628
rect 15749 10619 15807 10625
rect 15838 10616 15844 10628
rect 15896 10616 15902 10668
rect 15948 10665 15976 10696
rect 16758 10684 16764 10736
rect 16816 10724 16822 10736
rect 17218 10724 17224 10736
rect 16816 10696 17224 10724
rect 16816 10684 16822 10696
rect 17218 10684 17224 10696
rect 17276 10684 17282 10736
rect 18417 10727 18475 10733
rect 18417 10693 18429 10727
rect 18463 10724 18475 10727
rect 19702 10724 19708 10736
rect 18463 10696 19708 10724
rect 18463 10693 18475 10696
rect 18417 10687 18475 10693
rect 19702 10684 19708 10696
rect 19760 10684 19766 10736
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10625 15991 10659
rect 15933 10619 15991 10625
rect 16114 10616 16120 10668
rect 16172 10616 16178 10668
rect 16301 10659 16359 10665
rect 16301 10625 16313 10659
rect 16347 10656 16359 10659
rect 17034 10656 17040 10668
rect 16347 10628 17040 10656
rect 16347 10625 16359 10628
rect 16301 10619 16359 10625
rect 17034 10616 17040 10628
rect 17092 10656 17098 10668
rect 18506 10656 18512 10668
rect 17092 10628 18512 10656
rect 17092 10616 17098 10628
rect 18506 10616 18512 10628
rect 18564 10616 18570 10668
rect 18969 10659 19027 10665
rect 18969 10625 18981 10659
rect 19015 10656 19027 10659
rect 19242 10656 19248 10668
rect 19015 10628 19248 10656
rect 19015 10625 19027 10628
rect 18969 10619 19027 10625
rect 19242 10616 19248 10628
rect 19300 10616 19306 10668
rect 19610 10616 19616 10668
rect 19668 10656 19674 10668
rect 19797 10659 19855 10665
rect 19797 10656 19809 10659
rect 19668 10628 19809 10656
rect 19668 10616 19674 10628
rect 19797 10625 19809 10628
rect 19843 10656 19855 10659
rect 20073 10659 20131 10665
rect 20073 10656 20085 10659
rect 19843 10628 20085 10656
rect 19843 10625 19855 10628
rect 19797 10619 19855 10625
rect 20073 10625 20085 10628
rect 20119 10625 20131 10659
rect 20073 10619 20131 10625
rect 20257 10659 20315 10665
rect 20257 10625 20269 10659
rect 20303 10656 20315 10659
rect 20364 10656 20392 10764
rect 20714 10752 20720 10764
rect 20772 10752 20778 10804
rect 23658 10792 23664 10804
rect 20916 10764 23336 10792
rect 20441 10727 20499 10733
rect 20441 10693 20453 10727
rect 20487 10724 20499 10727
rect 20625 10727 20683 10733
rect 20625 10724 20637 10727
rect 20487 10696 20637 10724
rect 20487 10693 20499 10696
rect 20441 10687 20499 10693
rect 20625 10693 20637 10696
rect 20671 10693 20683 10727
rect 20916 10724 20944 10764
rect 20625 10687 20683 10693
rect 20732 10696 20944 10724
rect 20303 10628 20392 10656
rect 20303 10625 20315 10628
rect 20257 10619 20315 10625
rect 20530 10616 20536 10668
rect 20588 10616 20594 10668
rect 13096 10560 14596 10588
rect 11716 10492 12112 10520
rect 12342 10480 12348 10532
rect 12400 10520 12406 10532
rect 12400 10492 12940 10520
rect 12400 10480 12406 10492
rect 2225 10455 2283 10461
rect 2225 10452 2237 10455
rect 2188 10424 2237 10452
rect 2188 10412 2194 10424
rect 2225 10421 2237 10424
rect 2271 10421 2283 10455
rect 2225 10415 2283 10421
rect 8202 10412 8208 10464
rect 8260 10452 8266 10464
rect 10594 10452 10600 10464
rect 8260 10424 10600 10452
rect 8260 10412 8266 10424
rect 10594 10412 10600 10424
rect 10652 10412 10658 10464
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10452 12495 10455
rect 12802 10452 12808 10464
rect 12483 10424 12808 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 12912 10461 12940 10492
rect 12986 10480 12992 10532
rect 13044 10520 13050 10532
rect 13096 10529 13124 10560
rect 15378 10548 15384 10600
rect 15436 10548 15442 10600
rect 16025 10591 16083 10597
rect 16025 10557 16037 10591
rect 16071 10557 16083 10591
rect 16025 10551 16083 10557
rect 13081 10523 13139 10529
rect 13081 10520 13093 10523
rect 13044 10492 13093 10520
rect 13044 10480 13050 10492
rect 13081 10489 13093 10492
rect 13127 10489 13139 10523
rect 13081 10483 13139 10489
rect 13906 10480 13912 10532
rect 13964 10520 13970 10532
rect 16040 10520 16068 10551
rect 18690 10548 18696 10600
rect 18748 10548 18754 10600
rect 18782 10548 18788 10600
rect 18840 10548 18846 10600
rect 18874 10548 18880 10600
rect 18932 10548 18938 10600
rect 19978 10588 19984 10600
rect 18984 10560 19984 10588
rect 16666 10520 16672 10532
rect 13964 10492 16068 10520
rect 16408 10492 16672 10520
rect 13964 10480 13970 10492
rect 12897 10455 12955 10461
rect 12897 10421 12909 10455
rect 12943 10421 12955 10455
rect 12897 10415 12955 10421
rect 15473 10455 15531 10461
rect 15473 10421 15485 10455
rect 15519 10452 15531 10455
rect 16408 10452 16436 10492
rect 16666 10480 16672 10492
rect 16724 10480 16730 10532
rect 17310 10480 17316 10532
rect 17368 10520 17374 10532
rect 18984 10520 19012 10560
rect 19978 10548 19984 10560
rect 20036 10548 20042 10600
rect 20162 10548 20168 10600
rect 20220 10588 20226 10600
rect 20732 10588 20760 10696
rect 20990 10684 20996 10736
rect 21048 10724 21054 10736
rect 21361 10727 21419 10733
rect 21361 10724 21373 10727
rect 21048 10696 21373 10724
rect 21048 10684 21054 10696
rect 21192 10665 21220 10696
rect 21361 10693 21373 10696
rect 21407 10693 21419 10727
rect 21361 10687 21419 10693
rect 22830 10684 22836 10736
rect 22888 10684 22894 10736
rect 23106 10733 23112 10736
rect 23049 10727 23112 10733
rect 23049 10693 23061 10727
rect 23095 10693 23112 10727
rect 23049 10687 23112 10693
rect 23106 10684 23112 10687
rect 23164 10724 23170 10736
rect 23308 10724 23336 10764
rect 23584 10764 23664 10792
rect 23474 10724 23480 10736
rect 23164 10696 23244 10724
rect 23164 10684 23170 10696
rect 20809 10659 20867 10665
rect 20809 10625 20821 10659
rect 20855 10625 20867 10659
rect 20809 10619 20867 10625
rect 20901 10659 20959 10665
rect 20901 10625 20913 10659
rect 20947 10625 20959 10659
rect 20901 10619 20959 10625
rect 21085 10659 21143 10665
rect 21085 10625 21097 10659
rect 21131 10625 21143 10659
rect 21085 10619 21143 10625
rect 21177 10659 21235 10665
rect 21177 10625 21189 10659
rect 21223 10625 21235 10659
rect 21177 10619 21235 10625
rect 20220 10560 20760 10588
rect 20220 10548 20226 10560
rect 17368 10492 19012 10520
rect 17368 10480 17374 10492
rect 19242 10480 19248 10532
rect 19300 10520 19306 10532
rect 20824 10520 20852 10619
rect 19300 10492 20852 10520
rect 19300 10480 19306 10492
rect 15519 10424 16436 10452
rect 16485 10455 16543 10461
rect 15519 10421 15531 10424
rect 15473 10415 15531 10421
rect 16485 10421 16497 10455
rect 16531 10452 16543 10455
rect 16850 10452 16856 10464
rect 16531 10424 16856 10452
rect 16531 10421 16543 10424
rect 16485 10415 16543 10421
rect 16850 10412 16856 10424
rect 16908 10412 16914 10464
rect 18046 10412 18052 10464
rect 18104 10452 18110 10464
rect 18966 10452 18972 10464
rect 18104 10424 18972 10452
rect 18104 10412 18110 10424
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 19886 10412 19892 10464
rect 19944 10412 19950 10464
rect 19978 10412 19984 10464
rect 20036 10452 20042 10464
rect 20916 10452 20944 10619
rect 21100 10588 21128 10619
rect 21450 10616 21456 10668
rect 21508 10616 21514 10668
rect 21266 10588 21272 10600
rect 21100 10560 21272 10588
rect 21266 10548 21272 10560
rect 21324 10548 21330 10600
rect 23216 10588 23244 10696
rect 23308 10696 23480 10724
rect 23308 10665 23336 10696
rect 23474 10684 23480 10696
rect 23532 10684 23538 10736
rect 23584 10733 23612 10764
rect 23658 10752 23664 10764
rect 23716 10752 23722 10804
rect 23842 10752 23848 10804
rect 23900 10792 23906 10804
rect 23900 10764 25176 10792
rect 23900 10752 23906 10764
rect 23569 10727 23627 10733
rect 23569 10693 23581 10727
rect 23615 10693 23627 10727
rect 23569 10687 23627 10693
rect 24026 10684 24032 10736
rect 24084 10684 24090 10736
rect 25148 10665 25176 10764
rect 23293 10659 23351 10665
rect 23293 10625 23305 10659
rect 23339 10625 23351 10659
rect 23293 10619 23351 10625
rect 25133 10659 25191 10665
rect 25133 10625 25145 10659
rect 25179 10625 25191 10659
rect 25133 10619 25191 10625
rect 25314 10616 25320 10668
rect 25372 10616 25378 10668
rect 25225 10591 25283 10597
rect 25225 10588 25237 10591
rect 23216 10560 25237 10588
rect 25225 10557 25237 10560
rect 25271 10557 25283 10591
rect 25225 10551 25283 10557
rect 24578 10480 24584 10532
rect 24636 10520 24642 10532
rect 24762 10520 24768 10532
rect 24636 10492 24768 10520
rect 24636 10480 24642 10492
rect 24762 10480 24768 10492
rect 24820 10520 24826 10532
rect 25041 10523 25099 10529
rect 25041 10520 25053 10523
rect 24820 10492 25053 10520
rect 24820 10480 24826 10492
rect 25041 10489 25053 10492
rect 25087 10489 25099 10523
rect 25041 10483 25099 10489
rect 20036 10424 20944 10452
rect 20036 10412 20042 10424
rect 23014 10412 23020 10464
rect 23072 10412 23078 10464
rect 23201 10455 23259 10461
rect 23201 10421 23213 10455
rect 23247 10452 23259 10455
rect 24670 10452 24676 10464
rect 23247 10424 24676 10452
rect 23247 10421 23259 10424
rect 23201 10415 23259 10421
rect 24670 10412 24676 10424
rect 24728 10412 24734 10464
rect 1104 10362 28152 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 28152 10362
rect 1104 10288 28152 10310
rect 7653 10251 7711 10257
rect 7653 10217 7665 10251
rect 7699 10248 7711 10251
rect 8110 10248 8116 10260
rect 7699 10220 8116 10248
rect 7699 10217 7711 10220
rect 7653 10211 7711 10217
rect 8110 10208 8116 10220
rect 8168 10248 8174 10260
rect 8846 10248 8852 10260
rect 8168 10220 8852 10248
rect 8168 10208 8174 10220
rect 8846 10208 8852 10220
rect 8904 10208 8910 10260
rect 9125 10251 9183 10257
rect 9125 10217 9137 10251
rect 9171 10217 9183 10251
rect 9125 10211 9183 10217
rect 8202 10140 8208 10192
rect 8260 10140 8266 10192
rect 8386 10140 8392 10192
rect 8444 10180 8450 10192
rect 9140 10180 9168 10211
rect 9306 10208 9312 10260
rect 9364 10208 9370 10260
rect 9950 10208 9956 10260
rect 10008 10208 10014 10260
rect 10137 10251 10195 10257
rect 10137 10217 10149 10251
rect 10183 10248 10195 10251
rect 10594 10248 10600 10260
rect 10183 10220 10600 10248
rect 10183 10217 10195 10220
rect 10137 10211 10195 10217
rect 10594 10208 10600 10220
rect 10652 10208 10658 10260
rect 13906 10208 13912 10260
rect 13964 10208 13970 10260
rect 13998 10208 14004 10260
rect 14056 10248 14062 10260
rect 14056 10220 14412 10248
rect 14056 10208 14062 10220
rect 8444 10152 9168 10180
rect 12713 10183 12771 10189
rect 8444 10140 8450 10152
rect 12713 10149 12725 10183
rect 12759 10180 12771 10183
rect 12894 10180 12900 10192
rect 12759 10152 12900 10180
rect 12759 10149 12771 10152
rect 12713 10143 12771 10149
rect 12894 10140 12900 10152
rect 12952 10140 12958 10192
rect 13078 10140 13084 10192
rect 13136 10180 13142 10192
rect 13136 10152 14320 10180
rect 13136 10140 13142 10152
rect 2130 10072 2136 10124
rect 2188 10072 2194 10124
rect 7926 10072 7932 10124
rect 7984 10112 7990 10124
rect 12250 10112 12256 10124
rect 7984 10084 12256 10112
rect 7984 10072 7990 10084
rect 2225 10047 2283 10053
rect 2225 10013 2237 10047
rect 2271 10044 2283 10047
rect 2590 10044 2596 10056
rect 2271 10016 2596 10044
rect 2271 10013 2283 10016
rect 2225 10007 2283 10013
rect 2590 10004 2596 10016
rect 2648 10004 2654 10056
rect 7374 10004 7380 10056
rect 7432 10044 7438 10056
rect 7561 10047 7619 10053
rect 7561 10044 7573 10047
rect 7432 10016 7573 10044
rect 7432 10004 7438 10016
rect 7561 10013 7573 10016
rect 7607 10013 7619 10047
rect 7561 10007 7619 10013
rect 7650 10004 7656 10056
rect 7708 10044 7714 10056
rect 8036 10053 8064 10084
rect 12250 10072 12256 10084
rect 12308 10072 12314 10124
rect 12802 10072 12808 10124
rect 12860 10112 12866 10124
rect 12860 10084 13492 10112
rect 12860 10072 12866 10084
rect 7745 10047 7803 10053
rect 7745 10044 7757 10047
rect 7708 10016 7757 10044
rect 7708 10004 7714 10016
rect 7745 10013 7757 10016
rect 7791 10044 7803 10047
rect 7837 10047 7895 10053
rect 7837 10044 7849 10047
rect 7791 10016 7849 10044
rect 7791 10013 7803 10016
rect 7745 10007 7803 10013
rect 7837 10013 7849 10016
rect 7883 10013 7895 10047
rect 7837 10007 7895 10013
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10013 8079 10047
rect 8481 10047 8539 10053
rect 8481 10044 8493 10047
rect 8021 10007 8079 10013
rect 8128 10016 8493 10044
rect 7466 9936 7472 9988
rect 7524 9976 7530 9988
rect 8128 9976 8156 10016
rect 8481 10013 8493 10016
rect 8527 10013 8539 10047
rect 8481 10007 8539 10013
rect 8757 10047 8815 10053
rect 8757 10013 8769 10047
rect 8803 10044 8815 10047
rect 9769 10047 9827 10053
rect 9769 10044 9781 10047
rect 8803 10016 9781 10044
rect 8803 10013 8815 10016
rect 8757 10007 8815 10013
rect 9769 10013 9781 10016
rect 9815 10013 9827 10047
rect 9769 10007 9827 10013
rect 10045 10047 10103 10053
rect 10045 10013 10057 10047
rect 10091 10044 10103 10047
rect 10134 10044 10140 10056
rect 10091 10016 10140 10044
rect 10091 10013 10103 10016
rect 10045 10007 10103 10013
rect 10134 10004 10140 10016
rect 10192 10004 10198 10056
rect 11146 10004 11152 10056
rect 11204 10004 11210 10056
rect 12434 10004 12440 10056
rect 12492 10004 12498 10056
rect 12897 10047 12955 10053
rect 12897 10044 12909 10047
rect 12728 10016 12909 10044
rect 7524 9948 8156 9976
rect 7524 9936 7530 9948
rect 8294 9936 8300 9988
rect 8352 9976 8358 9988
rect 8941 9979 8999 9985
rect 8941 9976 8953 9979
rect 8352 9948 8953 9976
rect 8352 9936 8358 9948
rect 8941 9945 8953 9948
rect 8987 9945 8999 9979
rect 8941 9939 8999 9945
rect 9122 9936 9128 9988
rect 9180 9985 9186 9988
rect 9180 9979 9199 9985
rect 9187 9945 9199 9979
rect 9180 9939 9199 9945
rect 9401 9979 9459 9985
rect 9401 9945 9413 9979
rect 9447 9976 9459 9979
rect 9447 9948 9812 9976
rect 9447 9945 9459 9948
rect 9401 9939 9459 9945
rect 9180 9936 9186 9939
rect 9784 9920 9812 9948
rect 11422 9936 11428 9988
rect 11480 9976 11486 9988
rect 11974 9976 11980 9988
rect 11480 9948 11980 9976
rect 11480 9936 11486 9948
rect 11974 9936 11980 9948
rect 12032 9976 12038 9988
rect 12342 9976 12348 9988
rect 12032 9948 12348 9976
rect 12032 9936 12038 9948
rect 12342 9936 12348 9948
rect 12400 9976 12406 9988
rect 12529 9979 12587 9985
rect 12529 9976 12541 9979
rect 12400 9948 12541 9976
rect 12400 9936 12406 9948
rect 12529 9945 12541 9948
rect 12575 9945 12587 9979
rect 12529 9939 12587 9945
rect 12618 9936 12624 9988
rect 12676 9976 12682 9988
rect 12728 9985 12756 10016
rect 12897 10013 12909 10016
rect 12943 10013 12955 10047
rect 12897 10007 12955 10013
rect 13078 10004 13084 10056
rect 13136 10004 13142 10056
rect 13464 10053 13492 10084
rect 13265 10047 13323 10053
rect 13265 10013 13277 10047
rect 13311 10013 13323 10047
rect 13265 10007 13323 10013
rect 13449 10047 13507 10053
rect 13449 10013 13461 10047
rect 13495 10013 13507 10047
rect 13449 10007 13507 10013
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10044 13783 10047
rect 13771 10016 14044 10044
rect 13771 10013 13783 10016
rect 13725 10007 13783 10013
rect 12713 9979 12771 9985
rect 12713 9976 12725 9979
rect 12676 9948 12725 9976
rect 12676 9936 12682 9948
rect 12713 9945 12725 9948
rect 12759 9945 12771 9979
rect 13280 9976 13308 10007
rect 12713 9939 12771 9945
rect 13004 9948 13308 9976
rect 2593 9911 2651 9917
rect 2593 9877 2605 9911
rect 2639 9908 2651 9911
rect 2958 9908 2964 9920
rect 2639 9880 2964 9908
rect 2639 9877 2651 9880
rect 2593 9871 2651 9877
rect 2958 9868 2964 9880
rect 3016 9868 3022 9920
rect 7929 9911 7987 9917
rect 7929 9877 7941 9911
rect 7975 9908 7987 9911
rect 8389 9911 8447 9917
rect 8389 9908 8401 9911
rect 7975 9880 8401 9908
rect 7975 9877 7987 9880
rect 7929 9871 7987 9877
rect 8389 9877 8401 9880
rect 8435 9877 8447 9911
rect 8389 9871 8447 9877
rect 8573 9911 8631 9917
rect 8573 9877 8585 9911
rect 8619 9908 8631 9911
rect 8754 9908 8760 9920
rect 8619 9880 8760 9908
rect 8619 9877 8631 9880
rect 8573 9871 8631 9877
rect 8754 9868 8760 9880
rect 8812 9868 8818 9920
rect 9582 9868 9588 9920
rect 9640 9868 9646 9920
rect 9674 9868 9680 9920
rect 9732 9868 9738 9920
rect 9766 9868 9772 9920
rect 9824 9868 9830 9920
rect 11054 9868 11060 9920
rect 11112 9868 11118 9920
rect 12802 9868 12808 9920
rect 12860 9908 12866 9920
rect 13004 9917 13032 9948
rect 12989 9911 13047 9917
rect 12989 9908 13001 9911
rect 12860 9880 13001 9908
rect 12860 9868 12866 9880
rect 12989 9877 13001 9880
rect 13035 9877 13047 9911
rect 14016 9908 14044 10016
rect 14090 10004 14096 10056
rect 14148 10004 14154 10056
rect 14292 10053 14320 10152
rect 14384 10112 14412 10220
rect 14826 10208 14832 10260
rect 14884 10208 14890 10260
rect 15286 10257 15292 10260
rect 15280 10248 15292 10257
rect 15199 10220 15292 10248
rect 15280 10211 15292 10220
rect 15344 10248 15350 10260
rect 15746 10248 15752 10260
rect 15344 10220 15752 10248
rect 15286 10208 15292 10211
rect 15344 10208 15350 10220
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 16025 10251 16083 10257
rect 16025 10217 16037 10251
rect 16071 10248 16083 10251
rect 16206 10248 16212 10260
rect 16071 10220 16212 10248
rect 16071 10217 16083 10220
rect 16025 10211 16083 10217
rect 16206 10208 16212 10220
rect 16264 10208 16270 10260
rect 17129 10251 17187 10257
rect 17129 10217 17141 10251
rect 17175 10248 17187 10251
rect 18138 10248 18144 10260
rect 17175 10220 18144 10248
rect 17175 10217 17187 10220
rect 17129 10211 17187 10217
rect 18138 10208 18144 10220
rect 18196 10208 18202 10260
rect 18325 10251 18383 10257
rect 18325 10217 18337 10251
rect 18371 10248 18383 10251
rect 18782 10248 18788 10260
rect 18371 10220 18788 10248
rect 18371 10217 18383 10220
rect 18325 10211 18383 10217
rect 18782 10208 18788 10220
rect 18840 10208 18846 10260
rect 20990 10208 20996 10260
rect 21048 10248 21054 10260
rect 21450 10248 21456 10260
rect 21048 10220 21456 10248
rect 21048 10208 21054 10220
rect 21450 10208 21456 10220
rect 21508 10248 21514 10260
rect 21913 10251 21971 10257
rect 21913 10248 21925 10251
rect 21508 10220 21925 10248
rect 21508 10208 21514 10220
rect 21913 10217 21925 10220
rect 21959 10217 21971 10251
rect 21913 10211 21971 10217
rect 22554 10208 22560 10260
rect 22612 10248 22618 10260
rect 23293 10251 23351 10257
rect 23293 10248 23305 10251
rect 22612 10220 23305 10248
rect 22612 10208 22618 10220
rect 23293 10217 23305 10220
rect 23339 10217 23351 10251
rect 23293 10211 23351 10217
rect 23658 10208 23664 10260
rect 23716 10248 23722 10260
rect 23753 10251 23811 10257
rect 23753 10248 23765 10251
rect 23716 10220 23765 10248
rect 23716 10208 23722 10220
rect 23753 10217 23765 10220
rect 23799 10248 23811 10251
rect 23934 10248 23940 10260
rect 23799 10220 23940 10248
rect 23799 10217 23811 10220
rect 23753 10211 23811 10217
rect 23934 10208 23940 10220
rect 23992 10208 23998 10260
rect 15473 10183 15531 10189
rect 15473 10149 15485 10183
rect 15519 10149 15531 10183
rect 18598 10180 18604 10192
rect 15473 10143 15531 10149
rect 16408 10152 18604 10180
rect 15286 10112 15292 10124
rect 14384 10084 15292 10112
rect 14384 10053 14412 10084
rect 15286 10072 15292 10084
rect 15344 10072 15350 10124
rect 14277 10047 14335 10053
rect 14277 10013 14289 10047
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 14369 10047 14427 10053
rect 14369 10013 14381 10047
rect 14415 10013 14427 10047
rect 14369 10007 14427 10013
rect 14458 10004 14464 10056
rect 14516 10004 14522 10056
rect 14829 10047 14887 10053
rect 14829 10013 14841 10047
rect 14875 10044 14887 10047
rect 14918 10044 14924 10056
rect 14875 10016 14924 10044
rect 14875 10013 14887 10016
rect 14829 10007 14887 10013
rect 14918 10004 14924 10016
rect 14976 10004 14982 10056
rect 15013 10047 15071 10053
rect 15013 10013 15025 10047
rect 15059 10044 15071 10047
rect 15059 10016 15148 10044
rect 15059 10013 15071 10016
rect 15013 10007 15071 10013
rect 15120 9985 15148 10016
rect 15378 10004 15384 10056
rect 15436 10044 15442 10056
rect 15488 10044 15516 10143
rect 15436 10016 15516 10044
rect 16117 10047 16175 10053
rect 15436 10004 15442 10016
rect 16117 10013 16129 10047
rect 16163 10044 16175 10047
rect 16408 10044 16436 10152
rect 18598 10140 18604 10152
rect 18656 10140 18662 10192
rect 19886 10140 19892 10192
rect 19944 10180 19950 10192
rect 19944 10152 20300 10180
rect 19944 10140 19950 10152
rect 16850 10072 16856 10124
rect 16908 10112 16914 10124
rect 16908 10084 18184 10112
rect 16908 10072 16914 10084
rect 16163 10016 16436 10044
rect 16163 10013 16175 10016
rect 16117 10007 16175 10013
rect 16482 10004 16488 10056
rect 16540 10004 16546 10056
rect 16633 10047 16691 10053
rect 16633 10013 16645 10047
rect 16679 10044 16691 10047
rect 16679 10013 16712 10044
rect 16633 10007 16712 10013
rect 15105 9979 15163 9985
rect 15105 9945 15117 9979
rect 15151 9976 15163 9979
rect 16684 9976 16712 10007
rect 16942 10004 16948 10056
rect 17000 10053 17006 10056
rect 17000 10044 17008 10053
rect 17221 10047 17279 10053
rect 17000 10016 17045 10044
rect 17000 10007 17008 10016
rect 17221 10013 17233 10047
rect 17267 10044 17279 10047
rect 17310 10044 17316 10056
rect 17267 10016 17316 10044
rect 17267 10013 17279 10016
rect 17221 10007 17279 10013
rect 17000 10004 17006 10007
rect 17310 10004 17316 10016
rect 17368 10044 17374 10056
rect 17678 10044 17684 10056
rect 17368 10016 17684 10044
rect 17368 10004 17374 10016
rect 17678 10004 17684 10016
rect 17736 10004 17742 10056
rect 17954 10004 17960 10056
rect 18012 10004 18018 10056
rect 18156 10053 18184 10084
rect 18506 10072 18512 10124
rect 18564 10072 18570 10124
rect 20162 10072 20168 10124
rect 20220 10072 20226 10124
rect 20272 10112 20300 10152
rect 22462 10140 22468 10192
rect 22520 10180 22526 10192
rect 22520 10152 23520 10180
rect 22520 10140 22526 10152
rect 20441 10115 20499 10121
rect 20441 10112 20453 10115
rect 20272 10084 20453 10112
rect 20441 10081 20453 10084
rect 20487 10081 20499 10115
rect 20441 10075 20499 10081
rect 21634 10072 21640 10124
rect 21692 10112 21698 10124
rect 23385 10115 23443 10121
rect 23385 10112 23397 10115
rect 21692 10084 23397 10112
rect 21692 10072 21698 10084
rect 23385 10081 23397 10084
rect 23431 10081 23443 10115
rect 23385 10075 23443 10081
rect 18141 10047 18199 10053
rect 18141 10013 18153 10047
rect 18187 10013 18199 10047
rect 18141 10007 18199 10013
rect 18414 10004 18420 10056
rect 18472 10004 18478 10056
rect 22738 10004 22744 10056
rect 22796 10044 22802 10056
rect 23293 10047 23351 10053
rect 23293 10044 23305 10047
rect 22796 10016 23305 10044
rect 22796 10004 22802 10016
rect 23293 10013 23305 10016
rect 23339 10013 23351 10047
rect 23492 10044 23520 10152
rect 23566 10140 23572 10192
rect 23624 10180 23630 10192
rect 23624 10152 24440 10180
rect 23624 10140 23630 10152
rect 24412 10124 24440 10152
rect 23750 10072 23756 10124
rect 23808 10112 23814 10124
rect 24302 10112 24308 10124
rect 23808 10084 24308 10112
rect 23808 10072 23814 10084
rect 24044 10053 24072 10084
rect 24302 10072 24308 10084
rect 24360 10072 24366 10124
rect 24394 10072 24400 10124
rect 24452 10072 24458 10124
rect 24670 10072 24676 10124
rect 24728 10072 24734 10124
rect 23569 10047 23627 10053
rect 23569 10044 23581 10047
rect 23492 10016 23581 10044
rect 23293 10007 23351 10013
rect 23569 10013 23581 10016
rect 23615 10044 23627 10047
rect 23937 10047 23995 10053
rect 23937 10044 23949 10047
rect 23615 10016 23949 10044
rect 23615 10013 23627 10016
rect 23569 10007 23627 10013
rect 23937 10013 23949 10016
rect 23983 10013 23995 10047
rect 23937 10007 23995 10013
rect 24029 10047 24087 10053
rect 24029 10013 24041 10047
rect 24075 10013 24087 10047
rect 24029 10007 24087 10013
rect 15151 9948 16712 9976
rect 15151 9945 15163 9948
rect 15105 9939 15163 9945
rect 14645 9911 14703 9917
rect 14645 9908 14657 9911
rect 14016 9880 14657 9908
rect 12989 9871 13047 9877
rect 14645 9877 14657 9880
rect 14691 9908 14703 9911
rect 15010 9908 15016 9920
rect 14691 9880 15016 9908
rect 14691 9877 14703 9880
rect 14645 9871 14703 9877
rect 15010 9868 15016 9880
rect 15068 9868 15074 9920
rect 15194 9868 15200 9920
rect 15252 9908 15258 9920
rect 15305 9911 15363 9917
rect 15305 9908 15317 9911
rect 15252 9880 15317 9908
rect 15252 9868 15258 9880
rect 15305 9877 15317 9880
rect 15351 9877 15363 9911
rect 16684 9908 16712 9948
rect 16758 9936 16764 9988
rect 16816 9936 16822 9988
rect 16850 9936 16856 9988
rect 16908 9936 16914 9988
rect 17589 9979 17647 9985
rect 17589 9945 17601 9979
rect 17635 9976 17647 9979
rect 18046 9976 18052 9988
rect 17635 9948 18052 9976
rect 17635 9945 17647 9948
rect 17589 9939 17647 9945
rect 18046 9936 18052 9948
rect 18104 9936 18110 9988
rect 17126 9908 17132 9920
rect 16684 9880 17132 9908
rect 15305 9871 15363 9877
rect 17126 9868 17132 9880
rect 17184 9908 17190 9920
rect 18432 9908 18460 10004
rect 20898 9976 20904 9988
rect 17184 9880 18460 9908
rect 20824 9948 20904 9976
rect 20824 9908 20852 9948
rect 20898 9936 20904 9948
rect 20956 9936 20962 9988
rect 24946 9976 24952 9988
rect 21836 9948 24952 9976
rect 21836 9908 21864 9948
rect 24946 9936 24952 9948
rect 25004 9976 25010 9988
rect 25130 9976 25136 9988
rect 25004 9948 25136 9976
rect 25004 9936 25010 9948
rect 25130 9936 25136 9948
rect 25188 9936 25194 9988
rect 20824 9880 21864 9908
rect 17184 9868 17190 9880
rect 22830 9868 22836 9920
rect 22888 9908 22894 9920
rect 23566 9908 23572 9920
rect 22888 9880 23572 9908
rect 22888 9868 22894 9880
rect 23566 9868 23572 9880
rect 23624 9868 23630 9920
rect 24210 9868 24216 9920
rect 24268 9908 24274 9920
rect 26145 9911 26203 9917
rect 26145 9908 26157 9911
rect 24268 9880 26157 9908
rect 24268 9868 24274 9880
rect 26145 9877 26157 9880
rect 26191 9877 26203 9911
rect 26145 9871 26203 9877
rect 1104 9818 28152 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 28152 9818
rect 1104 9744 28152 9766
rect 5537 9707 5595 9713
rect 5537 9673 5549 9707
rect 5583 9704 5595 9707
rect 5626 9704 5632 9716
rect 5583 9676 5632 9704
rect 5583 9673 5595 9676
rect 5537 9667 5595 9673
rect 5626 9664 5632 9676
rect 5684 9664 5690 9716
rect 8294 9704 8300 9716
rect 6932 9676 8300 9704
rect 6932 9636 6960 9676
rect 8294 9664 8300 9676
rect 8352 9664 8358 9716
rect 8754 9664 8760 9716
rect 8812 9704 8818 9716
rect 14458 9704 14464 9716
rect 8812 9676 14464 9704
rect 8812 9664 8818 9676
rect 14458 9664 14464 9676
rect 14516 9664 14522 9716
rect 14734 9664 14740 9716
rect 14792 9704 14798 9716
rect 15470 9704 15476 9716
rect 14792 9676 15476 9704
rect 14792 9664 14798 9676
rect 15470 9664 15476 9676
rect 15528 9664 15534 9716
rect 15749 9707 15807 9713
rect 15749 9673 15761 9707
rect 15795 9704 15807 9707
rect 16482 9704 16488 9716
rect 15795 9676 16488 9704
rect 15795 9673 15807 9676
rect 15749 9667 15807 9673
rect 16482 9664 16488 9676
rect 16540 9664 16546 9716
rect 17954 9664 17960 9716
rect 18012 9704 18018 9716
rect 18325 9707 18383 9713
rect 18325 9704 18337 9707
rect 18012 9676 18337 9704
rect 18012 9664 18018 9676
rect 18325 9673 18337 9676
rect 18371 9673 18383 9707
rect 18325 9667 18383 9673
rect 18874 9664 18880 9716
rect 18932 9704 18938 9716
rect 18969 9707 19027 9713
rect 18969 9704 18981 9707
rect 18932 9676 18981 9704
rect 18932 9664 18938 9676
rect 18969 9673 18981 9676
rect 19015 9673 19027 9707
rect 18969 9667 19027 9673
rect 4080 9608 4752 9636
rect 4080 9577 4108 9608
rect 4724 9580 4752 9608
rect 5368 9608 6960 9636
rect 4065 9571 4123 9577
rect 4065 9537 4077 9571
rect 4111 9537 4123 9571
rect 4065 9531 4123 9537
rect 4525 9571 4583 9577
rect 4525 9537 4537 9571
rect 4571 9537 4583 9571
rect 4525 9531 4583 9537
rect 3970 9460 3976 9512
rect 4028 9500 4034 9512
rect 4540 9500 4568 9531
rect 4706 9528 4712 9580
rect 4764 9528 4770 9580
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9537 5135 9571
rect 5077 9531 5135 9537
rect 4028 9472 4568 9500
rect 4617 9503 4675 9509
rect 4028 9460 4034 9472
rect 4617 9469 4629 9503
rect 4663 9500 4675 9503
rect 5092 9500 5120 9531
rect 5258 9528 5264 9580
rect 5316 9568 5322 9580
rect 5368 9577 5396 9608
rect 7466 9596 7472 9648
rect 7524 9596 7530 9648
rect 8202 9596 8208 9648
rect 8260 9636 8266 9648
rect 8573 9639 8631 9645
rect 8573 9636 8585 9639
rect 8260 9608 8585 9636
rect 8260 9596 8266 9608
rect 8573 9605 8585 9608
rect 8619 9605 8631 9639
rect 14642 9636 14648 9648
rect 8573 9599 8631 9605
rect 12820 9608 14648 9636
rect 5353 9571 5411 9577
rect 5353 9568 5365 9571
rect 5316 9540 5365 9568
rect 5316 9528 5322 9540
rect 5353 9537 5365 9540
rect 5399 9537 5411 9571
rect 5353 9531 5411 9537
rect 7374 9528 7380 9580
rect 7432 9528 7438 9580
rect 7561 9571 7619 9577
rect 7561 9537 7573 9571
rect 7607 9568 7619 9571
rect 7607 9540 8064 9568
rect 7607 9537 7619 9540
rect 7561 9531 7619 9537
rect 4663 9472 5120 9500
rect 4663 9469 4675 9472
rect 4617 9463 4675 9469
rect 6638 9460 6644 9512
rect 6696 9500 6702 9512
rect 7576 9500 7604 9531
rect 6696 9472 7604 9500
rect 6696 9460 6702 9472
rect 7926 9460 7932 9512
rect 7984 9460 7990 9512
rect 8036 9500 8064 9540
rect 8110 9528 8116 9580
rect 8168 9528 8174 9580
rect 12820 9577 12848 9608
rect 14642 9596 14648 9608
rect 14700 9596 14706 9648
rect 15838 9596 15844 9648
rect 15896 9636 15902 9648
rect 16209 9639 16267 9645
rect 16209 9636 16221 9639
rect 15896 9608 16221 9636
rect 15896 9596 15902 9608
rect 16209 9605 16221 9608
rect 16255 9605 16267 9639
rect 18892 9636 18920 9664
rect 16209 9599 16267 9605
rect 18156 9608 18920 9636
rect 20349 9639 20407 9645
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9568 8355 9571
rect 8389 9571 8447 9577
rect 8389 9568 8401 9571
rect 8343 9540 8401 9568
rect 8343 9537 8355 9540
rect 8297 9531 8355 9537
rect 8389 9537 8401 9540
rect 8435 9537 8447 9571
rect 8389 9531 8447 9537
rect 12805 9571 12863 9577
rect 12805 9537 12817 9571
rect 12851 9537 12863 9571
rect 12805 9531 12863 9537
rect 12894 9528 12900 9580
rect 12952 9528 12958 9580
rect 12986 9528 12992 9580
rect 13044 9528 13050 9580
rect 13262 9528 13268 9580
rect 13320 9528 13326 9580
rect 15105 9571 15163 9577
rect 15105 9537 15117 9571
rect 15151 9568 15163 9571
rect 15194 9568 15200 9580
rect 15151 9540 15200 9568
rect 15151 9537 15163 9540
rect 15105 9531 15163 9537
rect 10042 9500 10048 9512
rect 8036 9472 10048 9500
rect 10042 9460 10048 9472
rect 10100 9460 10106 9512
rect 13004 9500 13032 9528
rect 15120 9500 15148 9531
rect 15194 9528 15200 9540
rect 15252 9528 15258 9580
rect 15286 9528 15292 9580
rect 15344 9528 15350 9580
rect 15378 9528 15384 9580
rect 15436 9528 15442 9580
rect 15562 9528 15568 9580
rect 15620 9528 15626 9580
rect 16114 9528 16120 9580
rect 16172 9528 16178 9580
rect 16301 9571 16359 9577
rect 16301 9537 16313 9571
rect 16347 9568 16359 9571
rect 16850 9568 16856 9580
rect 16347 9540 16856 9568
rect 16347 9537 16359 9540
rect 16301 9531 16359 9537
rect 16850 9528 16856 9540
rect 16908 9568 16914 9580
rect 18156 9577 18184 9608
rect 20349 9605 20361 9639
rect 20395 9605 20407 9639
rect 20349 9599 20407 9605
rect 20579 9605 20637 9611
rect 18141 9571 18199 9577
rect 16908 9540 17632 9568
rect 16908 9528 16914 9540
rect 13004 9472 15148 9500
rect 16132 9500 16160 9528
rect 17604 9512 17632 9540
rect 18141 9537 18153 9571
rect 18187 9537 18199 9571
rect 18141 9531 18199 9537
rect 18877 9571 18935 9577
rect 18877 9537 18889 9571
rect 18923 9537 18935 9571
rect 18877 9531 18935 9537
rect 19061 9571 19119 9577
rect 19061 9537 19073 9571
rect 19107 9568 19119 9571
rect 19426 9568 19432 9580
rect 19107 9540 19432 9568
rect 19107 9537 19119 9540
rect 19061 9531 19119 9537
rect 16942 9500 16948 9512
rect 16132 9472 16948 9500
rect 16942 9460 16948 9472
rect 17000 9460 17006 9512
rect 17586 9460 17592 9512
rect 17644 9500 17650 9512
rect 17865 9503 17923 9509
rect 17865 9500 17877 9503
rect 17644 9472 17877 9500
rect 17644 9460 17650 9472
rect 17865 9469 17877 9472
rect 17911 9469 17923 9503
rect 17865 9463 17923 9469
rect 18230 9460 18236 9512
rect 18288 9460 18294 9512
rect 18322 9460 18328 9512
rect 18380 9460 18386 9512
rect 4433 9435 4491 9441
rect 4433 9401 4445 9435
rect 4479 9432 4491 9435
rect 5166 9432 5172 9444
rect 4479 9404 5172 9432
rect 4479 9401 4491 9404
rect 4433 9395 4491 9401
rect 5166 9392 5172 9404
rect 5224 9392 5230 9444
rect 5261 9435 5319 9441
rect 5261 9401 5273 9435
rect 5307 9432 5319 9435
rect 5350 9432 5356 9444
rect 5307 9404 5356 9432
rect 5307 9401 5319 9404
rect 5261 9395 5319 9401
rect 5350 9392 5356 9404
rect 5408 9392 5414 9444
rect 9674 9392 9680 9444
rect 9732 9432 9738 9444
rect 16850 9432 16856 9444
rect 9732 9404 16856 9432
rect 9732 9392 9738 9404
rect 16850 9392 16856 9404
rect 16908 9392 16914 9444
rect 16960 9432 16988 9460
rect 17957 9435 18015 9441
rect 17957 9432 17969 9435
rect 16960 9404 17969 9432
rect 17957 9401 17969 9404
rect 18003 9401 18015 9435
rect 17957 9395 18015 9401
rect 18892 9432 18920 9531
rect 19426 9528 19432 9540
rect 19484 9528 19490 9580
rect 20364 9500 20392 9599
rect 20579 9571 20591 9605
rect 20625 9602 20637 9605
rect 20625 9580 20668 9602
rect 20714 9596 20720 9648
rect 20772 9636 20778 9648
rect 20809 9639 20867 9645
rect 20809 9636 20821 9639
rect 20772 9608 20821 9636
rect 20772 9596 20778 9608
rect 20809 9605 20821 9608
rect 20855 9605 20867 9639
rect 20809 9599 20867 9605
rect 20625 9571 20628 9580
rect 20579 9565 20628 9571
rect 20622 9528 20628 9565
rect 20680 9528 20686 9580
rect 20898 9528 20904 9580
rect 20956 9568 20962 9580
rect 21085 9571 21143 9577
rect 21085 9568 21097 9571
rect 20956 9540 21097 9568
rect 20956 9528 20962 9540
rect 21085 9537 21097 9540
rect 21131 9568 21143 9571
rect 21450 9568 21456 9580
rect 21131 9540 21456 9568
rect 21131 9537 21143 9540
rect 21085 9531 21143 9537
rect 21450 9528 21456 9540
rect 21508 9528 21514 9580
rect 21545 9571 21603 9577
rect 21545 9537 21557 9571
rect 21591 9568 21603 9571
rect 23290 9568 23296 9580
rect 21591 9540 23296 9568
rect 21591 9537 21603 9540
rect 21545 9531 21603 9537
rect 23290 9528 23296 9540
rect 23348 9528 23354 9580
rect 24210 9528 24216 9580
rect 24268 9528 24274 9580
rect 20990 9500 20996 9512
rect 20364 9472 20996 9500
rect 20990 9460 20996 9472
rect 21048 9460 21054 9512
rect 21358 9460 21364 9512
rect 21416 9460 21422 9512
rect 19702 9432 19708 9444
rect 18892 9404 19708 9432
rect 12434 9324 12440 9376
rect 12492 9364 12498 9376
rect 12529 9367 12587 9373
rect 12529 9364 12541 9367
rect 12492 9336 12541 9364
rect 12492 9324 12498 9336
rect 12529 9333 12541 9336
rect 12575 9333 12587 9367
rect 12529 9327 12587 9333
rect 13081 9367 13139 9373
rect 13081 9333 13093 9367
rect 13127 9364 13139 9367
rect 13354 9364 13360 9376
rect 13127 9336 13360 9364
rect 13127 9333 13139 9336
rect 13081 9327 13139 9333
rect 13354 9324 13360 9336
rect 13412 9324 13418 9376
rect 14918 9324 14924 9376
rect 14976 9324 14982 9376
rect 15010 9324 15016 9376
rect 15068 9364 15074 9376
rect 15381 9367 15439 9373
rect 15381 9364 15393 9367
rect 15068 9336 15393 9364
rect 15068 9324 15074 9336
rect 15381 9333 15393 9336
rect 15427 9333 15439 9367
rect 15381 9327 15439 9333
rect 15746 9324 15752 9376
rect 15804 9364 15810 9376
rect 18892 9364 18920 9404
rect 19702 9392 19708 9404
rect 19760 9392 19766 9444
rect 20717 9435 20775 9441
rect 20717 9401 20729 9435
rect 20763 9432 20775 9435
rect 21082 9432 21088 9444
rect 20763 9404 21088 9432
rect 20763 9401 20775 9404
rect 20717 9395 20775 9401
rect 21082 9392 21088 9404
rect 21140 9432 21146 9444
rect 21269 9435 21327 9441
rect 21269 9432 21281 9435
rect 21140 9404 21281 9432
rect 21140 9392 21146 9404
rect 21269 9401 21281 9404
rect 21315 9401 21327 9435
rect 21269 9395 21327 9401
rect 15804 9336 18920 9364
rect 15804 9324 15810 9336
rect 19426 9324 19432 9376
rect 19484 9364 19490 9376
rect 20533 9367 20591 9373
rect 20533 9364 20545 9367
rect 19484 9336 20545 9364
rect 19484 9324 19490 9336
rect 20533 9333 20545 9336
rect 20579 9364 20591 9367
rect 20806 9364 20812 9376
rect 20579 9336 20812 9364
rect 20579 9333 20591 9336
rect 20533 9327 20591 9333
rect 20806 9324 20812 9336
rect 20864 9324 20870 9376
rect 21174 9324 21180 9376
rect 21232 9324 21238 9376
rect 23474 9324 23480 9376
rect 23532 9364 23538 9376
rect 23842 9364 23848 9376
rect 23532 9336 23848 9364
rect 23532 9324 23538 9336
rect 23842 9324 23848 9336
rect 23900 9364 23906 9376
rect 24305 9367 24363 9373
rect 24305 9364 24317 9367
rect 23900 9336 24317 9364
rect 23900 9324 23906 9336
rect 24305 9333 24317 9336
rect 24351 9333 24363 9367
rect 24305 9327 24363 9333
rect 1104 9274 28152 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 28152 9274
rect 1104 9200 28152 9222
rect 4433 9163 4491 9169
rect 4433 9129 4445 9163
rect 4479 9160 4491 9163
rect 4706 9160 4712 9172
rect 4479 9132 4712 9160
rect 4479 9129 4491 9132
rect 4433 9123 4491 9129
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 8113 9163 8171 9169
rect 8113 9129 8125 9163
rect 8159 9160 8171 9163
rect 8202 9160 8208 9172
rect 8159 9132 8208 9160
rect 8159 9129 8171 9132
rect 8113 9123 8171 9129
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 11790 9120 11796 9172
rect 11848 9160 11854 9172
rect 12437 9163 12495 9169
rect 12437 9160 12449 9163
rect 11848 9132 12449 9160
rect 11848 9120 11854 9132
rect 12437 9129 12449 9132
rect 12483 9129 12495 9163
rect 12437 9123 12495 9129
rect 12989 9163 13047 9169
rect 12989 9129 13001 9163
rect 13035 9160 13047 9163
rect 15378 9160 15384 9172
rect 13035 9132 15384 9160
rect 13035 9129 13047 9132
rect 12989 9123 13047 9129
rect 15378 9120 15384 9132
rect 15436 9120 15442 9172
rect 18509 9163 18567 9169
rect 18509 9129 18521 9163
rect 18555 9160 18567 9163
rect 18690 9160 18696 9172
rect 18555 9132 18696 9160
rect 18555 9129 18567 9132
rect 18509 9123 18567 9129
rect 18690 9120 18696 9132
rect 18748 9120 18754 9172
rect 20993 9163 21051 9169
rect 20993 9129 21005 9163
rect 21039 9160 21051 9163
rect 21174 9160 21180 9172
rect 21039 9132 21180 9160
rect 21039 9129 21051 9132
rect 20993 9123 21051 9129
rect 21174 9120 21180 9132
rect 21232 9120 21238 9172
rect 5258 9092 5264 9104
rect 4080 9064 5264 9092
rect 3329 9027 3387 9033
rect 3329 8993 3341 9027
rect 3375 8993 3387 9027
rect 3329 8987 3387 8993
rect 3605 9027 3663 9033
rect 3605 8993 3617 9027
rect 3651 9024 3663 9027
rect 3878 9024 3884 9036
rect 3651 8996 3884 9024
rect 3651 8993 3663 8996
rect 3605 8987 3663 8993
rect 2682 8916 2688 8968
rect 2740 8956 2746 8968
rect 3237 8959 3295 8965
rect 3237 8956 3249 8959
rect 2740 8928 3249 8956
rect 2740 8916 2746 8928
rect 3237 8925 3249 8928
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 3344 8888 3372 8987
rect 3878 8984 3884 8996
rect 3936 8984 3942 9036
rect 4080 9033 4108 9064
rect 5258 9052 5264 9064
rect 5316 9052 5322 9104
rect 11977 9095 12035 9101
rect 11977 9061 11989 9095
rect 12023 9092 12035 9095
rect 12066 9092 12072 9104
rect 12023 9064 12072 9092
rect 12023 9061 12035 9064
rect 11977 9055 12035 9061
rect 12066 9052 12072 9064
rect 12124 9052 12130 9104
rect 4065 9027 4123 9033
rect 4065 8993 4077 9027
rect 4111 8993 4123 9027
rect 4065 8987 4123 8993
rect 5166 8984 5172 9036
rect 5224 8984 5230 9036
rect 10505 9027 10563 9033
rect 10505 8993 10517 9027
rect 10551 9024 10563 9027
rect 11054 9024 11060 9036
rect 10551 8996 11060 9024
rect 10551 8993 10563 8996
rect 10505 8987 10563 8993
rect 11054 8984 11060 8996
rect 11112 8984 11118 9036
rect 18230 8984 18236 9036
rect 18288 9024 18294 9036
rect 19245 9027 19303 9033
rect 19245 9024 19257 9027
rect 18288 8996 19257 9024
rect 18288 8984 18294 8996
rect 3970 8916 3976 8968
rect 4028 8916 4034 8968
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8925 4215 8959
rect 4157 8919 4215 8925
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8956 4307 8959
rect 4706 8956 4712 8968
rect 4295 8928 4712 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 4172 8888 4200 8919
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 5261 8959 5319 8965
rect 5261 8925 5273 8959
rect 5307 8956 5319 8959
rect 5442 8956 5448 8968
rect 5307 8928 5448 8956
rect 5307 8925 5319 8928
rect 5261 8919 5319 8925
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 7926 8916 7932 8968
rect 7984 8916 7990 8968
rect 8110 8916 8116 8968
rect 8168 8916 8174 8968
rect 10226 8916 10232 8968
rect 10284 8916 10290 8968
rect 12710 8916 12716 8968
rect 12768 8916 12774 8968
rect 12802 8916 12808 8968
rect 12860 8916 12866 8968
rect 18432 8965 18460 8996
rect 19245 8993 19257 8996
rect 19291 8993 19303 9027
rect 19245 8987 19303 8993
rect 18417 8959 18475 8965
rect 18417 8925 18429 8959
rect 18463 8925 18475 8959
rect 18417 8919 18475 8925
rect 18506 8916 18512 8968
rect 18564 8916 18570 8968
rect 19426 8916 19432 8968
rect 19484 8916 19490 8968
rect 20714 8916 20720 8968
rect 20772 8916 20778 8968
rect 20806 8916 20812 8968
rect 20864 8916 20870 8968
rect 20990 8916 20996 8968
rect 21048 8916 21054 8968
rect 23474 8916 23480 8968
rect 23532 8916 23538 8968
rect 23658 8916 23664 8968
rect 23716 8916 23722 8968
rect 23937 8959 23995 8965
rect 23937 8925 23949 8959
rect 23983 8956 23995 8959
rect 25038 8956 25044 8968
rect 23983 8928 25044 8956
rect 23983 8925 23995 8928
rect 23937 8919 23995 8925
rect 25038 8916 25044 8928
rect 25096 8916 25102 8968
rect 3344 8860 4200 8888
rect 4172 8820 4200 8860
rect 5350 8848 5356 8900
rect 5408 8888 5414 8900
rect 10134 8888 10140 8900
rect 5408 8860 10140 8888
rect 5408 8848 5414 8860
rect 10134 8848 10140 8860
rect 10192 8848 10198 8900
rect 12066 8888 12072 8900
rect 11730 8860 12072 8888
rect 12066 8848 12072 8860
rect 12124 8848 12130 8900
rect 12342 8848 12348 8900
rect 12400 8848 12406 8900
rect 16850 8848 16856 8900
rect 16908 8888 16914 8900
rect 17770 8888 17776 8900
rect 16908 8860 17776 8888
rect 16908 8848 16914 8860
rect 17770 8848 17776 8860
rect 17828 8888 17834 8900
rect 18233 8891 18291 8897
rect 18233 8888 18245 8891
rect 17828 8860 18245 8888
rect 17828 8848 17834 8860
rect 18233 8857 18245 8860
rect 18279 8857 18291 8891
rect 18233 8851 18291 8857
rect 19613 8891 19671 8897
rect 19613 8857 19625 8891
rect 19659 8888 19671 8891
rect 19702 8888 19708 8900
rect 19659 8860 19708 8888
rect 19659 8857 19671 8860
rect 19613 8851 19671 8857
rect 19702 8848 19708 8860
rect 19760 8848 19766 8900
rect 24302 8888 24308 8900
rect 23768 8860 24308 8888
rect 5534 8820 5540 8832
rect 4172 8792 5540 8820
rect 5534 8780 5540 8792
rect 5592 8780 5598 8832
rect 5629 8823 5687 8829
rect 5629 8789 5641 8823
rect 5675 8820 5687 8823
rect 6914 8820 6920 8832
rect 5675 8792 6920 8820
rect 5675 8789 5687 8792
rect 5629 8783 5687 8789
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 23290 8780 23296 8832
rect 23348 8820 23354 8832
rect 23768 8829 23796 8860
rect 24302 8848 24308 8860
rect 24360 8848 24366 8900
rect 23753 8823 23811 8829
rect 23753 8820 23765 8823
rect 23348 8792 23765 8820
rect 23348 8780 23354 8792
rect 23753 8789 23765 8792
rect 23799 8789 23811 8823
rect 23753 8783 23811 8789
rect 23934 8780 23940 8832
rect 23992 8820 23998 8832
rect 24762 8820 24768 8832
rect 23992 8792 24768 8820
rect 23992 8780 23998 8792
rect 24762 8780 24768 8792
rect 24820 8780 24826 8832
rect 1104 8730 28152 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 28152 8730
rect 1104 8656 28152 8678
rect 3605 8619 3663 8625
rect 3605 8585 3617 8619
rect 3651 8616 3663 8619
rect 3970 8616 3976 8628
rect 3651 8588 3976 8616
rect 3651 8585 3663 8588
rect 3605 8579 3663 8585
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 5442 8576 5448 8628
rect 5500 8576 5506 8628
rect 6914 8576 6920 8628
rect 6972 8616 6978 8628
rect 7745 8619 7803 8625
rect 6972 8588 7696 8616
rect 6972 8576 6978 8588
rect 4614 8548 4620 8560
rect 3068 8520 3740 8548
rect 3068 8489 3096 8520
rect 3712 8489 3740 8520
rect 3804 8520 4620 8548
rect 3804 8489 3832 8520
rect 4614 8508 4620 8520
rect 4672 8508 4678 8560
rect 5258 8508 5264 8560
rect 5316 8548 5322 8560
rect 7193 8551 7251 8557
rect 5316 8520 5580 8548
rect 5316 8508 5322 8520
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 3513 8483 3571 8489
rect 3513 8449 3525 8483
rect 3559 8449 3571 8483
rect 3513 8443 3571 8449
rect 3697 8483 3755 8489
rect 3697 8449 3709 8483
rect 3743 8449 3755 8483
rect 3697 8443 3755 8449
rect 3789 8483 3847 8489
rect 3789 8449 3801 8483
rect 3835 8449 3847 8483
rect 3789 8443 3847 8449
rect 2958 8372 2964 8424
rect 3016 8412 3022 8424
rect 3528 8412 3556 8443
rect 3016 8384 3556 8412
rect 3016 8372 3022 8384
rect 3421 8347 3479 8353
rect 3421 8313 3433 8347
rect 3467 8344 3479 8347
rect 3712 8344 3740 8443
rect 3878 8440 3884 8492
rect 3936 8480 3942 8492
rect 3973 8483 4031 8489
rect 3973 8480 3985 8483
rect 3936 8452 3985 8480
rect 3936 8440 3942 8452
rect 3973 8449 3985 8452
rect 4019 8449 4031 8483
rect 3973 8443 4031 8449
rect 5350 8440 5356 8492
rect 5408 8440 5414 8492
rect 5552 8489 5580 8520
rect 7193 8517 7205 8551
rect 7239 8548 7251 8551
rect 7668 8548 7696 8588
rect 7745 8585 7757 8619
rect 7791 8616 7803 8619
rect 7926 8616 7932 8628
rect 7791 8588 7932 8616
rect 7791 8585 7803 8588
rect 7745 8579 7803 8585
rect 7926 8576 7932 8588
rect 7984 8576 7990 8628
rect 8021 8619 8079 8625
rect 8021 8585 8033 8619
rect 8067 8616 8079 8619
rect 8386 8616 8392 8628
rect 8067 8588 8392 8616
rect 8067 8585 8079 8588
rect 8021 8579 8079 8585
rect 8386 8576 8392 8588
rect 8444 8576 8450 8628
rect 10134 8576 10140 8628
rect 10192 8616 10198 8628
rect 10778 8616 10784 8628
rect 10192 8588 10784 8616
rect 10192 8576 10198 8588
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 11882 8576 11888 8628
rect 11940 8576 11946 8628
rect 14918 8576 14924 8628
rect 14976 8616 14982 8628
rect 14976 8588 16804 8616
rect 14976 8576 14982 8588
rect 10321 8551 10379 8557
rect 7239 8520 7604 8548
rect 7668 8520 7880 8548
rect 7239 8517 7251 8520
rect 7193 8511 7251 8517
rect 5537 8483 5595 8489
rect 5537 8449 5549 8483
rect 5583 8449 5595 8483
rect 5537 8443 5595 8449
rect 7006 8440 7012 8492
rect 7064 8440 7070 8492
rect 7098 8440 7104 8492
rect 7156 8480 7162 8492
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 7156 8452 7389 8480
rect 7156 8440 7162 8452
rect 7377 8449 7389 8452
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 7466 8440 7472 8492
rect 7524 8440 7530 8492
rect 7576 8489 7604 8520
rect 7852 8489 7880 8520
rect 10321 8517 10333 8551
rect 10367 8548 10379 8551
rect 11054 8548 11060 8560
rect 10367 8520 11060 8548
rect 10367 8517 10379 8520
rect 10321 8511 10379 8517
rect 11054 8508 11060 8520
rect 11112 8508 11118 8560
rect 16669 8551 16727 8557
rect 16669 8517 16681 8551
rect 16715 8517 16727 8551
rect 16776 8548 16804 8588
rect 17126 8576 17132 8628
rect 17184 8616 17190 8628
rect 17221 8619 17279 8625
rect 17221 8616 17233 8619
rect 17184 8588 17233 8616
rect 17184 8576 17190 8588
rect 17221 8585 17233 8588
rect 17267 8585 17279 8619
rect 17221 8579 17279 8585
rect 18233 8619 18291 8625
rect 18233 8585 18245 8619
rect 18279 8616 18291 8619
rect 18322 8616 18328 8628
rect 18279 8588 18328 8616
rect 18279 8585 18291 8588
rect 18233 8579 18291 8585
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 22922 8576 22928 8628
rect 22980 8616 22986 8628
rect 23017 8619 23075 8625
rect 23017 8616 23029 8619
rect 22980 8588 23029 8616
rect 22980 8576 22986 8588
rect 23017 8585 23029 8588
rect 23063 8585 23075 8619
rect 23017 8579 23075 8585
rect 24118 8576 24124 8628
rect 24176 8616 24182 8628
rect 24670 8616 24676 8628
rect 24176 8588 24676 8616
rect 24176 8576 24182 8588
rect 24670 8576 24676 8588
rect 24728 8576 24734 8628
rect 24762 8576 24768 8628
rect 24820 8616 24826 8628
rect 24820 8588 25176 8616
rect 24820 8576 24826 8588
rect 16885 8551 16943 8557
rect 16885 8548 16897 8551
rect 16776 8520 16897 8548
rect 16669 8511 16727 8517
rect 16885 8517 16897 8520
rect 16931 8548 16943 8551
rect 16931 8520 17172 8548
rect 16931 8517 16943 8520
rect 16885 8511 16943 8517
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8449 7803 8483
rect 7745 8443 7803 8449
rect 7837 8483 7895 8489
rect 7837 8449 7849 8483
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 7024 8412 7052 8440
rect 7193 8415 7251 8421
rect 7193 8412 7205 8415
rect 7024 8384 7205 8412
rect 7193 8381 7205 8384
rect 7239 8381 7251 8415
rect 7193 8375 7251 8381
rect 3881 8347 3939 8353
rect 3881 8344 3893 8347
rect 3467 8316 3648 8344
rect 3712 8316 3893 8344
rect 3467 8313 3479 8316
rect 3421 8307 3479 8313
rect 3620 8276 3648 8316
rect 3881 8313 3893 8316
rect 3927 8313 3939 8347
rect 3881 8307 3939 8313
rect 6733 8347 6791 8353
rect 6733 8313 6745 8347
rect 6779 8344 6791 8347
rect 7006 8344 7012 8356
rect 6779 8316 7012 8344
rect 6779 8313 6791 8316
rect 6733 8307 6791 8313
rect 7006 8304 7012 8316
rect 7064 8344 7070 8356
rect 7760 8344 7788 8443
rect 8018 8440 8024 8492
rect 8076 8440 8082 8492
rect 9122 8440 9128 8492
rect 9180 8440 9186 8492
rect 9306 8440 9312 8492
rect 9364 8440 9370 8492
rect 10042 8440 10048 8492
rect 10100 8440 10106 8492
rect 10502 8440 10508 8492
rect 10560 8480 10566 8492
rect 10689 8483 10747 8489
rect 10689 8480 10701 8483
rect 10560 8452 10701 8480
rect 10560 8440 10566 8452
rect 10689 8449 10701 8452
rect 10735 8449 10747 8483
rect 10689 8443 10747 8449
rect 10778 8440 10784 8492
rect 10836 8440 10842 8492
rect 11790 8440 11796 8492
rect 11848 8440 11854 8492
rect 11974 8440 11980 8492
rect 12032 8480 12038 8492
rect 12342 8480 12348 8492
rect 12032 8452 12348 8480
rect 12032 8440 12038 8452
rect 12342 8440 12348 8452
rect 12400 8440 12406 8492
rect 10413 8415 10471 8421
rect 10413 8381 10425 8415
rect 10459 8412 10471 8415
rect 10594 8412 10600 8424
rect 10459 8384 10600 8412
rect 10459 8381 10471 8384
rect 10413 8375 10471 8381
rect 10594 8372 10600 8384
rect 10652 8372 10658 8424
rect 16684 8412 16712 8511
rect 17144 8489 17172 8520
rect 23290 8508 23296 8560
rect 23348 8508 23354 8560
rect 24213 8551 24271 8557
rect 24213 8517 24225 8551
rect 24259 8548 24271 8551
rect 24933 8551 24991 8557
rect 24933 8548 24945 8551
rect 24259 8520 24945 8548
rect 24259 8517 24271 8520
rect 24213 8511 24271 8517
rect 24933 8517 24945 8520
rect 24979 8548 24991 8551
rect 25038 8548 25044 8560
rect 24979 8520 25044 8548
rect 24979 8517 24991 8520
rect 24933 8511 24991 8517
rect 25038 8508 25044 8520
rect 25096 8508 25102 8560
rect 25148 8557 25176 8588
rect 25133 8551 25191 8557
rect 25133 8517 25145 8551
rect 25179 8517 25191 8551
rect 25133 8511 25191 8517
rect 17129 8483 17187 8489
rect 17129 8449 17141 8483
rect 17175 8449 17187 8483
rect 17129 8443 17187 8449
rect 17405 8483 17463 8489
rect 17405 8449 17417 8483
rect 17451 8480 17463 8483
rect 17586 8480 17592 8492
rect 17451 8452 17592 8480
rect 17451 8449 17463 8452
rect 17405 8443 17463 8449
rect 17420 8412 17448 8443
rect 17586 8440 17592 8452
rect 17644 8440 17650 8492
rect 17865 8483 17923 8489
rect 17865 8449 17877 8483
rect 17911 8480 17923 8483
rect 18046 8480 18052 8492
rect 17911 8452 18052 8480
rect 17911 8449 17923 8452
rect 17865 8443 17923 8449
rect 18046 8440 18052 8452
rect 18104 8440 18110 8492
rect 23201 8483 23259 8489
rect 23201 8449 23213 8483
rect 23247 8449 23259 8483
rect 23201 8443 23259 8449
rect 16684 8384 17448 8412
rect 17770 8372 17776 8424
rect 17828 8372 17834 8424
rect 23216 8412 23244 8443
rect 23382 8440 23388 8492
rect 23440 8440 23446 8492
rect 23566 8440 23572 8492
rect 23624 8480 23630 8492
rect 23842 8480 23848 8492
rect 23624 8452 23848 8480
rect 23624 8440 23630 8452
rect 23842 8440 23848 8452
rect 23900 8440 23906 8492
rect 23934 8440 23940 8492
rect 23992 8440 23998 8492
rect 24044 8452 24256 8480
rect 24044 8424 24072 8452
rect 24026 8412 24032 8424
rect 23216 8384 24032 8412
rect 24026 8372 24032 8384
rect 24084 8372 24090 8424
rect 24121 8415 24179 8421
rect 24121 8381 24133 8415
rect 24167 8381 24179 8415
rect 24228 8412 24256 8452
rect 24302 8440 24308 8492
rect 24360 8440 24366 8492
rect 24489 8483 24547 8489
rect 24489 8449 24501 8483
rect 24535 8449 24547 8483
rect 24489 8443 24547 8449
rect 24504 8412 24532 8443
rect 25222 8440 25228 8492
rect 25280 8480 25286 8492
rect 27706 8480 27712 8492
rect 25280 8452 27712 8480
rect 25280 8440 25286 8452
rect 27706 8440 27712 8452
rect 27764 8440 27770 8492
rect 24228 8384 24532 8412
rect 24121 8375 24179 8381
rect 7064 8316 7788 8344
rect 9217 8347 9275 8353
rect 7064 8304 7070 8316
rect 9217 8313 9229 8347
rect 9263 8344 9275 8347
rect 9674 8344 9680 8356
rect 9263 8316 9680 8344
rect 9263 8313 9275 8316
rect 9217 8307 9275 8313
rect 9674 8304 9680 8316
rect 9732 8304 9738 8356
rect 10965 8347 11023 8353
rect 10965 8313 10977 8347
rect 11011 8344 11023 8347
rect 15194 8344 15200 8356
rect 11011 8316 15200 8344
rect 11011 8313 11023 8316
rect 10965 8307 11023 8313
rect 15194 8304 15200 8316
rect 15252 8304 15258 8356
rect 17126 8344 17132 8356
rect 16868 8316 17132 8344
rect 4706 8276 4712 8288
rect 3620 8248 4712 8276
rect 4706 8236 4712 8248
rect 4764 8236 4770 8288
rect 7101 8279 7159 8285
rect 7101 8245 7113 8279
rect 7147 8276 7159 8279
rect 7466 8276 7472 8288
rect 7147 8248 7472 8276
rect 7147 8245 7159 8248
rect 7101 8239 7159 8245
rect 7466 8236 7472 8248
rect 7524 8236 7530 8288
rect 16868 8285 16896 8316
rect 17126 8304 17132 8316
rect 17184 8304 17190 8356
rect 21082 8344 21088 8356
rect 20548 8316 21088 8344
rect 16853 8279 16911 8285
rect 16853 8245 16865 8279
rect 16899 8245 16911 8279
rect 16853 8239 16911 8245
rect 17034 8236 17040 8288
rect 17092 8236 17098 8288
rect 17402 8236 17408 8288
rect 17460 8236 17466 8288
rect 18874 8236 18880 8288
rect 18932 8276 18938 8288
rect 20548 8276 20576 8316
rect 21082 8304 21088 8316
rect 21140 8304 21146 8356
rect 23750 8304 23756 8356
rect 23808 8304 23814 8356
rect 24136 8344 24164 8375
rect 24670 8372 24676 8424
rect 24728 8412 24734 8424
rect 24728 8384 24900 8412
rect 24728 8372 24734 8384
rect 24302 8344 24308 8356
rect 24136 8316 24308 8344
rect 24302 8304 24308 8316
rect 24360 8304 24366 8356
rect 24765 8347 24823 8353
rect 24765 8344 24777 8347
rect 24412 8316 24777 8344
rect 18932 8248 20576 8276
rect 18932 8236 18938 8248
rect 24118 8236 24124 8288
rect 24176 8236 24182 8288
rect 24210 8236 24216 8288
rect 24268 8276 24274 8288
rect 24412 8276 24440 8316
rect 24765 8313 24777 8316
rect 24811 8313 24823 8347
rect 24765 8307 24823 8313
rect 24268 8248 24440 8276
rect 24268 8236 24274 8248
rect 24670 8236 24676 8288
rect 24728 8236 24734 8288
rect 24872 8276 24900 8384
rect 25130 8304 25136 8356
rect 25188 8344 25194 8356
rect 25409 8347 25467 8353
rect 25409 8344 25421 8347
rect 25188 8316 25421 8344
rect 25188 8304 25194 8316
rect 25409 8313 25421 8316
rect 25455 8313 25467 8347
rect 25409 8307 25467 8313
rect 24949 8279 25007 8285
rect 24949 8276 24961 8279
rect 24872 8248 24961 8276
rect 24949 8245 24961 8248
rect 24995 8245 25007 8279
rect 24949 8239 25007 8245
rect 1104 8186 28152 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 28152 8186
rect 1104 8112 28152 8134
rect 8481 8075 8539 8081
rect 8481 8041 8493 8075
rect 8527 8072 8539 8075
rect 9122 8072 9128 8084
rect 8527 8044 9128 8072
rect 8527 8041 8539 8044
rect 8481 8035 8539 8041
rect 9122 8032 9128 8044
rect 9180 8032 9186 8084
rect 9306 8032 9312 8084
rect 9364 8032 9370 8084
rect 11974 8032 11980 8084
rect 12032 8032 12038 8084
rect 12710 8032 12716 8084
rect 12768 8032 12774 8084
rect 15378 8032 15384 8084
rect 15436 8032 15442 8084
rect 15838 8032 15844 8084
rect 15896 8032 15902 8084
rect 16574 8032 16580 8084
rect 16632 8072 16638 8084
rect 17221 8075 17279 8081
rect 17221 8072 17233 8075
rect 16632 8044 17233 8072
rect 16632 8032 16638 8044
rect 17221 8041 17233 8044
rect 17267 8041 17279 8075
rect 17221 8035 17279 8041
rect 4341 8007 4399 8013
rect 4341 7973 4353 8007
rect 4387 8004 4399 8007
rect 5626 8004 5632 8016
rect 4387 7976 5632 8004
rect 4387 7973 4399 7976
rect 4341 7967 4399 7973
rect 5626 7964 5632 7976
rect 5684 7964 5690 8016
rect 8018 8004 8024 8016
rect 7208 7976 8024 8004
rect 3878 7896 3884 7948
rect 3936 7896 3942 7948
rect 4522 7936 4528 7948
rect 3988 7908 4528 7936
rect 3988 7877 4016 7908
rect 4522 7896 4528 7908
rect 4580 7896 4586 7948
rect 4706 7896 4712 7948
rect 4764 7896 4770 7948
rect 6914 7896 6920 7948
rect 6972 7896 6978 7948
rect 7208 7880 7236 7976
rect 8018 7964 8024 7976
rect 8076 7964 8082 8016
rect 11790 7964 11796 8016
rect 11848 8004 11854 8016
rect 17236 8004 17264 8035
rect 18322 8032 18328 8084
rect 18380 8072 18386 8084
rect 18380 8044 21496 8072
rect 18380 8032 18386 8044
rect 17862 8004 17868 8016
rect 11848 7976 13216 8004
rect 17236 7976 17868 8004
rect 11848 7964 11854 7976
rect 7377 7939 7435 7945
rect 7377 7905 7389 7939
rect 7423 7905 7435 7939
rect 11517 7939 11575 7945
rect 7377 7899 7435 7905
rect 8404 7908 9168 7936
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4338 7828 4344 7880
rect 4396 7868 4402 7880
rect 4617 7871 4675 7877
rect 4617 7868 4629 7871
rect 4396 7840 4629 7868
rect 4396 7828 4402 7840
rect 4617 7837 4629 7840
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7868 7067 7871
rect 7190 7868 7196 7880
rect 7055 7840 7196 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 7392 7868 7420 7899
rect 8404 7877 8432 7908
rect 8389 7871 8447 7877
rect 8389 7868 8401 7871
rect 7392 7840 8401 7868
rect 8389 7837 8401 7840
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 8570 7828 8576 7880
rect 8628 7868 8634 7880
rect 9140 7877 9168 7908
rect 11517 7905 11529 7939
rect 11563 7936 11575 7939
rect 11974 7936 11980 7948
rect 11563 7908 11980 7936
rect 11563 7905 11575 7908
rect 11517 7899 11575 7905
rect 11974 7896 11980 7908
rect 12032 7896 12038 7948
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8628 7840 8953 7868
rect 8628 7828 8634 7840
rect 8941 7837 8953 7840
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 9125 7871 9183 7877
rect 9125 7837 9137 7871
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 10778 7828 10784 7880
rect 10836 7868 10842 7880
rect 11425 7871 11483 7877
rect 11425 7868 11437 7871
rect 10836 7840 11437 7868
rect 10836 7828 10842 7840
rect 11425 7837 11437 7840
rect 11471 7837 11483 7871
rect 11425 7831 11483 7837
rect 11701 7871 11759 7877
rect 11701 7837 11713 7871
rect 11747 7837 11759 7871
rect 11701 7831 11759 7837
rect 11793 7871 11851 7877
rect 11793 7837 11805 7871
rect 11839 7868 11851 7871
rect 12710 7868 12716 7880
rect 11839 7840 12716 7868
rect 11839 7837 11851 7840
rect 11793 7831 11851 7837
rect 10134 7760 10140 7812
rect 10192 7800 10198 7812
rect 11716 7800 11744 7831
rect 12710 7828 12716 7840
rect 12768 7868 12774 7880
rect 13188 7877 13216 7976
rect 17862 7964 17868 7976
rect 17920 7964 17926 8016
rect 18414 7964 18420 8016
rect 18472 8004 18478 8016
rect 19242 8004 19248 8016
rect 18472 7976 19248 8004
rect 18472 7964 18478 7976
rect 19242 7964 19248 7976
rect 19300 8004 19306 8016
rect 19300 7976 20576 8004
rect 19300 7964 19306 7976
rect 13354 7896 13360 7948
rect 13412 7936 13418 7948
rect 14458 7936 14464 7948
rect 13412 7908 14464 7936
rect 13412 7896 13418 7908
rect 14458 7896 14464 7908
rect 14516 7936 14522 7948
rect 14516 7908 16988 7936
rect 14516 7896 14522 7908
rect 12897 7871 12955 7877
rect 12897 7868 12909 7871
rect 12768 7840 12909 7868
rect 12768 7828 12774 7840
rect 12897 7837 12909 7840
rect 12943 7837 12955 7871
rect 12897 7831 12955 7837
rect 12989 7871 13047 7877
rect 12989 7837 13001 7871
rect 13035 7837 13047 7871
rect 12989 7831 13047 7837
rect 13173 7871 13231 7877
rect 13173 7837 13185 7871
rect 13219 7837 13231 7871
rect 13173 7831 13231 7837
rect 13004 7800 13032 7831
rect 13262 7828 13268 7880
rect 13320 7828 13326 7880
rect 15194 7828 15200 7880
rect 15252 7868 15258 7880
rect 15381 7871 15439 7877
rect 15381 7868 15393 7871
rect 15252 7840 15393 7868
rect 15252 7828 15258 7840
rect 15381 7837 15393 7840
rect 15427 7837 15439 7871
rect 15381 7831 15439 7837
rect 15562 7828 15568 7880
rect 15620 7828 15626 7880
rect 15654 7828 15660 7880
rect 15712 7828 15718 7880
rect 16960 7877 16988 7908
rect 17034 7896 17040 7948
rect 17092 7936 17098 7948
rect 19613 7939 19671 7945
rect 17092 7908 19472 7936
rect 17092 7896 17098 7908
rect 16945 7871 17003 7877
rect 16945 7837 16957 7871
rect 16991 7837 17003 7871
rect 16945 7831 17003 7837
rect 17221 7871 17279 7877
rect 17221 7837 17233 7871
rect 17267 7868 17279 7871
rect 17402 7868 17408 7880
rect 17267 7840 17408 7868
rect 17267 7837 17279 7840
rect 17221 7831 17279 7837
rect 14274 7800 14280 7812
rect 10192 7772 14280 7800
rect 10192 7760 10198 7772
rect 14274 7760 14280 7772
rect 14332 7760 14338 7812
rect 16960 7800 16988 7831
rect 17402 7828 17408 7840
rect 17460 7828 17466 7880
rect 18046 7828 18052 7880
rect 18104 7828 18110 7880
rect 18138 7828 18144 7880
rect 18196 7828 18202 7880
rect 18322 7828 18328 7880
rect 18380 7828 18386 7880
rect 18414 7828 18420 7880
rect 18472 7828 18478 7880
rect 18506 7828 18512 7880
rect 18564 7868 18570 7880
rect 18892 7877 18920 7908
rect 18693 7871 18751 7877
rect 18693 7868 18705 7871
rect 18564 7840 18705 7868
rect 18564 7828 18570 7840
rect 18693 7837 18705 7840
rect 18739 7837 18751 7871
rect 18693 7831 18751 7837
rect 18871 7871 18929 7877
rect 18871 7837 18883 7871
rect 18917 7837 18929 7871
rect 18871 7831 18929 7837
rect 16960 7772 17448 7800
rect 4985 7735 5043 7741
rect 4985 7701 4997 7735
rect 5031 7732 5043 7735
rect 5442 7732 5448 7744
rect 5031 7704 5448 7732
rect 5031 7701 5043 7704
rect 4985 7695 5043 7701
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 12250 7692 12256 7744
rect 12308 7732 12314 7744
rect 13814 7732 13820 7744
rect 12308 7704 13820 7732
rect 12308 7692 12314 7704
rect 13814 7692 13820 7704
rect 13872 7732 13878 7744
rect 15010 7732 15016 7744
rect 13872 7704 15016 7732
rect 13872 7692 13878 7704
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 16761 7735 16819 7741
rect 16761 7701 16773 7735
rect 16807 7732 16819 7735
rect 17310 7732 17316 7744
rect 16807 7704 17316 7732
rect 16807 7701 16819 7704
rect 16761 7695 16819 7701
rect 17310 7692 17316 7704
rect 17368 7692 17374 7744
rect 17420 7732 17448 7772
rect 17678 7760 17684 7812
rect 17736 7800 17742 7812
rect 18340 7800 18368 7828
rect 17736 7772 18368 7800
rect 17736 7760 17742 7772
rect 18506 7732 18512 7744
rect 17420 7704 18512 7732
rect 18506 7692 18512 7704
rect 18564 7692 18570 7744
rect 18598 7692 18604 7744
rect 18656 7692 18662 7744
rect 18708 7732 18736 7831
rect 19242 7828 19248 7880
rect 19300 7828 19306 7880
rect 19444 7877 19472 7908
rect 19613 7905 19625 7939
rect 19659 7936 19671 7939
rect 20070 7936 20076 7948
rect 19659 7908 20076 7936
rect 19659 7905 19671 7908
rect 19613 7899 19671 7905
rect 20070 7896 20076 7908
rect 20128 7896 20134 7948
rect 20548 7880 20576 7976
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7837 19487 7871
rect 19429 7831 19487 7837
rect 19702 7828 19708 7880
rect 19760 7828 19766 7880
rect 19797 7871 19855 7877
rect 19797 7837 19809 7871
rect 19843 7868 19855 7871
rect 20438 7868 20444 7880
rect 19843 7840 20444 7868
rect 19843 7837 19855 7840
rect 19797 7831 19855 7837
rect 20438 7828 20444 7840
rect 20496 7828 20502 7880
rect 20530 7828 20536 7880
rect 20588 7828 20594 7880
rect 20640 7877 20668 8044
rect 21269 8007 21327 8013
rect 21269 7973 21281 8007
rect 21315 8004 21327 8007
rect 21358 8004 21364 8016
rect 21315 7976 21364 8004
rect 21315 7973 21327 7976
rect 21269 7967 21327 7973
rect 21358 7964 21364 7976
rect 21416 7964 21422 8016
rect 21468 8004 21496 8044
rect 21818 8032 21824 8084
rect 21876 8072 21882 8084
rect 22554 8072 22560 8084
rect 21876 8044 22560 8072
rect 21876 8032 21882 8044
rect 22554 8032 22560 8044
rect 22612 8032 22618 8084
rect 24026 8032 24032 8084
rect 24084 8072 24090 8084
rect 24121 8075 24179 8081
rect 24121 8072 24133 8075
rect 24084 8044 24133 8072
rect 24084 8032 24090 8044
rect 24121 8041 24133 8044
rect 24167 8041 24179 8075
rect 24121 8035 24179 8041
rect 25038 8032 25044 8084
rect 25096 8072 25102 8084
rect 26145 8075 26203 8081
rect 26145 8072 26157 8075
rect 25096 8044 26157 8072
rect 25096 8032 25102 8044
rect 26145 8041 26157 8044
rect 26191 8041 26203 8075
rect 26145 8035 26203 8041
rect 22922 8004 22928 8016
rect 21468 7976 22928 8004
rect 22922 7964 22928 7976
rect 22980 7964 22986 8016
rect 21634 7936 21640 7948
rect 21192 7908 21640 7936
rect 21192 7880 21220 7908
rect 21634 7896 21640 7908
rect 21692 7896 21698 7948
rect 22002 7896 22008 7948
rect 22060 7936 22066 7948
rect 22060 7908 23980 7936
rect 22060 7896 22066 7908
rect 20625 7871 20683 7877
rect 20625 7837 20637 7871
rect 20671 7837 20683 7871
rect 20625 7831 20683 7837
rect 20806 7828 20812 7880
rect 20864 7828 20870 7880
rect 20898 7828 20904 7880
rect 20956 7828 20962 7880
rect 21174 7828 21180 7880
rect 21232 7828 21238 7880
rect 21358 7828 21364 7880
rect 21416 7828 21422 7880
rect 21450 7828 21456 7880
rect 21508 7868 21514 7880
rect 22738 7868 22744 7880
rect 21508 7840 22744 7868
rect 21508 7828 21514 7840
rect 22738 7828 22744 7840
rect 22796 7868 22802 7880
rect 22833 7871 22891 7877
rect 22833 7868 22845 7871
rect 22796 7840 22845 7868
rect 22796 7828 22802 7840
rect 22833 7837 22845 7840
rect 22879 7837 22891 7871
rect 22833 7831 22891 7837
rect 23382 7828 23388 7880
rect 23440 7868 23446 7880
rect 23661 7871 23719 7877
rect 23661 7868 23673 7871
rect 23440 7840 23673 7868
rect 23440 7828 23446 7840
rect 23661 7837 23673 7840
rect 23707 7837 23719 7871
rect 23661 7831 23719 7837
rect 23842 7828 23848 7880
rect 23900 7828 23906 7880
rect 23952 7877 23980 7908
rect 24394 7896 24400 7948
rect 24452 7896 24458 7948
rect 24670 7896 24676 7948
rect 24728 7896 24734 7948
rect 23937 7871 23995 7877
rect 23937 7837 23949 7871
rect 23983 7837 23995 7871
rect 23937 7831 23995 7837
rect 24118 7828 24124 7880
rect 24176 7828 24182 7880
rect 18785 7803 18843 7809
rect 18785 7769 18797 7803
rect 18831 7800 18843 7803
rect 19978 7800 19984 7812
rect 18831 7772 19984 7800
rect 18831 7769 18843 7772
rect 18785 7763 18843 7769
rect 19978 7760 19984 7772
rect 20036 7760 20042 7812
rect 20162 7760 20168 7812
rect 20220 7800 20226 7812
rect 21468 7800 21496 7828
rect 20220 7772 21496 7800
rect 20220 7760 20226 7772
rect 21726 7760 21732 7812
rect 21784 7760 21790 7812
rect 22646 7760 22652 7812
rect 22704 7800 22710 7812
rect 23293 7803 23351 7809
rect 23293 7800 23305 7803
rect 22704 7772 23305 7800
rect 22704 7760 22710 7772
rect 23293 7769 23305 7772
rect 23339 7769 23351 7803
rect 23293 7763 23351 7769
rect 25130 7760 25136 7812
rect 25188 7760 25194 7812
rect 19242 7732 19248 7744
rect 18708 7704 19248 7732
rect 19242 7692 19248 7704
rect 19300 7692 19306 7744
rect 20254 7692 20260 7744
rect 20312 7732 20318 7744
rect 20349 7735 20407 7741
rect 20349 7732 20361 7735
rect 20312 7704 20361 7732
rect 20312 7692 20318 7704
rect 20349 7701 20361 7704
rect 20395 7701 20407 7735
rect 20349 7695 20407 7701
rect 20806 7692 20812 7744
rect 20864 7732 20870 7744
rect 20993 7735 21051 7741
rect 20993 7732 21005 7735
rect 20864 7704 21005 7732
rect 20864 7692 20870 7704
rect 20993 7701 21005 7704
rect 21039 7701 21051 7735
rect 20993 7695 21051 7701
rect 21082 7692 21088 7744
rect 21140 7732 21146 7744
rect 21818 7732 21824 7744
rect 21140 7704 21824 7732
rect 21140 7692 21146 7704
rect 21818 7692 21824 7704
rect 21876 7692 21882 7744
rect 23014 7692 23020 7744
rect 23072 7692 23078 7744
rect 23474 7692 23480 7744
rect 23532 7692 23538 7744
rect 1104 7642 28152 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 28152 7642
rect 1104 7568 28152 7590
rect 4338 7488 4344 7540
rect 4396 7488 4402 7540
rect 6457 7531 6515 7537
rect 6457 7497 6469 7531
rect 6503 7528 6515 7531
rect 7282 7528 7288 7540
rect 6503 7500 7288 7528
rect 6503 7497 6515 7500
rect 6457 7491 6515 7497
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 9582 7528 9588 7540
rect 9324 7500 9588 7528
rect 6641 7463 6699 7469
rect 6641 7429 6653 7463
rect 6687 7460 6699 7463
rect 6825 7463 6883 7469
rect 6825 7460 6837 7463
rect 6687 7432 6837 7460
rect 6687 7429 6699 7432
rect 6641 7423 6699 7429
rect 6825 7429 6837 7432
rect 6871 7429 6883 7463
rect 6825 7423 6883 7429
rect 8386 7420 8392 7472
rect 8444 7460 8450 7472
rect 9324 7469 9352 7500
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 11241 7531 11299 7537
rect 11241 7497 11253 7531
rect 11287 7528 11299 7531
rect 14182 7528 14188 7540
rect 11287 7500 14188 7528
rect 11287 7497 11299 7500
rect 11241 7491 11299 7497
rect 14182 7488 14188 7500
rect 14240 7488 14246 7540
rect 15562 7488 15568 7540
rect 15620 7528 15626 7540
rect 15657 7531 15715 7537
rect 15657 7528 15669 7531
rect 15620 7500 15669 7528
rect 15620 7488 15626 7500
rect 15657 7497 15669 7500
rect 15703 7497 15715 7531
rect 15657 7491 15715 7497
rect 17494 7488 17500 7540
rect 17552 7528 17558 7540
rect 17957 7531 18015 7537
rect 17957 7528 17969 7531
rect 17552 7500 17969 7528
rect 17552 7488 17558 7500
rect 17957 7497 17969 7500
rect 18003 7497 18015 7531
rect 17957 7491 18015 7497
rect 18506 7488 18512 7540
rect 18564 7528 18570 7540
rect 20993 7531 21051 7537
rect 18564 7500 20392 7528
rect 18564 7488 18570 7500
rect 8665 7463 8723 7469
rect 8665 7460 8677 7463
rect 8444 7432 8677 7460
rect 8444 7420 8450 7432
rect 8665 7429 8677 7432
rect 8711 7429 8723 7463
rect 8665 7423 8723 7429
rect 9309 7463 9367 7469
rect 9309 7429 9321 7463
rect 9355 7429 9367 7463
rect 9309 7423 9367 7429
rect 9766 7420 9772 7472
rect 9824 7420 9830 7472
rect 10042 7420 10048 7472
rect 10100 7460 10106 7472
rect 11609 7463 11667 7469
rect 10100 7432 11560 7460
rect 10100 7420 10106 7432
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 5258 7392 5264 7404
rect 4387 7364 5264 7392
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 4172 7324 4200 7355
rect 5258 7352 5264 7364
rect 5316 7352 5322 7404
rect 6270 7352 6276 7404
rect 6328 7392 6334 7404
rect 6365 7395 6423 7401
rect 6365 7392 6377 7395
rect 6328 7364 6377 7392
rect 6328 7352 6334 7364
rect 6365 7361 6377 7364
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 5534 7324 5540 7336
rect 4172 7296 5540 7324
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 5626 7284 5632 7336
rect 5684 7324 5690 7336
rect 6748 7324 6776 7355
rect 6914 7352 6920 7404
rect 6972 7352 6978 7404
rect 8202 7352 8208 7404
rect 8260 7392 8266 7404
rect 8481 7395 8539 7401
rect 8481 7392 8493 7395
rect 8260 7364 8493 7392
rect 8260 7352 8266 7364
rect 8481 7361 8493 7364
rect 8527 7361 8539 7395
rect 8481 7355 8539 7361
rect 8849 7395 8907 7401
rect 8849 7361 8861 7395
rect 8895 7392 8907 7395
rect 8941 7395 8999 7401
rect 8941 7392 8953 7395
rect 8895 7364 8953 7392
rect 8895 7361 8907 7364
rect 8849 7355 8907 7361
rect 8941 7361 8953 7364
rect 8987 7361 8999 7395
rect 8941 7355 8999 7361
rect 9122 7352 9128 7404
rect 9180 7352 9186 7404
rect 9398 7352 9404 7404
rect 9456 7352 9462 7404
rect 9585 7395 9643 7401
rect 9585 7361 9597 7395
rect 9631 7361 9643 7395
rect 9585 7355 9643 7361
rect 5684 7296 6776 7324
rect 5684 7284 5690 7296
rect 8570 7284 8576 7336
rect 8628 7324 8634 7336
rect 9600 7324 9628 7355
rect 10318 7352 10324 7404
rect 10376 7392 10382 7404
rect 10689 7395 10747 7401
rect 10689 7392 10701 7395
rect 10376 7364 10701 7392
rect 10376 7352 10382 7364
rect 10689 7361 10701 7364
rect 10735 7361 10747 7395
rect 10689 7355 10747 7361
rect 10778 7352 10784 7404
rect 10836 7352 10842 7404
rect 10962 7352 10968 7404
rect 11020 7352 11026 7404
rect 11054 7352 11060 7404
rect 11112 7352 11118 7404
rect 11532 7401 11560 7432
rect 11609 7429 11621 7463
rect 11655 7460 11667 7463
rect 11790 7460 11796 7472
rect 11655 7432 11796 7460
rect 11655 7429 11667 7432
rect 11609 7423 11667 7429
rect 11790 7420 11796 7432
rect 11848 7420 11854 7472
rect 12161 7463 12219 7469
rect 12161 7429 12173 7463
rect 12207 7429 12219 7463
rect 12161 7423 12219 7429
rect 12377 7463 12435 7469
rect 12377 7429 12389 7463
rect 12423 7460 12435 7463
rect 12894 7460 12900 7472
rect 12423 7432 12900 7460
rect 12423 7429 12435 7432
rect 12377 7423 12435 7429
rect 11517 7395 11575 7401
rect 11517 7361 11529 7395
rect 11563 7361 11575 7395
rect 11517 7355 11575 7361
rect 11701 7395 11759 7401
rect 11701 7361 11713 7395
rect 11747 7392 11759 7395
rect 11747 7364 11928 7392
rect 11747 7361 11759 7364
rect 11701 7355 11759 7361
rect 8628 7296 9628 7324
rect 8628 7284 8634 7296
rect 11900 7268 11928 7364
rect 11974 7352 11980 7404
rect 12032 7392 12038 7404
rect 12176 7392 12204 7423
rect 12894 7420 12900 7432
rect 12952 7420 12958 7472
rect 14274 7420 14280 7472
rect 14332 7460 14338 7472
rect 15219 7463 15277 7469
rect 14332 7432 14964 7460
rect 14332 7420 14338 7432
rect 12032 7364 12204 7392
rect 12032 7352 12038 7364
rect 12618 7352 12624 7404
rect 12676 7392 12682 7404
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12676 7364 13001 7392
rect 12676 7352 12682 7364
rect 12989 7361 13001 7364
rect 13035 7392 13047 7395
rect 13262 7392 13268 7404
rect 13035 7364 13268 7392
rect 13035 7361 13047 7364
rect 12989 7355 13047 7361
rect 13262 7352 13268 7364
rect 13320 7352 13326 7404
rect 14461 7395 14519 7401
rect 14461 7361 14473 7395
rect 14507 7392 14519 7395
rect 14550 7392 14556 7404
rect 14507 7364 14556 7392
rect 14507 7361 14519 7364
rect 14461 7355 14519 7361
rect 14550 7352 14556 7364
rect 14608 7352 14614 7404
rect 14734 7352 14740 7404
rect 14792 7352 14798 7404
rect 14826 7352 14832 7404
rect 14884 7352 14890 7404
rect 14936 7401 14964 7432
rect 15219 7429 15231 7463
rect 15265 7460 15277 7463
rect 15378 7460 15384 7472
rect 15265 7432 15384 7460
rect 15265 7429 15277 7432
rect 15219 7423 15277 7429
rect 15378 7420 15384 7432
rect 15436 7420 15442 7472
rect 16114 7460 16120 7472
rect 15856 7432 16120 7460
rect 14921 7395 14979 7401
rect 14921 7361 14933 7395
rect 14967 7361 14979 7395
rect 15856 7392 15884 7432
rect 16114 7420 16120 7432
rect 16172 7460 16178 7472
rect 16209 7463 16267 7469
rect 16209 7460 16221 7463
rect 16172 7432 16221 7460
rect 16172 7420 16178 7432
rect 16209 7429 16221 7432
rect 16255 7429 16267 7463
rect 16209 7423 16267 7429
rect 18046 7420 18052 7472
rect 18104 7460 18110 7472
rect 18782 7460 18788 7472
rect 18104 7432 18788 7460
rect 18104 7420 18110 7432
rect 18782 7420 18788 7432
rect 18840 7460 18846 7472
rect 18840 7432 19012 7460
rect 18840 7420 18846 7432
rect 14921 7355 14979 7361
rect 15120 7364 15884 7392
rect 15933 7395 15991 7401
rect 11992 7296 14596 7324
rect 11882 7216 11888 7268
rect 11940 7216 11946 7268
rect 5902 7148 5908 7200
rect 5960 7188 5966 7200
rect 6641 7191 6699 7197
rect 6641 7188 6653 7191
rect 5960 7160 6653 7188
rect 5960 7148 5966 7160
rect 6641 7157 6653 7160
rect 6687 7157 6699 7191
rect 6641 7151 6699 7157
rect 9766 7148 9772 7200
rect 9824 7188 9830 7200
rect 11992 7188 12020 7296
rect 12710 7256 12716 7268
rect 12360 7228 12716 7256
rect 12360 7197 12388 7228
rect 12710 7216 12716 7228
rect 12768 7216 12774 7268
rect 12986 7216 12992 7268
rect 13044 7256 13050 7268
rect 13354 7256 13360 7268
rect 13044 7228 13360 7256
rect 13044 7216 13050 7228
rect 13354 7216 13360 7228
rect 13412 7216 13418 7268
rect 14568 7256 14596 7296
rect 14642 7284 14648 7336
rect 14700 7284 14706 7336
rect 15120 7333 15148 7364
rect 15933 7361 15945 7395
rect 15979 7392 15991 7395
rect 17405 7395 17463 7401
rect 15979 7364 17356 7392
rect 15979 7361 15991 7364
rect 15933 7355 15991 7361
rect 15105 7327 15163 7333
rect 15105 7293 15117 7327
rect 15151 7293 15163 7327
rect 15105 7287 15163 7293
rect 15120 7256 15148 7287
rect 15746 7284 15752 7336
rect 15804 7324 15810 7336
rect 15841 7327 15899 7333
rect 15841 7324 15853 7327
rect 15804 7296 15853 7324
rect 15804 7284 15810 7296
rect 15841 7293 15853 7296
rect 15887 7293 15899 7327
rect 16301 7327 16359 7333
rect 16301 7324 16313 7327
rect 15841 7287 15899 7293
rect 16224 7296 16313 7324
rect 14568 7228 15148 7256
rect 15289 7259 15347 7265
rect 15289 7225 15301 7259
rect 15335 7256 15347 7259
rect 16224 7256 16252 7296
rect 16301 7293 16313 7296
rect 16347 7324 16359 7327
rect 16758 7324 16764 7336
rect 16347 7296 16764 7324
rect 16347 7293 16359 7296
rect 16301 7287 16359 7293
rect 16758 7284 16764 7296
rect 16816 7284 16822 7336
rect 15335 7228 16252 7256
rect 17328 7256 17356 7364
rect 17405 7361 17417 7395
rect 17451 7392 17463 7395
rect 17586 7392 17592 7404
rect 17451 7364 17592 7392
rect 17451 7361 17463 7364
rect 17405 7355 17463 7361
rect 17586 7352 17592 7364
rect 17644 7352 17650 7404
rect 17865 7395 17923 7401
rect 17865 7361 17877 7395
rect 17911 7392 17923 7395
rect 17954 7392 17960 7404
rect 17911 7364 17960 7392
rect 17911 7361 17923 7364
rect 17865 7355 17923 7361
rect 17954 7352 17960 7364
rect 18012 7352 18018 7404
rect 18598 7352 18604 7404
rect 18656 7352 18662 7404
rect 18984 7401 19012 7432
rect 20364 7404 20392 7500
rect 20993 7497 21005 7531
rect 21039 7528 21051 7531
rect 21082 7528 21088 7540
rect 21039 7500 21088 7528
rect 21039 7497 21051 7500
rect 20993 7491 21051 7497
rect 21082 7488 21088 7500
rect 21140 7488 21146 7540
rect 21358 7488 21364 7540
rect 21416 7528 21422 7540
rect 21637 7531 21695 7537
rect 21637 7528 21649 7531
rect 21416 7500 21649 7528
rect 21416 7488 21422 7500
rect 21637 7497 21649 7500
rect 21683 7497 21695 7531
rect 21637 7491 21695 7497
rect 21910 7488 21916 7540
rect 21968 7528 21974 7540
rect 23017 7531 23075 7537
rect 23017 7528 23029 7531
rect 21968 7500 23029 7528
rect 21968 7488 21974 7500
rect 23017 7497 23029 7500
rect 23063 7497 23075 7531
rect 23017 7491 23075 7497
rect 23109 7531 23167 7537
rect 23109 7497 23121 7531
rect 23155 7528 23167 7531
rect 24210 7528 24216 7540
rect 23155 7500 24216 7528
rect 23155 7497 23167 7500
rect 23109 7491 23167 7497
rect 24210 7488 24216 7500
rect 24268 7488 24274 7540
rect 21821 7463 21879 7469
rect 21821 7460 21833 7463
rect 20548 7432 21833 7460
rect 20548 7404 20576 7432
rect 21821 7429 21833 7432
rect 21867 7429 21879 7463
rect 22189 7463 22247 7469
rect 22189 7460 22201 7463
rect 21821 7423 21879 7429
rect 21928 7432 22201 7460
rect 18969 7395 19027 7401
rect 18969 7361 18981 7395
rect 19015 7361 19027 7395
rect 18969 7355 19027 7361
rect 19889 7395 19947 7401
rect 19889 7361 19901 7395
rect 19935 7392 19947 7395
rect 20162 7392 20168 7404
rect 19935 7364 20168 7392
rect 19935 7361 19947 7364
rect 19889 7355 19947 7361
rect 20162 7352 20168 7364
rect 20220 7352 20226 7404
rect 20346 7352 20352 7404
rect 20404 7352 20410 7404
rect 20438 7352 20444 7404
rect 20496 7352 20502 7404
rect 20530 7352 20536 7404
rect 20588 7352 20594 7404
rect 20717 7395 20775 7401
rect 20717 7361 20729 7395
rect 20763 7361 20775 7395
rect 20717 7355 20775 7361
rect 18693 7327 18751 7333
rect 18693 7293 18705 7327
rect 18739 7293 18751 7327
rect 18693 7287 18751 7293
rect 18708 7256 18736 7287
rect 18874 7284 18880 7336
rect 18932 7284 18938 7336
rect 19702 7284 19708 7336
rect 19760 7324 19766 7336
rect 20254 7324 20260 7336
rect 19760 7296 20260 7324
rect 19760 7284 19766 7296
rect 20254 7284 20260 7296
rect 20312 7324 20318 7336
rect 20732 7324 20760 7355
rect 20806 7352 20812 7404
rect 20864 7352 20870 7404
rect 20990 7352 20996 7404
rect 21048 7392 21054 7404
rect 21269 7395 21327 7401
rect 21269 7392 21281 7395
rect 21048 7364 21281 7392
rect 21048 7352 21054 7364
rect 21269 7361 21281 7364
rect 21315 7392 21327 7395
rect 21542 7392 21548 7404
rect 21315 7364 21548 7392
rect 21315 7361 21327 7364
rect 21269 7355 21327 7361
rect 21542 7352 21548 7364
rect 21600 7352 21606 7404
rect 21177 7327 21235 7333
rect 21177 7324 21189 7327
rect 20312 7296 20760 7324
rect 20824 7296 21189 7324
rect 20312 7284 20318 7296
rect 19613 7259 19671 7265
rect 19613 7256 19625 7259
rect 17328 7228 18644 7256
rect 18708 7228 19625 7256
rect 15335 7225 15347 7228
rect 15289 7219 15347 7225
rect 9824 7160 12020 7188
rect 12345 7191 12403 7197
rect 9824 7148 9830 7160
rect 12345 7157 12357 7191
rect 12391 7157 12403 7191
rect 12345 7151 12403 7157
rect 12526 7148 12532 7200
rect 12584 7148 12590 7200
rect 12802 7148 12808 7200
rect 12860 7188 12866 7200
rect 12897 7191 12955 7197
rect 12897 7188 12909 7191
rect 12860 7160 12909 7188
rect 12860 7148 12866 7160
rect 12897 7157 12909 7160
rect 12943 7157 12955 7191
rect 12897 7151 12955 7157
rect 14366 7148 14372 7200
rect 14424 7188 14430 7200
rect 14461 7191 14519 7197
rect 14461 7188 14473 7191
rect 14424 7160 14473 7188
rect 14424 7148 14430 7160
rect 14461 7157 14473 7160
rect 14507 7188 14519 7191
rect 15013 7191 15071 7197
rect 15013 7188 15025 7191
rect 14507 7160 15025 7188
rect 14507 7157 14519 7160
rect 14461 7151 14519 7157
rect 15013 7157 15025 7160
rect 15059 7157 15071 7191
rect 15013 7151 15071 7157
rect 17497 7191 17555 7197
rect 17497 7157 17509 7191
rect 17543 7188 17555 7191
rect 18046 7188 18052 7200
rect 17543 7160 18052 7188
rect 17543 7157 17555 7160
rect 17497 7151 17555 7157
rect 18046 7148 18052 7160
rect 18104 7148 18110 7200
rect 18616 7188 18644 7228
rect 19613 7225 19625 7228
rect 19659 7225 19671 7259
rect 19613 7219 19671 7225
rect 19978 7216 19984 7268
rect 20036 7216 20042 7268
rect 20070 7216 20076 7268
rect 20128 7256 20134 7268
rect 20714 7256 20720 7268
rect 20128 7228 20720 7256
rect 20128 7216 20134 7228
rect 20714 7216 20720 7228
rect 20772 7256 20778 7268
rect 20824 7256 20852 7296
rect 21177 7293 21189 7296
rect 21223 7293 21235 7327
rect 21177 7287 21235 7293
rect 20772 7228 20852 7256
rect 20772 7216 20778 7228
rect 20898 7216 20904 7268
rect 20956 7256 20962 7268
rect 21928 7256 21956 7432
rect 22189 7429 22201 7432
rect 22235 7429 22247 7463
rect 22189 7423 22247 7429
rect 22738 7420 22744 7472
rect 22796 7420 22802 7472
rect 22922 7420 22928 7472
rect 22980 7420 22986 7472
rect 23768 7432 24348 7460
rect 22002 7352 22008 7404
rect 22060 7352 22066 7404
rect 22281 7395 22339 7401
rect 22281 7361 22293 7395
rect 22327 7392 22339 7395
rect 22554 7392 22560 7404
rect 22327 7364 22560 7392
rect 22327 7361 22339 7364
rect 22281 7355 22339 7361
rect 22554 7352 22560 7364
rect 22612 7352 22618 7404
rect 23768 7401 23796 7432
rect 24320 7404 24348 7432
rect 22649 7395 22707 7401
rect 22649 7361 22661 7395
rect 22695 7361 22707 7395
rect 22649 7355 22707 7361
rect 23753 7395 23811 7401
rect 23753 7361 23765 7395
rect 23799 7361 23811 7395
rect 23753 7355 23811 7361
rect 20956 7228 21956 7256
rect 22465 7259 22523 7265
rect 20956 7216 20962 7228
rect 22465 7225 22477 7259
rect 22511 7256 22523 7259
rect 22554 7256 22560 7268
rect 22511 7228 22560 7256
rect 22511 7225 22523 7228
rect 22465 7219 22523 7225
rect 22554 7216 22560 7228
rect 22612 7216 22618 7268
rect 19334 7188 19340 7200
rect 18616 7160 19340 7188
rect 19334 7148 19340 7160
rect 19392 7148 19398 7200
rect 19702 7148 19708 7200
rect 19760 7188 19766 7200
rect 20165 7191 20223 7197
rect 20165 7188 20177 7191
rect 19760 7160 20177 7188
rect 19760 7148 19766 7160
rect 20165 7157 20177 7160
rect 20211 7157 20223 7191
rect 22664 7188 22692 7355
rect 24210 7352 24216 7404
rect 24268 7352 24274 7404
rect 24302 7352 24308 7404
rect 24360 7352 24366 7404
rect 23382 7284 23388 7336
rect 23440 7284 23446 7336
rect 23845 7327 23903 7333
rect 23845 7293 23857 7327
rect 23891 7324 23903 7327
rect 24118 7324 24124 7336
rect 23891 7296 24124 7324
rect 23891 7293 23903 7296
rect 23845 7287 23903 7293
rect 23293 7259 23351 7265
rect 23293 7225 23305 7259
rect 23339 7256 23351 7259
rect 23860 7256 23888 7287
rect 24118 7284 24124 7296
rect 24176 7284 24182 7336
rect 27614 7256 27620 7268
rect 23339 7228 23888 7256
rect 23952 7228 27620 7256
rect 23339 7225 23351 7228
rect 23293 7219 23351 7225
rect 23952 7188 23980 7228
rect 27614 7216 27620 7228
rect 27672 7216 27678 7268
rect 22664 7160 23980 7188
rect 20165 7151 20223 7157
rect 24026 7148 24032 7200
rect 24084 7148 24090 7200
rect 1104 7098 28152 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 28152 7098
rect 1104 7024 28152 7046
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 5592 6956 7880 6984
rect 5592 6944 5598 6956
rect 5442 6876 5448 6928
rect 5500 6876 5506 6928
rect 5626 6808 5632 6860
rect 5684 6848 5690 6860
rect 5997 6851 6055 6857
rect 5684 6820 5948 6848
rect 5684 6808 5690 6820
rect 5169 6783 5227 6789
rect 5169 6749 5181 6783
rect 5215 6780 5227 6783
rect 5810 6780 5816 6792
rect 5215 6752 5816 6780
rect 5215 6749 5227 6752
rect 5169 6743 5227 6749
rect 5810 6740 5816 6752
rect 5868 6740 5874 6792
rect 5920 6789 5948 6820
rect 5997 6817 6009 6851
rect 6043 6817 6055 6851
rect 5997 6811 6055 6817
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6749 5963 6783
rect 5905 6743 5963 6749
rect 6012 6712 6040 6811
rect 6270 6808 6276 6860
rect 6328 6808 6334 6860
rect 6380 6857 6408 6956
rect 7852 6925 7880 6956
rect 8570 6944 8576 6996
rect 8628 6984 8634 6996
rect 8665 6987 8723 6993
rect 8665 6984 8677 6987
rect 8628 6956 8677 6984
rect 8628 6944 8634 6956
rect 8665 6953 8677 6956
rect 8711 6953 8723 6987
rect 8665 6947 8723 6953
rect 9309 6987 9367 6993
rect 9309 6953 9321 6987
rect 9355 6984 9367 6987
rect 9398 6984 9404 6996
rect 9355 6956 9404 6984
rect 9355 6953 9367 6956
rect 9309 6947 9367 6953
rect 9398 6944 9404 6956
rect 9456 6944 9462 6996
rect 10413 6987 10471 6993
rect 10413 6953 10425 6987
rect 10459 6984 10471 6987
rect 10502 6984 10508 6996
rect 10459 6956 10508 6984
rect 10459 6953 10471 6956
rect 10413 6947 10471 6953
rect 10502 6944 10508 6956
rect 10560 6944 10566 6996
rect 10778 6944 10784 6996
rect 10836 6944 10842 6996
rect 11164 6956 12020 6984
rect 7377 6919 7435 6925
rect 7377 6885 7389 6919
rect 7423 6885 7435 6919
rect 7377 6879 7435 6885
rect 7837 6919 7895 6925
rect 7837 6885 7849 6919
rect 7883 6916 7895 6919
rect 10042 6916 10048 6928
rect 7883 6888 10048 6916
rect 7883 6885 7895 6888
rect 7837 6879 7895 6885
rect 6365 6851 6423 6857
rect 6365 6817 6377 6851
rect 6411 6817 6423 6851
rect 6365 6811 6423 6817
rect 6454 6808 6460 6860
rect 6512 6848 6518 6860
rect 6917 6851 6975 6857
rect 6917 6848 6929 6851
rect 6512 6820 6929 6848
rect 6512 6808 6518 6820
rect 6917 6817 6929 6820
rect 6963 6817 6975 6851
rect 7392 6848 7420 6879
rect 8941 6851 8999 6857
rect 8941 6848 8953 6851
rect 7392 6820 8953 6848
rect 6917 6811 6975 6817
rect 6549 6783 6607 6789
rect 6549 6749 6561 6783
rect 6595 6780 6607 6783
rect 6638 6780 6644 6792
rect 6595 6752 6644 6780
rect 6595 6749 6607 6752
rect 6549 6743 6607 6749
rect 6638 6740 6644 6752
rect 6696 6740 6702 6792
rect 6733 6783 6791 6789
rect 6733 6749 6745 6783
rect 6779 6780 6791 6783
rect 7009 6783 7067 6789
rect 7009 6780 7021 6783
rect 6779 6752 7021 6780
rect 6779 6749 6791 6752
rect 6733 6743 6791 6749
rect 7009 6749 7021 6752
rect 7055 6780 7067 6783
rect 7098 6780 7104 6792
rect 7055 6752 7104 6780
rect 7055 6749 7067 6752
rect 7009 6743 7067 6749
rect 7098 6740 7104 6752
rect 7156 6740 7162 6792
rect 8202 6740 8208 6792
rect 8260 6740 8266 6792
rect 8386 6740 8392 6792
rect 8444 6740 8450 6792
rect 8496 6789 8524 6820
rect 8941 6817 8953 6820
rect 8987 6817 8999 6851
rect 8941 6811 8999 6817
rect 8481 6783 8539 6789
rect 8481 6749 8493 6783
rect 8527 6749 8539 6783
rect 8481 6743 8539 6749
rect 8665 6783 8723 6789
rect 8665 6749 8677 6783
rect 8711 6780 8723 6783
rect 9122 6780 9128 6792
rect 8711 6752 9128 6780
rect 8711 6749 8723 6752
rect 8665 6743 8723 6749
rect 6914 6712 6920 6724
rect 6012 6684 6920 6712
rect 6914 6672 6920 6684
rect 6972 6672 6978 6724
rect 7558 6672 7564 6724
rect 7616 6712 7622 6724
rect 8297 6715 8355 6721
rect 7616 6684 8248 6712
rect 7616 6672 7622 6684
rect 5629 6647 5687 6653
rect 5629 6613 5641 6647
rect 5675 6644 5687 6647
rect 6638 6644 6644 6656
rect 5675 6616 6644 6644
rect 5675 6613 5687 6616
rect 5629 6607 5687 6613
rect 6638 6604 6644 6616
rect 6696 6604 6702 6656
rect 8220 6644 8248 6684
rect 8297 6681 8309 6715
rect 8343 6712 8355 6715
rect 8680 6712 8708 6743
rect 9122 6740 9128 6752
rect 9180 6740 9186 6792
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6780 9459 6783
rect 9508 6780 9536 6888
rect 10042 6876 10048 6888
rect 10100 6876 10106 6928
rect 10796 6848 10824 6944
rect 11054 6848 11060 6860
rect 10428 6820 10824 6848
rect 10888 6820 11060 6848
rect 9447 6752 9536 6780
rect 9585 6783 9643 6789
rect 9447 6749 9459 6752
rect 9401 6743 9459 6749
rect 9585 6749 9597 6783
rect 9631 6780 9643 6783
rect 10134 6780 10140 6792
rect 9631 6752 10140 6780
rect 9631 6749 9643 6752
rect 9585 6743 9643 6749
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10428 6789 10456 6820
rect 10413 6783 10471 6789
rect 10413 6749 10425 6783
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 10689 6783 10747 6789
rect 10689 6749 10701 6783
rect 10735 6780 10747 6783
rect 10888 6780 10916 6820
rect 11054 6808 11060 6820
rect 11112 6808 11118 6860
rect 10735 6752 10916 6780
rect 10965 6783 11023 6789
rect 10735 6749 10747 6752
rect 10689 6743 10747 6749
rect 10965 6749 10977 6783
rect 11011 6780 11023 6783
rect 11164 6780 11192 6956
rect 11238 6876 11244 6928
rect 11296 6916 11302 6928
rect 11882 6916 11888 6928
rect 11296 6888 11888 6916
rect 11296 6876 11302 6888
rect 11882 6876 11888 6888
rect 11940 6876 11946 6928
rect 11011 6752 11192 6780
rect 11241 6783 11299 6789
rect 11011 6749 11023 6752
rect 10965 6743 11023 6749
rect 11241 6749 11253 6783
rect 11287 6780 11299 6783
rect 11422 6780 11428 6792
rect 11287 6752 11428 6780
rect 11287 6749 11299 6752
rect 11241 6743 11299 6749
rect 11422 6740 11428 6752
rect 11480 6740 11486 6792
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6749 11575 6783
rect 11517 6743 11575 6749
rect 11609 6783 11667 6789
rect 11609 6749 11621 6783
rect 11655 6780 11667 6783
rect 11698 6780 11704 6792
rect 11655 6752 11704 6780
rect 11655 6749 11667 6752
rect 11609 6743 11667 6749
rect 10318 6712 10324 6724
rect 8343 6684 8708 6712
rect 9416 6684 10324 6712
rect 8343 6681 8355 6684
rect 8297 6675 8355 6681
rect 9416 6644 9444 6684
rect 10318 6672 10324 6684
rect 10376 6672 10382 6724
rect 11146 6672 11152 6724
rect 11204 6672 11210 6724
rect 11532 6712 11560 6743
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 11790 6740 11796 6792
rect 11848 6740 11854 6792
rect 11900 6789 11928 6876
rect 11992 6857 12020 6956
rect 14274 6944 14280 6996
rect 14332 6944 14338 6996
rect 17678 6984 17684 6996
rect 14660 6956 17684 6984
rect 13078 6876 13084 6928
rect 13136 6916 13142 6928
rect 13136 6888 13308 6916
rect 13136 6876 13142 6888
rect 11977 6851 12035 6857
rect 11977 6817 11989 6851
rect 12023 6848 12035 6851
rect 12250 6848 12256 6860
rect 12023 6820 12256 6848
rect 12023 6817 12035 6820
rect 11977 6811 12035 6817
rect 12250 6808 12256 6820
rect 12308 6808 12314 6860
rect 12342 6808 12348 6860
rect 12400 6848 12406 6860
rect 12529 6851 12587 6857
rect 12529 6848 12541 6851
rect 12400 6820 12541 6848
rect 12400 6808 12406 6820
rect 12529 6817 12541 6820
rect 12575 6817 12587 6851
rect 12529 6811 12587 6817
rect 12618 6808 12624 6860
rect 12676 6848 12682 6860
rect 12713 6851 12771 6857
rect 12713 6848 12725 6851
rect 12676 6820 12725 6848
rect 12676 6808 12682 6820
rect 12713 6817 12725 6820
rect 12759 6817 12771 6851
rect 12713 6811 12771 6817
rect 11885 6783 11943 6789
rect 11885 6749 11897 6783
rect 11931 6749 11943 6783
rect 11885 6743 11943 6749
rect 12069 6783 12127 6789
rect 12069 6749 12081 6783
rect 12115 6780 12127 6783
rect 12158 6780 12164 6792
rect 12115 6752 12164 6780
rect 12115 6749 12127 6752
rect 12069 6743 12127 6749
rect 12158 6740 12164 6752
rect 12216 6740 12222 6792
rect 12437 6783 12495 6789
rect 12437 6780 12449 6783
rect 12360 6752 12449 6780
rect 12360 6724 12388 6752
rect 12437 6749 12449 6752
rect 12483 6749 12495 6783
rect 12437 6743 12495 6749
rect 12802 6740 12808 6792
rect 12860 6780 12866 6792
rect 13173 6783 13231 6789
rect 12860 6774 13032 6780
rect 13071 6777 13129 6783
rect 13071 6774 13083 6777
rect 12860 6752 13083 6774
rect 12860 6740 12866 6752
rect 13004 6746 13083 6752
rect 13071 6743 13083 6746
rect 13117 6743 13129 6777
rect 13173 6749 13185 6783
rect 13219 6782 13231 6783
rect 13280 6782 13308 6888
rect 13354 6876 13360 6928
rect 13412 6916 13418 6928
rect 14660 6916 14688 6956
rect 15197 6919 15255 6925
rect 15197 6916 15209 6919
rect 13412 6888 14688 6916
rect 14752 6888 15209 6916
rect 13412 6876 13418 6888
rect 14752 6860 14780 6888
rect 15197 6885 15209 6888
rect 15243 6885 15255 6919
rect 15197 6879 15255 6885
rect 14734 6808 14740 6860
rect 14792 6808 14798 6860
rect 14826 6808 14832 6860
rect 14884 6848 14890 6860
rect 14884 6820 14964 6848
rect 14884 6808 14890 6820
rect 13219 6754 13308 6782
rect 13219 6749 13231 6754
rect 13173 6743 13231 6749
rect 13071 6737 13129 6743
rect 13354 6740 13360 6792
rect 13412 6740 13418 6792
rect 13446 6740 13452 6792
rect 13504 6740 13510 6792
rect 14090 6740 14096 6792
rect 14148 6780 14154 6792
rect 14185 6783 14243 6789
rect 14185 6780 14197 6783
rect 14148 6752 14197 6780
rect 14148 6740 14154 6752
rect 14185 6749 14197 6752
rect 14231 6780 14243 6783
rect 14461 6783 14519 6789
rect 14461 6780 14473 6783
rect 14231 6752 14473 6780
rect 14231 6749 14243 6752
rect 14185 6743 14243 6749
rect 14461 6749 14473 6752
rect 14507 6749 14519 6783
rect 14461 6743 14519 6749
rect 14550 6740 14556 6792
rect 14608 6740 14614 6792
rect 14752 6780 14780 6808
rect 14936 6789 14964 6820
rect 15488 6789 15516 6956
rect 17678 6944 17684 6956
rect 17736 6944 17742 6996
rect 17862 6944 17868 6996
rect 17920 6984 17926 6996
rect 17920 6956 18552 6984
rect 17920 6944 17926 6956
rect 16206 6916 16212 6928
rect 15580 6888 16212 6916
rect 14921 6783 14979 6789
rect 14752 6752 14872 6780
rect 11532 6684 11652 6712
rect 11624 6656 11652 6684
rect 12342 6672 12348 6724
rect 12400 6672 12406 6724
rect 13630 6672 13636 6724
rect 13688 6672 13694 6724
rect 13814 6672 13820 6724
rect 13872 6712 13878 6724
rect 14734 6712 14740 6724
rect 13872 6684 14740 6712
rect 13872 6672 13878 6684
rect 14734 6672 14740 6684
rect 14792 6672 14798 6724
rect 14844 6721 14872 6752
rect 14921 6749 14933 6783
rect 14967 6749 14979 6783
rect 15381 6783 15439 6789
rect 15381 6780 15393 6783
rect 14921 6743 14979 6749
rect 15028 6752 15393 6780
rect 14829 6715 14887 6721
rect 14829 6681 14841 6715
rect 14875 6681 14887 6715
rect 14829 6675 14887 6681
rect 8220 6616 9444 6644
rect 9490 6604 9496 6656
rect 9548 6604 9554 6656
rect 10597 6647 10655 6653
rect 10597 6613 10609 6647
rect 10643 6644 10655 6647
rect 10962 6644 10968 6656
rect 10643 6616 10968 6644
rect 10643 6613 10655 6616
rect 10597 6607 10655 6613
rect 10962 6604 10968 6616
rect 11020 6644 11026 6656
rect 11333 6647 11391 6653
rect 11333 6644 11345 6647
rect 11020 6616 11345 6644
rect 11020 6604 11026 6616
rect 11333 6613 11345 6616
rect 11379 6613 11391 6647
rect 11333 6607 11391 6613
rect 11606 6604 11612 6656
rect 11664 6604 11670 6656
rect 11698 6604 11704 6656
rect 11756 6644 11762 6656
rect 13354 6644 13360 6656
rect 11756 6616 13360 6644
rect 11756 6604 11762 6616
rect 13354 6604 13360 6616
rect 13412 6604 13418 6656
rect 13538 6604 13544 6656
rect 13596 6644 13602 6656
rect 15028 6644 15056 6752
rect 15381 6749 15393 6752
rect 15427 6749 15439 6783
rect 15381 6743 15439 6749
rect 15473 6783 15531 6789
rect 15473 6749 15485 6783
rect 15519 6749 15531 6783
rect 15473 6743 15531 6749
rect 15396 6712 15424 6743
rect 15580 6712 15608 6888
rect 16206 6876 16212 6888
rect 16264 6916 16270 6928
rect 18414 6916 18420 6928
rect 16264 6888 18420 6916
rect 16264 6876 16270 6888
rect 15933 6851 15991 6857
rect 15933 6848 15945 6851
rect 15764 6820 15945 6848
rect 15764 6792 15792 6820
rect 15933 6817 15945 6820
rect 15979 6817 15991 6851
rect 15933 6811 15991 6817
rect 16758 6808 16764 6860
rect 16816 6808 16822 6860
rect 17221 6851 17279 6857
rect 17221 6817 17233 6851
rect 17267 6848 17279 6851
rect 17497 6851 17555 6857
rect 17497 6848 17509 6851
rect 17267 6820 17509 6848
rect 17267 6817 17279 6820
rect 17221 6811 17279 6817
rect 17497 6817 17509 6820
rect 17543 6817 17555 6851
rect 17497 6811 17555 6817
rect 15654 6740 15660 6792
rect 15712 6740 15718 6792
rect 15746 6740 15752 6792
rect 15804 6740 15810 6792
rect 15838 6740 15844 6792
rect 15896 6740 15902 6792
rect 16666 6740 16672 6792
rect 16724 6740 16730 6792
rect 17034 6740 17040 6792
rect 17092 6740 17098 6792
rect 17310 6740 17316 6792
rect 17368 6740 17374 6792
rect 17696 6789 17724 6888
rect 18414 6876 18420 6888
rect 18472 6876 18478 6928
rect 18524 6916 18552 6956
rect 18782 6944 18788 6996
rect 18840 6944 18846 6996
rect 19334 6944 19340 6996
rect 19392 6984 19398 6996
rect 19429 6987 19487 6993
rect 19429 6984 19441 6987
rect 19392 6956 19441 6984
rect 19392 6944 19398 6956
rect 19429 6953 19441 6956
rect 19475 6984 19487 6987
rect 20054 6987 20112 6993
rect 20054 6984 20066 6987
rect 19475 6956 20066 6984
rect 19475 6953 19487 6956
rect 19429 6947 19487 6953
rect 20054 6953 20066 6956
rect 20100 6953 20112 6987
rect 20054 6947 20112 6953
rect 21542 6944 21548 6996
rect 21600 6944 21606 6996
rect 21726 6944 21732 6996
rect 21784 6984 21790 6996
rect 21821 6987 21879 6993
rect 21821 6984 21833 6987
rect 21784 6956 21833 6984
rect 21784 6944 21790 6956
rect 21821 6953 21833 6956
rect 21867 6953 21879 6987
rect 21821 6947 21879 6953
rect 22728 6987 22786 6993
rect 22728 6953 22740 6987
rect 22774 6984 22786 6987
rect 23474 6984 23480 6996
rect 22774 6956 23480 6984
rect 22774 6953 22786 6956
rect 22728 6947 22786 6953
rect 23474 6944 23480 6956
rect 23532 6944 23538 6996
rect 24213 6987 24271 6993
rect 24213 6953 24225 6987
rect 24259 6984 24271 6987
rect 24302 6984 24308 6996
rect 24259 6956 24308 6984
rect 24259 6953 24271 6956
rect 24213 6947 24271 6953
rect 24302 6944 24308 6956
rect 24360 6944 24366 6996
rect 19702 6916 19708 6928
rect 18524 6888 19708 6916
rect 19702 6876 19708 6888
rect 19760 6876 19766 6928
rect 18138 6848 18144 6860
rect 17972 6820 18144 6848
rect 17681 6783 17739 6789
rect 17681 6749 17693 6783
rect 17727 6749 17739 6783
rect 17681 6743 17739 6749
rect 17770 6740 17776 6792
rect 17828 6740 17834 6792
rect 17972 6789 18000 6820
rect 18138 6808 18144 6820
rect 18196 6808 18202 6860
rect 19797 6851 19855 6857
rect 19797 6817 19809 6851
rect 19843 6848 19855 6851
rect 22465 6851 22523 6857
rect 22465 6848 22477 6851
rect 19843 6820 22477 6848
rect 19843 6817 19855 6820
rect 19797 6811 19855 6817
rect 22465 6817 22477 6820
rect 22511 6848 22523 6851
rect 24394 6848 24400 6860
rect 22511 6820 24400 6848
rect 22511 6817 22523 6820
rect 22465 6811 22523 6817
rect 24394 6808 24400 6820
rect 24452 6808 24458 6860
rect 17957 6783 18015 6789
rect 17957 6749 17969 6783
rect 18003 6749 18015 6783
rect 17957 6743 18015 6749
rect 15396 6684 15608 6712
rect 15672 6712 15700 6740
rect 17972 6712 18000 6743
rect 18046 6740 18052 6792
rect 18104 6740 18110 6792
rect 18322 6740 18328 6792
rect 18380 6740 18386 6792
rect 18414 6740 18420 6792
rect 18472 6780 18478 6792
rect 18601 6783 18659 6789
rect 18601 6780 18613 6783
rect 18472 6752 18613 6780
rect 18472 6740 18478 6752
rect 18601 6749 18613 6752
rect 18647 6780 18659 6783
rect 18782 6780 18788 6792
rect 18647 6752 18788 6780
rect 18647 6749 18659 6752
rect 18601 6743 18659 6749
rect 18782 6740 18788 6752
rect 18840 6740 18846 6792
rect 18877 6783 18935 6789
rect 18877 6749 18889 6783
rect 18923 6780 18935 6783
rect 19242 6780 19248 6792
rect 18923 6752 19248 6780
rect 18923 6749 18935 6752
rect 18877 6743 18935 6749
rect 19242 6740 19248 6752
rect 19300 6740 19306 6792
rect 19426 6740 19432 6792
rect 19484 6740 19490 6792
rect 19610 6740 19616 6792
rect 19668 6740 19674 6792
rect 19705 6783 19763 6789
rect 19705 6749 19717 6783
rect 19751 6749 19763 6783
rect 19705 6743 19763 6749
rect 15672 6684 18000 6712
rect 18064 6712 18092 6740
rect 18509 6715 18567 6721
rect 18509 6712 18521 6715
rect 18064 6684 18521 6712
rect 18509 6681 18521 6684
rect 18555 6681 18567 6715
rect 18509 6675 18567 6681
rect 13596 6616 15056 6644
rect 13596 6604 13602 6616
rect 15102 6604 15108 6656
rect 15160 6604 15166 6656
rect 16666 6604 16672 6656
rect 16724 6644 16730 6656
rect 18141 6647 18199 6653
rect 18141 6644 18153 6647
rect 16724 6616 18153 6644
rect 16724 6604 16730 6616
rect 18141 6613 18153 6616
rect 18187 6613 18199 6647
rect 19720 6644 19748 6743
rect 22002 6740 22008 6792
rect 22060 6740 22066 6792
rect 25130 6712 25136 6724
rect 21298 6684 22094 6712
rect 23966 6684 25136 6712
rect 20806 6644 20812 6656
rect 19720 6616 20812 6644
rect 18141 6607 18199 6613
rect 20806 6604 20812 6616
rect 20864 6604 20870 6656
rect 22066 6644 22094 6684
rect 24044 6644 24072 6684
rect 25130 6672 25136 6684
rect 25188 6672 25194 6724
rect 22066 6616 24072 6644
rect 1104 6554 28152 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 28152 6554
rect 1104 6480 28152 6502
rect 6181 6443 6239 6449
rect 6181 6409 6193 6443
rect 6227 6440 6239 6443
rect 6454 6440 6460 6452
rect 6227 6412 6460 6440
rect 6227 6409 6239 6412
rect 6181 6403 6239 6409
rect 6454 6400 6460 6412
rect 6512 6400 6518 6452
rect 6549 6443 6607 6449
rect 6549 6409 6561 6443
rect 6595 6440 6607 6443
rect 7098 6440 7104 6452
rect 6595 6412 7104 6440
rect 6595 6409 6607 6412
rect 6549 6403 6607 6409
rect 7098 6400 7104 6412
rect 7156 6400 7162 6452
rect 11054 6400 11060 6452
rect 11112 6440 11118 6452
rect 11793 6443 11851 6449
rect 11793 6440 11805 6443
rect 11112 6412 11805 6440
rect 11112 6400 11118 6412
rect 11793 6409 11805 6412
rect 11839 6409 11851 6443
rect 11793 6403 11851 6409
rect 12158 6400 12164 6452
rect 12216 6440 12222 6452
rect 13170 6440 13176 6452
rect 12216 6412 13176 6440
rect 12216 6400 12222 6412
rect 13170 6400 13176 6412
rect 13228 6400 13234 6452
rect 14826 6400 14832 6452
rect 14884 6400 14890 6452
rect 15289 6443 15347 6449
rect 15289 6409 15301 6443
rect 15335 6440 15347 6443
rect 15746 6440 15752 6452
rect 15335 6412 15752 6440
rect 15335 6409 15347 6412
rect 15289 6403 15347 6409
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 17494 6400 17500 6452
rect 17552 6400 17558 6452
rect 17862 6400 17868 6452
rect 17920 6400 17926 6452
rect 19153 6443 19211 6449
rect 19153 6409 19165 6443
rect 19199 6440 19211 6443
rect 19242 6440 19248 6452
rect 19199 6412 19248 6440
rect 19199 6409 19211 6412
rect 19153 6403 19211 6409
rect 19242 6400 19248 6412
rect 19300 6400 19306 6452
rect 19426 6400 19432 6452
rect 19484 6440 19490 6452
rect 20530 6440 20536 6452
rect 19484 6412 20536 6440
rect 19484 6400 19490 6412
rect 20530 6400 20536 6412
rect 20588 6400 20594 6452
rect 20898 6400 20904 6452
rect 20956 6440 20962 6452
rect 20993 6443 21051 6449
rect 20993 6440 21005 6443
rect 20956 6412 21005 6440
rect 20956 6400 20962 6412
rect 20993 6409 21005 6412
rect 21039 6409 21051 6443
rect 20993 6403 21051 6409
rect 22002 6400 22008 6452
rect 22060 6440 22066 6452
rect 23017 6443 23075 6449
rect 23017 6440 23029 6443
rect 22060 6412 23029 6440
rect 22060 6400 22066 6412
rect 23017 6409 23029 6412
rect 23063 6409 23075 6443
rect 23017 6403 23075 6409
rect 27614 6400 27620 6452
rect 27672 6400 27678 6452
rect 6917 6375 6975 6381
rect 6917 6341 6929 6375
rect 6963 6372 6975 6375
rect 7190 6372 7196 6384
rect 6963 6344 7196 6372
rect 6963 6341 6975 6344
rect 6917 6335 6975 6341
rect 7190 6332 7196 6344
rect 7248 6332 7254 6384
rect 11974 6332 11980 6384
rect 12032 6372 12038 6384
rect 12621 6375 12679 6381
rect 12621 6372 12633 6375
rect 12032 6344 12633 6372
rect 12032 6332 12038 6344
rect 12621 6341 12633 6344
rect 12667 6341 12679 6375
rect 12621 6335 12679 6341
rect 12710 6332 12716 6384
rect 12768 6372 12774 6384
rect 12805 6375 12863 6381
rect 12805 6372 12817 6375
rect 12768 6344 12817 6372
rect 12768 6332 12774 6344
rect 12805 6341 12817 6344
rect 12851 6372 12863 6375
rect 14274 6372 14280 6384
rect 12851 6344 14280 6372
rect 12851 6341 12863 6344
rect 12805 6335 12863 6341
rect 5442 6264 5448 6316
rect 5500 6304 5506 6316
rect 5813 6307 5871 6313
rect 5813 6304 5825 6307
rect 5500 6276 5825 6304
rect 5500 6264 5506 6276
rect 5813 6273 5825 6276
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 6454 6264 6460 6316
rect 6512 6264 6518 6316
rect 6638 6264 6644 6316
rect 6696 6304 6702 6316
rect 6733 6307 6791 6313
rect 6733 6304 6745 6307
rect 6696 6276 6745 6304
rect 6696 6264 6702 6276
rect 6733 6273 6745 6276
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 7282 6264 7288 6316
rect 7340 6304 7346 6316
rect 9490 6304 9496 6316
rect 7340 6276 9496 6304
rect 7340 6264 7346 6276
rect 9490 6264 9496 6276
rect 9548 6264 9554 6316
rect 12069 6307 12127 6313
rect 12069 6273 12081 6307
rect 12115 6273 12127 6307
rect 12069 6267 12127 6273
rect 12253 6307 12311 6313
rect 12253 6273 12265 6307
rect 12299 6304 12311 6307
rect 12434 6304 12440 6316
rect 12299 6276 12440 6304
rect 12299 6273 12311 6276
rect 12253 6267 12311 6273
rect 5902 6196 5908 6248
rect 5960 6196 5966 6248
rect 6270 6196 6276 6248
rect 6328 6236 6334 6248
rect 7193 6239 7251 6245
rect 7193 6236 7205 6239
rect 6328 6208 7205 6236
rect 6328 6196 6334 6208
rect 7193 6205 7205 6208
rect 7239 6205 7251 6239
rect 7193 6199 7251 6205
rect 7653 6239 7711 6245
rect 7653 6205 7665 6239
rect 7699 6236 7711 6239
rect 8386 6236 8392 6248
rect 7699 6208 8392 6236
rect 7699 6205 7711 6208
rect 7653 6199 7711 6205
rect 8386 6196 8392 6208
rect 8444 6196 8450 6248
rect 12084 6236 12112 6267
rect 12434 6264 12440 6276
rect 12492 6264 12498 6316
rect 12529 6307 12587 6313
rect 12529 6273 12541 6307
rect 12575 6304 12587 6307
rect 12575 6276 12848 6304
rect 12575 6273 12587 6276
rect 12529 6267 12587 6273
rect 12820 6236 12848 6276
rect 12894 6264 12900 6316
rect 12952 6304 12958 6316
rect 13832 6313 13860 6344
rect 14274 6332 14280 6344
rect 14332 6332 14338 6384
rect 14550 6332 14556 6384
rect 14608 6372 14614 6384
rect 14921 6375 14979 6381
rect 14921 6372 14933 6375
rect 14608 6344 14933 6372
rect 14608 6332 14614 6344
rect 14921 6341 14933 6344
rect 14967 6341 14979 6375
rect 17512 6372 17540 6400
rect 17681 6375 17739 6381
rect 17681 6372 17693 6375
rect 17512 6344 17693 6372
rect 14921 6335 14979 6341
rect 17681 6341 17693 6344
rect 17727 6341 17739 6375
rect 17880 6372 17908 6400
rect 17880 6344 18170 6372
rect 17681 6335 17739 6341
rect 13817 6307 13875 6313
rect 12952 6276 13768 6304
rect 12952 6264 12958 6276
rect 12986 6236 12992 6248
rect 12084 6208 12756 6236
rect 12820 6208 12992 6236
rect 12161 6171 12219 6177
rect 12161 6137 12173 6171
rect 12207 6168 12219 6171
rect 12621 6171 12679 6177
rect 12621 6168 12633 6171
rect 12207 6140 12633 6168
rect 12207 6137 12219 6140
rect 12161 6131 12219 6137
rect 12621 6137 12633 6140
rect 12667 6137 12679 6171
rect 12728 6168 12756 6208
rect 12986 6196 12992 6208
rect 13044 6196 13050 6248
rect 13740 6245 13768 6276
rect 13817 6273 13829 6307
rect 13863 6273 13875 6307
rect 14449 6307 14507 6313
rect 14449 6304 14461 6307
rect 13817 6267 13875 6273
rect 14200 6276 14461 6304
rect 13725 6239 13783 6245
rect 13725 6205 13737 6239
rect 13771 6205 13783 6239
rect 13725 6199 13783 6205
rect 13814 6168 13820 6180
rect 12728 6140 13820 6168
rect 12621 6131 12679 6137
rect 13814 6128 13820 6140
rect 13872 6128 13878 6180
rect 14200 6177 14228 6276
rect 14449 6273 14461 6276
rect 14495 6273 14507 6307
rect 14449 6267 14507 6273
rect 15102 6264 15108 6316
rect 15160 6264 15166 6316
rect 15378 6264 15384 6316
rect 15436 6304 15442 6316
rect 16390 6304 16396 6316
rect 15436 6276 16396 6304
rect 15436 6264 15442 6276
rect 16390 6264 16396 6276
rect 16448 6264 16454 6316
rect 21085 6307 21143 6313
rect 21085 6273 21097 6307
rect 21131 6304 21143 6307
rect 21542 6304 21548 6316
rect 21131 6276 21548 6304
rect 21131 6273 21143 6276
rect 21085 6267 21143 6273
rect 21542 6264 21548 6276
rect 21600 6264 21606 6316
rect 22925 6307 22983 6313
rect 22925 6273 22937 6307
rect 22971 6304 22983 6307
rect 23014 6304 23020 6316
rect 22971 6276 23020 6304
rect 22971 6273 22983 6276
rect 22925 6267 22983 6273
rect 23014 6264 23020 6276
rect 23072 6264 23078 6316
rect 27798 6264 27804 6316
rect 27856 6264 27862 6316
rect 14550 6196 14556 6248
rect 14608 6196 14614 6248
rect 17218 6196 17224 6248
rect 17276 6236 17282 6248
rect 17405 6239 17463 6245
rect 17405 6236 17417 6239
rect 17276 6208 17417 6236
rect 17276 6196 17282 6208
rect 17405 6205 17417 6208
rect 17451 6205 17463 6239
rect 17405 6199 17463 6205
rect 17678 6196 17684 6248
rect 17736 6236 17742 6248
rect 24026 6236 24032 6248
rect 17736 6208 24032 6236
rect 17736 6196 17742 6208
rect 24026 6196 24032 6208
rect 24084 6196 24090 6248
rect 14185 6171 14243 6177
rect 14185 6137 14197 6171
rect 14231 6137 14243 6171
rect 14185 6131 14243 6137
rect 14274 6128 14280 6180
rect 14332 6168 14338 6180
rect 15838 6168 15844 6180
rect 14332 6140 15844 6168
rect 14332 6128 14338 6140
rect 15838 6128 15844 6140
rect 15896 6128 15902 6180
rect 16574 6168 16580 6180
rect 16132 6140 16580 6168
rect 12342 6060 12348 6112
rect 12400 6060 12406 6112
rect 14642 6060 14648 6112
rect 14700 6100 14706 6112
rect 16132 6100 16160 6140
rect 16574 6128 16580 6140
rect 16632 6128 16638 6180
rect 14700 6072 16160 6100
rect 14700 6060 14706 6072
rect 16390 6060 16396 6112
rect 16448 6100 16454 6112
rect 18414 6100 18420 6112
rect 16448 6072 18420 6100
rect 16448 6060 16454 6072
rect 18414 6060 18420 6072
rect 18472 6060 18478 6112
rect 18690 6060 18696 6112
rect 18748 6100 18754 6112
rect 23014 6100 23020 6112
rect 18748 6072 23020 6100
rect 18748 6060 18754 6072
rect 23014 6060 23020 6072
rect 23072 6060 23078 6112
rect 1104 6010 28152 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 28152 6010
rect 1104 5936 28152 5958
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7374 5896 7380 5908
rect 6972 5868 7380 5896
rect 6972 5856 6978 5868
rect 7374 5856 7380 5868
rect 7432 5896 7438 5908
rect 8662 5896 8668 5908
rect 7432 5868 8668 5896
rect 7432 5856 7438 5868
rect 8662 5856 8668 5868
rect 8720 5896 8726 5908
rect 8720 5868 11560 5896
rect 8720 5856 8726 5868
rect 11532 5828 11560 5868
rect 11974 5856 11980 5908
rect 12032 5856 12038 5908
rect 12618 5856 12624 5908
rect 12676 5896 12682 5908
rect 15378 5896 15384 5908
rect 12676 5868 15384 5896
rect 12676 5856 12682 5868
rect 15378 5856 15384 5868
rect 15436 5856 15442 5908
rect 15838 5856 15844 5908
rect 15896 5856 15902 5908
rect 17586 5856 17592 5908
rect 17644 5896 17650 5908
rect 17957 5899 18015 5905
rect 17957 5896 17969 5899
rect 17644 5868 17969 5896
rect 17644 5856 17650 5868
rect 17957 5865 17969 5868
rect 18003 5865 18015 5899
rect 17957 5859 18015 5865
rect 27617 5899 27675 5905
rect 27617 5865 27629 5899
rect 27663 5896 27675 5899
rect 27706 5896 27712 5908
rect 27663 5868 27712 5896
rect 27663 5865 27675 5868
rect 27617 5859 27675 5865
rect 27706 5856 27712 5868
rect 27764 5856 27770 5908
rect 13998 5828 14004 5840
rect 11532 5800 14004 5828
rect 13998 5788 14004 5800
rect 14056 5788 14062 5840
rect 10226 5720 10232 5772
rect 10284 5760 10290 5772
rect 11514 5760 11520 5772
rect 10284 5732 11520 5760
rect 10284 5720 10290 5732
rect 11514 5720 11520 5732
rect 11572 5760 11578 5772
rect 14093 5763 14151 5769
rect 14093 5760 14105 5763
rect 11572 5732 14105 5760
rect 11572 5720 11578 5732
rect 14093 5729 14105 5732
rect 14139 5760 14151 5763
rect 16209 5763 16267 5769
rect 16209 5760 16221 5763
rect 14139 5732 16221 5760
rect 14139 5729 14151 5732
rect 14093 5723 14151 5729
rect 16209 5729 16221 5732
rect 16255 5760 16267 5763
rect 17218 5760 17224 5772
rect 16255 5732 17224 5760
rect 16255 5729 16267 5732
rect 16209 5723 16267 5729
rect 17218 5720 17224 5732
rect 17276 5720 17282 5772
rect 27522 5652 27528 5704
rect 27580 5692 27586 5704
rect 27801 5695 27859 5701
rect 27801 5692 27813 5695
rect 27580 5664 27813 5692
rect 27580 5652 27586 5664
rect 27801 5661 27813 5664
rect 27847 5661 27859 5695
rect 27801 5655 27859 5661
rect 10502 5584 10508 5636
rect 10560 5584 10566 5636
rect 12066 5624 12072 5636
rect 11730 5596 12072 5624
rect 12066 5584 12072 5596
rect 12124 5624 12130 5636
rect 13078 5624 13084 5636
rect 12124 5596 13084 5624
rect 12124 5584 12130 5596
rect 13078 5584 13084 5596
rect 13136 5584 13142 5636
rect 14366 5584 14372 5636
rect 14424 5584 14430 5636
rect 16485 5627 16543 5633
rect 15594 5596 15700 5624
rect 15672 5568 15700 5596
rect 16485 5593 16497 5627
rect 16531 5624 16543 5627
rect 16758 5624 16764 5636
rect 16531 5596 16764 5624
rect 16531 5593 16543 5596
rect 16485 5587 16543 5593
rect 16758 5584 16764 5596
rect 16816 5584 16822 5636
rect 17862 5624 17868 5636
rect 17710 5596 17868 5624
rect 15654 5516 15660 5568
rect 15712 5556 15718 5568
rect 17788 5556 17816 5596
rect 17862 5584 17868 5596
rect 17920 5584 17926 5636
rect 15712 5528 17816 5556
rect 15712 5516 15718 5528
rect 1104 5466 28152 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 28152 5466
rect 1104 5392 28152 5414
rect 12158 5352 12164 5364
rect 11808 5324 12164 5352
rect 11808 5293 11836 5324
rect 12158 5312 12164 5324
rect 12216 5312 12222 5364
rect 13262 5312 13268 5364
rect 13320 5312 13326 5364
rect 11793 5287 11851 5293
rect 11793 5253 11805 5287
rect 11839 5253 11851 5287
rect 13078 5284 13084 5296
rect 13018 5256 13084 5284
rect 11793 5247 11851 5253
rect 13078 5244 13084 5256
rect 13136 5284 13142 5296
rect 15654 5284 15660 5296
rect 13136 5256 15660 5284
rect 13136 5244 13142 5256
rect 15654 5244 15660 5256
rect 15712 5244 15718 5296
rect 11514 5176 11520 5228
rect 11572 5176 11578 5228
rect 1104 4922 28152 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 28152 4922
rect 1104 4848 28152 4870
rect 1104 4378 28152 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 28152 4378
rect 1104 4304 28152 4326
rect 1104 3834 28152 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 28152 3834
rect 1104 3760 28152 3782
rect 1104 3290 28152 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 28152 3290
rect 1104 3216 28152 3238
rect 1104 2746 28152 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 28152 2746
rect 1104 2672 28152 2694
rect 6089 2635 6147 2641
rect 6089 2601 6101 2635
rect 6135 2632 6147 2635
rect 7558 2632 7564 2644
rect 6135 2604 7564 2632
rect 6135 2601 6147 2604
rect 6089 2595 6147 2601
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 8662 2592 8668 2644
rect 8720 2592 8726 2644
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5868 2400 5917 2428
rect 5868 2388 5874 2400
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 8481 2431 8539 2437
rect 8481 2428 8493 2431
rect 8444 2400 8493 2428
rect 8444 2388 8450 2400
rect 8481 2397 8493 2400
rect 8527 2397 8539 2431
rect 8481 2391 8539 2397
rect 1104 2202 28152 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 28152 2202
rect 1104 2128 28152 2150
<< via1 >>
rect 16764 28908 16816 28960
rect 17500 28908 17552 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 12900 28704 12952 28756
rect 13544 28747 13596 28756
rect 13544 28713 13553 28747
rect 13553 28713 13587 28747
rect 13587 28713 13596 28747
rect 13544 28704 13596 28713
rect 14372 28747 14424 28756
rect 14372 28713 14381 28747
rect 14381 28713 14415 28747
rect 14415 28713 14424 28747
rect 14372 28704 14424 28713
rect 14832 28704 14884 28756
rect 15660 28747 15712 28756
rect 15660 28713 15669 28747
rect 15669 28713 15703 28747
rect 15703 28713 15712 28747
rect 15660 28704 15712 28713
rect 16120 28704 16172 28756
rect 17408 28704 17460 28756
rect 18052 28704 18104 28756
rect 19340 28704 19392 28756
rect 20628 28704 20680 28756
rect 21916 28704 21968 28756
rect 17224 28636 17276 28688
rect 17132 28500 17184 28552
rect 17500 28679 17552 28688
rect 17500 28645 17509 28679
rect 17509 28645 17543 28679
rect 17543 28645 17552 28679
rect 17500 28636 17552 28645
rect 18696 28636 18748 28688
rect 19984 28636 20036 28688
rect 21272 28636 21324 28688
rect 22560 28704 22612 28756
rect 23204 28704 23256 28756
rect 23848 28704 23900 28756
rect 25136 28704 25188 28756
rect 25780 28704 25832 28756
rect 26424 28704 26476 28756
rect 24492 28636 24544 28688
rect 26056 28500 26108 28552
rect 13268 28475 13320 28484
rect 13268 28441 13277 28475
rect 13277 28441 13311 28475
rect 13311 28441 13320 28475
rect 13268 28432 13320 28441
rect 14648 28475 14700 28484
rect 14648 28441 14657 28475
rect 14657 28441 14691 28475
rect 14691 28441 14700 28475
rect 14648 28432 14700 28441
rect 16856 28432 16908 28484
rect 17776 28364 17828 28416
rect 18144 28475 18196 28484
rect 18144 28441 18153 28475
rect 18153 28441 18187 28475
rect 18187 28441 18196 28475
rect 18144 28432 18196 28441
rect 18420 28475 18472 28484
rect 18420 28441 18429 28475
rect 18429 28441 18463 28475
rect 18463 28441 18472 28475
rect 18420 28432 18472 28441
rect 19340 28475 19392 28484
rect 19340 28441 19349 28475
rect 19349 28441 19383 28475
rect 19383 28441 19392 28475
rect 19340 28432 19392 28441
rect 20076 28432 20128 28484
rect 20444 28475 20496 28484
rect 20444 28441 20453 28475
rect 20453 28441 20487 28475
rect 20487 28441 20496 28475
rect 20444 28432 20496 28441
rect 20996 28475 21048 28484
rect 20996 28441 21005 28475
rect 21005 28441 21039 28475
rect 21039 28441 21048 28475
rect 20996 28432 21048 28441
rect 21456 28432 21508 28484
rect 22468 28475 22520 28484
rect 22468 28441 22477 28475
rect 22477 28441 22511 28475
rect 22511 28441 22520 28475
rect 22468 28432 22520 28441
rect 23020 28475 23072 28484
rect 23020 28441 23029 28475
rect 23029 28441 23063 28475
rect 23063 28441 23072 28475
rect 23020 28432 23072 28441
rect 23112 28432 23164 28484
rect 24492 28475 24544 28484
rect 24492 28441 24501 28475
rect 24501 28441 24535 28475
rect 24535 28441 24544 28475
rect 24492 28432 24544 28441
rect 25044 28475 25096 28484
rect 25044 28441 25053 28475
rect 25053 28441 25087 28475
rect 25087 28441 25096 28475
rect 25044 28432 25096 28441
rect 25596 28475 25648 28484
rect 25596 28441 25605 28475
rect 25605 28441 25639 28475
rect 25639 28441 25648 28475
rect 25596 28432 25648 28441
rect 26424 28475 26476 28484
rect 26424 28441 26433 28475
rect 26433 28441 26467 28475
rect 26467 28441 26476 28475
rect 26424 28432 26476 28441
rect 22008 28364 22060 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 18420 28160 18472 28212
rect 10140 28092 10192 28144
rect 6368 28024 6420 28076
rect 6920 28024 6972 28076
rect 10968 28067 11020 28076
rect 10968 28033 10977 28067
rect 10977 28033 11011 28067
rect 11011 28033 11020 28067
rect 10968 28024 11020 28033
rect 11796 28067 11848 28076
rect 9404 27956 9456 28008
rect 11796 28033 11804 28067
rect 11804 28033 11838 28067
rect 11838 28033 11848 28067
rect 11796 28024 11848 28033
rect 13268 28092 13320 28144
rect 19984 28160 20036 28212
rect 20076 28203 20128 28212
rect 20076 28169 20085 28203
rect 20085 28169 20119 28203
rect 20119 28169 20128 28203
rect 20076 28160 20128 28169
rect 20444 28160 20496 28212
rect 23020 28160 23072 28212
rect 27068 28160 27120 28212
rect 12256 28024 12308 28076
rect 17960 28067 18012 28076
rect 17960 28033 17969 28067
rect 17969 28033 18003 28067
rect 18003 28033 18012 28067
rect 17960 28024 18012 28033
rect 12072 27956 12124 28008
rect 17592 27956 17644 28008
rect 19156 27956 19208 28008
rect 19432 28135 19484 28144
rect 19432 28101 19441 28135
rect 19441 28101 19475 28135
rect 19475 28101 19484 28135
rect 19432 28092 19484 28101
rect 19616 28092 19668 28144
rect 19708 28067 19760 28076
rect 19708 28033 19717 28067
rect 19717 28033 19751 28067
rect 19751 28033 19760 28067
rect 19708 28024 19760 28033
rect 19800 28067 19852 28076
rect 19800 28033 19809 28067
rect 19809 28033 19843 28067
rect 19843 28033 19852 28067
rect 19800 28024 19852 28033
rect 20904 28092 20956 28144
rect 21916 28092 21968 28144
rect 21180 28067 21232 28076
rect 21180 28033 21189 28067
rect 21189 28033 21223 28067
rect 21223 28033 21232 28067
rect 21180 28024 21232 28033
rect 19064 27888 19116 27940
rect 19432 27888 19484 27940
rect 6460 27820 6512 27872
rect 7012 27863 7064 27872
rect 7012 27829 7021 27863
rect 7021 27829 7055 27863
rect 7055 27829 7064 27863
rect 7012 27820 7064 27829
rect 10232 27820 10284 27872
rect 10876 27820 10928 27872
rect 11704 27863 11756 27872
rect 11704 27829 11713 27863
rect 11713 27829 11747 27863
rect 11747 27829 11756 27863
rect 11704 27820 11756 27829
rect 19616 27820 19668 27872
rect 19984 27956 20036 28008
rect 22376 28024 22428 28076
rect 24584 28024 24636 28076
rect 24768 28024 24820 28076
rect 25780 28024 25832 28076
rect 24400 27956 24452 28008
rect 25228 27956 25280 28008
rect 19892 27888 19944 27940
rect 20628 27888 20680 27940
rect 25136 27888 25188 27940
rect 26332 28024 26384 28076
rect 29000 28024 29052 28076
rect 26148 27888 26200 27940
rect 24860 27863 24912 27872
rect 24860 27829 24869 27863
rect 24869 27829 24903 27863
rect 24903 27829 24912 27863
rect 24860 27820 24912 27829
rect 25320 27863 25372 27872
rect 25320 27829 25329 27863
rect 25329 27829 25363 27863
rect 25363 27829 25372 27863
rect 25320 27820 25372 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 2228 27480 2280 27532
rect 5264 27480 5316 27532
rect 5448 27548 5500 27600
rect 6368 27616 6420 27668
rect 6920 27548 6972 27600
rect 10876 27616 10928 27668
rect 11244 27616 11296 27668
rect 11796 27616 11848 27668
rect 3884 27412 3936 27464
rect 3976 27455 4028 27464
rect 3976 27421 3985 27455
rect 3985 27421 4019 27455
rect 4019 27421 4028 27455
rect 3976 27412 4028 27421
rect 4804 27412 4856 27464
rect 3700 27344 3752 27396
rect 6184 27412 6236 27464
rect 6460 27455 6512 27464
rect 6460 27421 6469 27455
rect 6469 27421 6503 27455
rect 6503 27421 6512 27455
rect 6460 27412 6512 27421
rect 6552 27412 6604 27464
rect 4068 27276 4120 27328
rect 4712 27276 4764 27328
rect 6000 27344 6052 27396
rect 5540 27276 5592 27328
rect 5816 27319 5868 27328
rect 5816 27285 5825 27319
rect 5825 27285 5859 27319
rect 5859 27285 5868 27319
rect 5816 27276 5868 27285
rect 6092 27319 6144 27328
rect 6092 27285 6101 27319
rect 6101 27285 6135 27319
rect 6135 27285 6144 27319
rect 6092 27276 6144 27285
rect 6460 27276 6512 27328
rect 7380 27276 7432 27328
rect 10140 27548 10192 27600
rect 10324 27591 10376 27600
rect 10324 27557 10333 27591
rect 10333 27557 10367 27591
rect 10367 27557 10376 27591
rect 10324 27548 10376 27557
rect 17224 27659 17276 27668
rect 17224 27625 17233 27659
rect 17233 27625 17267 27659
rect 17267 27625 17276 27659
rect 17224 27616 17276 27625
rect 18144 27616 18196 27668
rect 19064 27616 19116 27668
rect 7932 27412 7984 27464
rect 9404 27412 9456 27464
rect 10784 27523 10836 27532
rect 10784 27489 10793 27523
rect 10793 27489 10827 27523
rect 10827 27489 10836 27523
rect 10784 27480 10836 27489
rect 8300 27276 8352 27328
rect 9312 27276 9364 27328
rect 9496 27344 9548 27396
rect 10232 27412 10284 27464
rect 11336 27455 11388 27464
rect 11336 27421 11345 27455
rect 11345 27421 11379 27455
rect 11379 27421 11388 27455
rect 11336 27412 11388 27421
rect 11704 27412 11756 27464
rect 11796 27455 11848 27464
rect 11796 27421 11805 27455
rect 11805 27421 11839 27455
rect 11839 27421 11848 27455
rect 11796 27412 11848 27421
rect 12164 27412 12216 27464
rect 12256 27455 12308 27464
rect 17132 27548 17184 27600
rect 17776 27591 17828 27600
rect 17776 27557 17785 27591
rect 17785 27557 17819 27591
rect 17819 27557 17828 27591
rect 17776 27548 17828 27557
rect 12256 27421 12295 27455
rect 12295 27421 12308 27455
rect 12256 27412 12308 27421
rect 11888 27276 11940 27328
rect 11980 27276 12032 27328
rect 12808 27344 12860 27396
rect 17592 27412 17644 27464
rect 17868 27412 17920 27464
rect 18052 27455 18104 27464
rect 18052 27421 18061 27455
rect 18061 27421 18095 27455
rect 18095 27421 18104 27455
rect 18052 27412 18104 27421
rect 12992 27276 13044 27328
rect 18236 27276 18288 27328
rect 19432 27659 19484 27668
rect 19432 27625 19441 27659
rect 19441 27625 19475 27659
rect 19475 27625 19484 27659
rect 19432 27616 19484 27625
rect 20996 27616 21048 27668
rect 19524 27523 19576 27532
rect 19524 27489 19533 27523
rect 19533 27489 19567 27523
rect 19567 27489 19576 27523
rect 19524 27480 19576 27489
rect 19892 27548 19944 27600
rect 19984 27591 20036 27600
rect 19984 27557 19993 27591
rect 19993 27557 20027 27591
rect 20027 27557 20036 27591
rect 19984 27548 20036 27557
rect 20076 27548 20128 27600
rect 19800 27480 19852 27532
rect 20168 27480 20220 27532
rect 20352 27412 20404 27464
rect 21456 27591 21508 27600
rect 21456 27557 21465 27591
rect 21465 27557 21499 27591
rect 21499 27557 21508 27591
rect 21456 27548 21508 27557
rect 22468 27616 22520 27668
rect 24492 27616 24544 27668
rect 24584 27616 24636 27668
rect 24952 27616 25004 27668
rect 25136 27659 25188 27668
rect 25136 27625 25145 27659
rect 25145 27625 25179 27659
rect 25179 27625 25188 27659
rect 25136 27616 25188 27625
rect 25504 27616 25556 27668
rect 26424 27616 26476 27668
rect 19524 27344 19576 27396
rect 19800 27344 19852 27396
rect 20076 27344 20128 27396
rect 19432 27276 19484 27328
rect 20168 27319 20220 27328
rect 20168 27285 20177 27319
rect 20177 27285 20211 27319
rect 20211 27285 20220 27319
rect 20168 27276 20220 27285
rect 20260 27276 20312 27328
rect 20536 27387 20588 27396
rect 20536 27353 20545 27387
rect 20545 27353 20579 27387
rect 20579 27353 20588 27387
rect 20536 27344 20588 27353
rect 21640 27412 21692 27464
rect 22560 27412 22612 27464
rect 23112 27548 23164 27600
rect 25044 27548 25096 27600
rect 27712 27591 27764 27600
rect 27712 27557 27721 27591
rect 27721 27557 27755 27591
rect 27755 27557 27764 27591
rect 27712 27548 27764 27557
rect 21180 27344 21232 27396
rect 21916 27387 21968 27396
rect 21916 27353 21925 27387
rect 21925 27353 21959 27387
rect 21959 27353 21968 27387
rect 21916 27344 21968 27353
rect 22652 27319 22704 27328
rect 22652 27285 22661 27319
rect 22661 27285 22695 27319
rect 22695 27285 22704 27319
rect 22652 27276 22704 27285
rect 23020 27344 23072 27396
rect 23296 27455 23348 27464
rect 23296 27421 23305 27455
rect 23305 27421 23339 27455
rect 23339 27421 23348 27455
rect 23296 27412 23348 27421
rect 24032 27455 24084 27464
rect 24032 27421 24041 27455
rect 24041 27421 24075 27455
rect 24075 27421 24084 27455
rect 24032 27412 24084 27421
rect 24860 27480 24912 27532
rect 24492 27455 24544 27464
rect 24492 27421 24501 27455
rect 24501 27421 24535 27455
rect 24535 27421 24544 27455
rect 24492 27412 24544 27421
rect 23388 27344 23440 27396
rect 24308 27344 24360 27396
rect 24768 27412 24820 27464
rect 25044 27412 25096 27464
rect 25412 27455 25464 27464
rect 25412 27421 25421 27455
rect 25421 27421 25455 27455
rect 25455 27421 25464 27455
rect 25412 27412 25464 27421
rect 26148 27480 26200 27532
rect 26240 27455 26292 27464
rect 26240 27421 26249 27455
rect 26249 27421 26283 27455
rect 26283 27421 26292 27455
rect 26240 27412 26292 27421
rect 25872 27344 25924 27396
rect 24952 27276 25004 27328
rect 25136 27276 25188 27328
rect 25964 27319 26016 27328
rect 25964 27285 25973 27319
rect 25973 27285 26007 27319
rect 26007 27285 26016 27319
rect 25964 27276 26016 27285
rect 28356 27344 28408 27396
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 3976 27072 4028 27124
rect 5264 27115 5316 27124
rect 5264 27081 5273 27115
rect 5273 27081 5307 27115
rect 5307 27081 5316 27115
rect 5264 27072 5316 27081
rect 3148 27047 3200 27056
rect 3148 27013 3157 27047
rect 3157 27013 3191 27047
rect 3191 27013 3200 27047
rect 3148 27004 3200 27013
rect 2228 26936 2280 26988
rect 5724 27072 5776 27124
rect 1860 26868 1912 26920
rect 2320 26911 2372 26920
rect 2320 26877 2329 26911
rect 2329 26877 2363 26911
rect 2363 26877 2372 26911
rect 2320 26868 2372 26877
rect 2872 26732 2924 26784
rect 3700 26979 3752 26988
rect 3700 26945 3709 26979
rect 3709 26945 3743 26979
rect 3743 26945 3752 26979
rect 3700 26936 3752 26945
rect 4068 26979 4120 26988
rect 4068 26945 4077 26979
rect 4077 26945 4111 26979
rect 4111 26945 4120 26979
rect 4068 26936 4120 26945
rect 4620 26936 4672 26988
rect 5632 27004 5684 27056
rect 5816 27004 5868 27056
rect 6000 26936 6052 26988
rect 6552 26979 6604 26988
rect 6552 26945 6561 26979
rect 6561 26945 6595 26979
rect 6595 26945 6604 26979
rect 6552 26936 6604 26945
rect 6920 27072 6972 27124
rect 6736 26936 6788 26988
rect 7380 26979 7432 26988
rect 7380 26945 7389 26979
rect 7389 26945 7423 26979
rect 7423 26945 7432 26979
rect 7380 26936 7432 26945
rect 5264 26868 5316 26920
rect 4804 26800 4856 26852
rect 5724 26911 5776 26920
rect 5724 26877 5733 26911
rect 5733 26877 5767 26911
rect 5767 26877 5776 26911
rect 5724 26868 5776 26877
rect 3884 26775 3936 26784
rect 3884 26741 3893 26775
rect 3893 26741 3927 26775
rect 3927 26741 3936 26775
rect 3884 26732 3936 26741
rect 5724 26732 5776 26784
rect 6092 26868 6144 26920
rect 6368 26911 6420 26920
rect 6368 26877 6377 26911
rect 6377 26877 6411 26911
rect 6411 26877 6420 26911
rect 6368 26868 6420 26877
rect 7012 26868 7064 26920
rect 7932 26936 7984 26988
rect 10968 27072 11020 27124
rect 12072 27072 12124 27124
rect 16856 27072 16908 27124
rect 19340 27072 19392 27124
rect 19616 27072 19668 27124
rect 20168 27072 20220 27124
rect 8300 27004 8352 27056
rect 9128 26936 9180 26988
rect 10600 26936 10652 26988
rect 10232 26911 10284 26920
rect 10232 26877 10241 26911
rect 10241 26877 10275 26911
rect 10275 26877 10284 26911
rect 10232 26868 10284 26877
rect 6552 26800 6604 26852
rect 6000 26775 6052 26784
rect 6000 26741 6009 26775
rect 6009 26741 6043 26775
rect 6043 26741 6052 26775
rect 6000 26732 6052 26741
rect 6920 26732 6972 26784
rect 8208 26732 8260 26784
rect 10692 26732 10744 26784
rect 11336 27004 11388 27056
rect 11244 26979 11296 26988
rect 11244 26945 11253 26979
rect 11253 26945 11287 26979
rect 11287 26945 11296 26979
rect 11244 26936 11296 26945
rect 11704 26979 11756 26988
rect 11704 26945 11713 26979
rect 11713 26945 11747 26979
rect 11747 26945 11756 26979
rect 11704 26936 11756 26945
rect 11888 26936 11940 26988
rect 12532 27047 12584 27056
rect 12532 27013 12541 27047
rect 12541 27013 12575 27047
rect 12575 27013 12584 27047
rect 12532 27004 12584 27013
rect 12164 26936 12216 26988
rect 18972 27004 19024 27056
rect 19800 27004 19852 27056
rect 22008 27115 22060 27124
rect 22008 27081 22017 27115
rect 22017 27081 22051 27115
rect 22051 27081 22060 27115
rect 22008 27072 22060 27081
rect 18052 26936 18104 26988
rect 18236 26979 18288 26988
rect 18236 26945 18245 26979
rect 18245 26945 18279 26979
rect 18279 26945 18288 26979
rect 18236 26936 18288 26945
rect 19156 26979 19208 26988
rect 19156 26945 19164 26979
rect 19164 26945 19198 26979
rect 19198 26945 19208 26979
rect 19156 26936 19208 26945
rect 19248 26979 19300 26988
rect 19248 26945 19257 26979
rect 19257 26945 19291 26979
rect 19291 26945 19300 26979
rect 19248 26936 19300 26945
rect 19524 26979 19576 26988
rect 19524 26945 19533 26979
rect 19533 26945 19567 26979
rect 19567 26945 19576 26979
rect 19524 26936 19576 26945
rect 20168 26936 20220 26988
rect 11336 26800 11388 26852
rect 12440 26800 12492 26852
rect 19340 26868 19392 26920
rect 11980 26775 12032 26784
rect 11980 26741 11989 26775
rect 11989 26741 12023 26775
rect 12023 26741 12032 26775
rect 11980 26732 12032 26741
rect 12256 26732 12308 26784
rect 13084 26732 13136 26784
rect 19432 26732 19484 26784
rect 19800 26732 19852 26784
rect 20076 26843 20128 26852
rect 20076 26809 20085 26843
rect 20085 26809 20119 26843
rect 20119 26809 20128 26843
rect 20076 26800 20128 26809
rect 20444 26936 20496 26988
rect 23296 27072 23348 27124
rect 24860 27115 24912 27124
rect 24860 27081 24869 27115
rect 24869 27081 24903 27115
rect 24903 27081 24912 27115
rect 24860 27072 24912 27081
rect 25596 27072 25648 27124
rect 25872 27072 25924 27124
rect 26056 27115 26108 27124
rect 26056 27081 26065 27115
rect 26065 27081 26099 27115
rect 26099 27081 26108 27115
rect 26056 27072 26108 27081
rect 22836 27004 22888 27056
rect 23020 27004 23072 27056
rect 23112 27047 23164 27056
rect 23112 27013 23153 27047
rect 23153 27013 23164 27047
rect 23112 27004 23164 27013
rect 24492 27004 24544 27056
rect 26240 27072 26292 27124
rect 26332 27115 26384 27124
rect 26332 27081 26341 27115
rect 26341 27081 26375 27115
rect 26375 27081 26384 27115
rect 26332 27072 26384 27081
rect 20996 26979 21048 26988
rect 20996 26945 21005 26979
rect 21005 26945 21039 26979
rect 21039 26945 21048 26979
rect 20996 26936 21048 26945
rect 21640 26979 21692 26988
rect 21640 26945 21649 26979
rect 21649 26945 21683 26979
rect 21683 26945 21692 26979
rect 21640 26936 21692 26945
rect 22192 26936 22244 26988
rect 20352 26800 20404 26852
rect 20996 26800 21048 26852
rect 22284 26911 22336 26920
rect 22284 26877 22293 26911
rect 22293 26877 22327 26911
rect 22327 26877 22336 26911
rect 22284 26868 22336 26877
rect 24216 26979 24268 26988
rect 24216 26945 24225 26979
rect 24225 26945 24259 26979
rect 24259 26945 24268 26979
rect 24216 26936 24268 26945
rect 24400 26936 24452 26988
rect 24676 26979 24728 26988
rect 24676 26945 24685 26979
rect 24685 26945 24719 26979
rect 24719 26945 24728 26979
rect 24676 26936 24728 26945
rect 22652 26800 22704 26852
rect 24492 26911 24544 26920
rect 24492 26877 24501 26911
rect 24501 26877 24535 26911
rect 24535 26877 24544 26911
rect 24492 26868 24544 26877
rect 24952 26979 25004 26988
rect 24952 26945 24961 26979
rect 24961 26945 24995 26979
rect 24995 26945 25004 26979
rect 24952 26936 25004 26945
rect 25320 26936 25372 26988
rect 25780 26936 25832 26988
rect 25504 26868 25556 26920
rect 24032 26800 24084 26852
rect 25964 26979 26016 26988
rect 25964 26945 25973 26979
rect 25973 26945 26007 26979
rect 26007 26945 26016 26979
rect 25964 26936 26016 26945
rect 26516 26936 26568 26988
rect 26792 26800 26844 26852
rect 23112 26775 23164 26784
rect 23112 26741 23121 26775
rect 23121 26741 23155 26775
rect 23155 26741 23164 26775
rect 23112 26732 23164 26741
rect 23388 26732 23440 26784
rect 24308 26775 24360 26784
rect 24308 26741 24317 26775
rect 24317 26741 24351 26775
rect 24351 26741 24360 26775
rect 24308 26732 24360 26741
rect 24584 26732 24636 26784
rect 24676 26732 24728 26784
rect 27068 26732 27120 26784
rect 27712 26775 27764 26784
rect 27712 26741 27721 26775
rect 27721 26741 27755 26775
rect 27755 26741 27764 26775
rect 27712 26732 27764 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 2320 26528 2372 26580
rect 3148 26528 3200 26580
rect 3700 26528 3752 26580
rect 3976 26571 4028 26580
rect 3976 26537 3985 26571
rect 3985 26537 4019 26571
rect 4019 26537 4028 26571
rect 3976 26528 4028 26537
rect 4804 26528 4856 26580
rect 5172 26528 5224 26580
rect 6184 26528 6236 26580
rect 6920 26571 6972 26580
rect 6920 26537 6929 26571
rect 6929 26537 6963 26571
rect 6963 26537 6972 26571
rect 6920 26528 6972 26537
rect 9864 26528 9916 26580
rect 12532 26528 12584 26580
rect 17960 26528 18012 26580
rect 20168 26571 20220 26580
rect 20168 26537 20177 26571
rect 20177 26537 20211 26571
rect 20211 26537 20220 26571
rect 20168 26528 20220 26537
rect 20352 26571 20404 26580
rect 20352 26537 20361 26571
rect 20361 26537 20395 26571
rect 20395 26537 20404 26571
rect 20352 26528 20404 26537
rect 20996 26528 21048 26580
rect 22376 26571 22428 26580
rect 22376 26537 22385 26571
rect 22385 26537 22419 26571
rect 22419 26537 22428 26571
rect 22376 26528 22428 26537
rect 22928 26528 22980 26580
rect 24676 26528 24728 26580
rect 26792 26571 26844 26580
rect 26792 26537 26801 26571
rect 26801 26537 26835 26571
rect 26835 26537 26844 26571
rect 26792 26528 26844 26537
rect 4712 26460 4764 26512
rect 1860 26367 1912 26376
rect 1860 26333 1869 26367
rect 1869 26333 1903 26367
rect 1903 26333 1912 26367
rect 1860 26324 1912 26333
rect 1952 26324 2004 26376
rect 3056 26324 3108 26376
rect 3884 26324 3936 26376
rect 5080 26392 5132 26444
rect 2780 26256 2832 26308
rect 3424 26256 3476 26308
rect 5172 26367 5224 26376
rect 5172 26333 5181 26367
rect 5181 26333 5215 26367
rect 5215 26333 5224 26367
rect 5172 26324 5224 26333
rect 12624 26460 12676 26512
rect 23020 26460 23072 26512
rect 5540 26367 5592 26376
rect 5540 26333 5549 26367
rect 5549 26333 5583 26367
rect 5583 26333 5592 26367
rect 5540 26324 5592 26333
rect 5816 26367 5868 26376
rect 5816 26333 5825 26367
rect 5825 26333 5859 26367
rect 5859 26333 5868 26367
rect 5816 26324 5868 26333
rect 6460 26435 6512 26444
rect 6460 26401 6469 26435
rect 6469 26401 6503 26435
rect 6503 26401 6512 26435
rect 6460 26392 6512 26401
rect 6552 26392 6604 26444
rect 4620 26256 4672 26308
rect 6092 26299 6144 26308
rect 6092 26265 6101 26299
rect 6101 26265 6135 26299
rect 6135 26265 6144 26299
rect 6092 26256 6144 26265
rect 6736 26324 6788 26376
rect 6828 26188 6880 26240
rect 8852 26188 8904 26240
rect 9128 26367 9180 26376
rect 9128 26333 9137 26367
rect 9137 26333 9171 26367
rect 9171 26333 9180 26367
rect 9128 26324 9180 26333
rect 9312 26367 9364 26376
rect 9312 26333 9321 26367
rect 9321 26333 9355 26367
rect 9355 26333 9364 26367
rect 9312 26324 9364 26333
rect 10600 26367 10652 26376
rect 10600 26333 10609 26367
rect 10609 26333 10643 26367
rect 10643 26333 10652 26367
rect 10600 26324 10652 26333
rect 11244 26392 11296 26444
rect 11336 26324 11388 26376
rect 11980 26367 12032 26376
rect 11980 26333 11989 26367
rect 11989 26333 12023 26367
rect 12023 26333 12032 26367
rect 11980 26324 12032 26333
rect 12532 26367 12584 26376
rect 12532 26333 12541 26367
rect 12541 26333 12575 26367
rect 12575 26333 12584 26367
rect 12532 26324 12584 26333
rect 12992 26324 13044 26376
rect 13084 26367 13136 26376
rect 13084 26333 13093 26367
rect 13093 26333 13127 26367
rect 13127 26333 13136 26367
rect 13084 26324 13136 26333
rect 13176 26367 13228 26376
rect 13176 26333 13185 26367
rect 13185 26333 13219 26367
rect 13219 26333 13228 26367
rect 13176 26324 13228 26333
rect 20444 26392 20496 26444
rect 21640 26392 21692 26444
rect 23572 26503 23624 26512
rect 23572 26469 23581 26503
rect 23581 26469 23615 26503
rect 23615 26469 23624 26503
rect 23572 26460 23624 26469
rect 27528 26460 27580 26512
rect 23296 26435 23348 26444
rect 23296 26401 23305 26435
rect 23305 26401 23339 26435
rect 23339 26401 23348 26435
rect 23296 26392 23348 26401
rect 25044 26392 25096 26444
rect 25412 26392 25464 26444
rect 26240 26392 26292 26444
rect 19800 26324 19852 26376
rect 9772 26231 9824 26240
rect 9772 26197 9781 26231
rect 9781 26197 9815 26231
rect 9815 26197 9824 26231
rect 9772 26188 9824 26197
rect 10876 26231 10928 26240
rect 10876 26197 10885 26231
rect 10885 26197 10919 26231
rect 10919 26197 10928 26231
rect 10876 26188 10928 26197
rect 12716 26256 12768 26308
rect 22468 26367 22520 26376
rect 22468 26333 22477 26367
rect 22477 26333 22511 26367
rect 22511 26333 22520 26367
rect 22468 26324 22520 26333
rect 22652 26367 22704 26376
rect 22652 26333 22661 26367
rect 22661 26333 22695 26367
rect 22695 26333 22704 26367
rect 22652 26324 22704 26333
rect 22744 26324 22796 26376
rect 22928 26367 22980 26376
rect 22928 26333 22937 26367
rect 22937 26333 22971 26367
rect 22971 26333 22980 26367
rect 22928 26324 22980 26333
rect 24308 26324 24360 26376
rect 25136 26367 25188 26376
rect 25136 26333 25145 26367
rect 25145 26333 25179 26367
rect 25179 26333 25188 26367
rect 25136 26324 25188 26333
rect 22284 26256 22336 26308
rect 23112 26256 23164 26308
rect 12440 26188 12492 26240
rect 20168 26188 20220 26240
rect 20444 26188 20496 26240
rect 24400 26256 24452 26308
rect 24492 26256 24544 26308
rect 25228 26256 25280 26308
rect 25596 26324 25648 26376
rect 26332 26367 26384 26376
rect 26332 26333 26341 26367
rect 26341 26333 26375 26367
rect 26375 26333 26384 26367
rect 26332 26324 26384 26333
rect 26792 26324 26844 26376
rect 26424 26256 26476 26308
rect 25412 26231 25464 26240
rect 25412 26197 25421 26231
rect 25421 26197 25455 26231
rect 25455 26197 25464 26231
rect 25412 26188 25464 26197
rect 25688 26188 25740 26240
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 5448 25916 5500 25968
rect 2780 25891 2832 25900
rect 2780 25857 2789 25891
rect 2789 25857 2823 25891
rect 2823 25857 2832 25891
rect 2780 25848 2832 25857
rect 3148 25891 3200 25900
rect 3148 25857 3157 25891
rect 3157 25857 3191 25891
rect 3191 25857 3200 25891
rect 3148 25848 3200 25857
rect 6000 25848 6052 25900
rect 8208 25959 8260 25968
rect 8208 25925 8217 25959
rect 8217 25925 8251 25959
rect 8251 25925 8260 25959
rect 8208 25916 8260 25925
rect 12256 25984 12308 26036
rect 12440 26027 12492 26036
rect 12440 25993 12449 26027
rect 12449 25993 12483 26027
rect 12483 25993 12492 26027
rect 12440 25984 12492 25993
rect 13176 25984 13228 26036
rect 25412 25984 25464 26036
rect 26516 25984 26568 26036
rect 12808 25959 12860 25968
rect 12808 25925 12817 25959
rect 12817 25925 12851 25959
rect 12851 25925 12860 25959
rect 12808 25916 12860 25925
rect 22468 25916 22520 25968
rect 23020 25959 23072 25968
rect 23020 25925 23029 25959
rect 23029 25925 23063 25959
rect 23063 25925 23072 25959
rect 23020 25916 23072 25925
rect 23388 25916 23440 25968
rect 25136 25916 25188 25968
rect 25596 25959 25648 25968
rect 25596 25925 25605 25959
rect 25605 25925 25639 25959
rect 25639 25925 25648 25959
rect 25596 25916 25648 25925
rect 2872 25780 2924 25832
rect 6828 25823 6880 25832
rect 6828 25789 6837 25823
rect 6837 25789 6871 25823
rect 6871 25789 6880 25823
rect 6828 25780 6880 25789
rect 8852 25891 8904 25900
rect 8852 25857 8861 25891
rect 8861 25857 8895 25891
rect 8895 25857 8904 25891
rect 8852 25848 8904 25857
rect 12716 25848 12768 25900
rect 12624 25780 12676 25832
rect 12808 25780 12860 25832
rect 20444 25891 20496 25900
rect 20444 25857 20453 25891
rect 20453 25857 20487 25891
rect 20487 25857 20496 25891
rect 20444 25848 20496 25857
rect 20904 25848 20956 25900
rect 22008 25848 22060 25900
rect 22652 25891 22704 25900
rect 22652 25857 22661 25891
rect 22661 25857 22695 25891
rect 22695 25857 22704 25891
rect 22652 25848 22704 25857
rect 24216 25848 24268 25900
rect 24860 25848 24912 25900
rect 25044 25848 25096 25900
rect 26332 25848 26384 25900
rect 26424 25891 26476 25900
rect 26424 25857 26433 25891
rect 26433 25857 26467 25891
rect 26467 25857 26476 25891
rect 26424 25848 26476 25857
rect 26792 25780 26844 25832
rect 25504 25712 25556 25764
rect 25596 25712 25648 25764
rect 7564 25644 7616 25696
rect 7656 25687 7708 25696
rect 7656 25653 7665 25687
rect 7665 25653 7699 25687
rect 7699 25653 7708 25687
rect 7656 25644 7708 25653
rect 8668 25644 8720 25696
rect 12072 25687 12124 25696
rect 12072 25653 12081 25687
rect 12081 25653 12115 25687
rect 12115 25653 12124 25687
rect 12072 25644 12124 25653
rect 20536 25687 20588 25696
rect 20536 25653 20545 25687
rect 20545 25653 20579 25687
rect 20579 25653 20588 25687
rect 20536 25644 20588 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 12440 25440 12492 25492
rect 12992 25483 13044 25492
rect 12992 25449 13001 25483
rect 13001 25449 13035 25483
rect 13035 25449 13044 25483
rect 12992 25440 13044 25449
rect 17408 25440 17460 25492
rect 23020 25440 23072 25492
rect 25872 25440 25924 25492
rect 26332 25440 26384 25492
rect 20536 25372 20588 25424
rect 26240 25372 26292 25424
rect 9772 25236 9824 25288
rect 9864 25279 9916 25288
rect 9864 25245 9873 25279
rect 9873 25245 9907 25279
rect 9907 25245 9916 25279
rect 9864 25236 9916 25245
rect 10692 25279 10744 25288
rect 10692 25245 10701 25279
rect 10701 25245 10735 25279
rect 10735 25245 10744 25279
rect 10692 25236 10744 25245
rect 10876 25279 10928 25288
rect 10876 25245 10885 25279
rect 10885 25245 10919 25279
rect 10919 25245 10928 25279
rect 10876 25236 10928 25245
rect 13176 25304 13228 25356
rect 12440 25279 12492 25288
rect 12440 25245 12449 25279
rect 12449 25245 12483 25279
rect 12483 25245 12492 25279
rect 12440 25236 12492 25245
rect 12624 25279 12676 25288
rect 12624 25245 12633 25279
rect 12633 25245 12667 25279
rect 12667 25245 12676 25279
rect 12624 25236 12676 25245
rect 12716 25279 12768 25288
rect 12716 25245 12725 25279
rect 12725 25245 12759 25279
rect 12759 25245 12768 25279
rect 12716 25236 12768 25245
rect 15568 25279 15620 25288
rect 15568 25245 15577 25279
rect 15577 25245 15611 25279
rect 15611 25245 15620 25279
rect 15568 25236 15620 25245
rect 15660 25279 15712 25288
rect 15660 25245 15669 25279
rect 15669 25245 15703 25279
rect 15703 25245 15712 25279
rect 15660 25236 15712 25245
rect 15936 25236 15988 25288
rect 22008 25279 22060 25288
rect 22008 25245 22017 25279
rect 22017 25245 22051 25279
rect 22051 25245 22060 25279
rect 22008 25236 22060 25245
rect 25320 25236 25372 25288
rect 11060 25168 11112 25220
rect 9864 25143 9916 25152
rect 9864 25109 9873 25143
rect 9873 25109 9907 25143
rect 9907 25109 9916 25143
rect 9864 25100 9916 25109
rect 10692 25100 10744 25152
rect 10968 25100 11020 25152
rect 11888 25100 11940 25152
rect 12440 25100 12492 25152
rect 16120 25168 16172 25220
rect 17592 25168 17644 25220
rect 22192 25211 22244 25220
rect 22192 25177 22201 25211
rect 22201 25177 22235 25211
rect 22235 25177 22244 25211
rect 22192 25168 22244 25177
rect 27528 25279 27580 25288
rect 27528 25245 27537 25279
rect 27537 25245 27571 25279
rect 27571 25245 27580 25279
rect 27528 25236 27580 25245
rect 26332 25211 26384 25220
rect 26332 25177 26341 25211
rect 26341 25177 26375 25211
rect 26375 25177 26384 25211
rect 26332 25168 26384 25177
rect 27436 25168 27488 25220
rect 16948 25143 17000 25152
rect 16948 25109 16973 25143
rect 16973 25109 17000 25143
rect 16948 25100 17000 25109
rect 17132 25143 17184 25152
rect 17132 25109 17141 25143
rect 17141 25109 17175 25143
rect 17175 25109 17184 25143
rect 17132 25100 17184 25109
rect 25596 25100 25648 25152
rect 27068 25143 27120 25152
rect 27068 25109 27077 25143
rect 27077 25109 27111 25143
rect 27111 25109 27120 25143
rect 27068 25100 27120 25109
rect 27712 25143 27764 25152
rect 27712 25109 27721 25143
rect 27721 25109 27755 25143
rect 27755 25109 27764 25143
rect 27712 25100 27764 25109
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 10876 24896 10928 24948
rect 10968 24896 11020 24948
rect 11060 24896 11112 24948
rect 2872 24828 2924 24880
rect 848 24760 900 24812
rect 2504 24803 2556 24812
rect 2504 24769 2513 24803
rect 2513 24769 2547 24803
rect 2547 24769 2556 24803
rect 2504 24760 2556 24769
rect 2688 24803 2740 24812
rect 2688 24769 2697 24803
rect 2697 24769 2731 24803
rect 2731 24769 2740 24803
rect 2688 24760 2740 24769
rect 4068 24760 4120 24812
rect 4896 24828 4948 24880
rect 9864 24828 9916 24880
rect 5080 24803 5132 24812
rect 5080 24769 5089 24803
rect 5089 24769 5123 24803
rect 5123 24769 5132 24803
rect 5080 24760 5132 24769
rect 5264 24803 5316 24812
rect 5264 24769 5273 24803
rect 5273 24769 5307 24803
rect 5307 24769 5316 24803
rect 5264 24760 5316 24769
rect 5356 24803 5408 24812
rect 5356 24769 5365 24803
rect 5365 24769 5399 24803
rect 5399 24769 5408 24803
rect 5356 24760 5408 24769
rect 5448 24803 5500 24812
rect 5448 24769 5457 24803
rect 5457 24769 5491 24803
rect 5491 24769 5500 24803
rect 5448 24760 5500 24769
rect 7656 24760 7708 24812
rect 4712 24692 4764 24744
rect 8392 24803 8444 24812
rect 8392 24769 8401 24803
rect 8401 24769 8435 24803
rect 8435 24769 8444 24803
rect 8392 24760 8444 24769
rect 8668 24803 8720 24812
rect 8668 24769 8677 24803
rect 8677 24769 8711 24803
rect 8711 24769 8720 24803
rect 8668 24760 8720 24769
rect 10692 24760 10744 24812
rect 10876 24803 10928 24812
rect 10876 24769 10885 24803
rect 10885 24769 10919 24803
rect 10919 24769 10928 24803
rect 10876 24760 10928 24769
rect 5908 24624 5960 24676
rect 8392 24624 8444 24676
rect 10968 24624 11020 24676
rect 2136 24556 2188 24608
rect 2964 24599 3016 24608
rect 2964 24565 2973 24599
rect 2973 24565 3007 24599
rect 3007 24565 3016 24599
rect 2964 24556 3016 24565
rect 4620 24556 4672 24608
rect 9312 24556 9364 24608
rect 9404 24599 9456 24608
rect 9404 24565 9413 24599
rect 9413 24565 9447 24599
rect 9447 24565 9456 24599
rect 9404 24556 9456 24565
rect 10416 24556 10468 24608
rect 12072 24828 12124 24880
rect 15660 24896 15712 24948
rect 15936 24828 15988 24880
rect 16856 24939 16908 24948
rect 16856 24905 16865 24939
rect 16865 24905 16899 24939
rect 16899 24905 16908 24939
rect 16856 24896 16908 24905
rect 17408 24939 17460 24948
rect 17408 24905 17417 24939
rect 17417 24905 17451 24939
rect 17451 24905 17460 24939
rect 17408 24896 17460 24905
rect 22008 24896 22060 24948
rect 26332 24896 26384 24948
rect 14832 24803 14884 24812
rect 14832 24769 14841 24803
rect 14841 24769 14875 24803
rect 14875 24769 14884 24803
rect 14832 24760 14884 24769
rect 11980 24692 12032 24744
rect 12348 24692 12400 24744
rect 12532 24692 12584 24744
rect 15568 24760 15620 24812
rect 15660 24760 15712 24812
rect 16120 24803 16172 24812
rect 16120 24769 16129 24803
rect 16129 24769 16163 24803
rect 16163 24769 16172 24803
rect 16120 24760 16172 24769
rect 19156 24828 19208 24880
rect 22192 24828 22244 24880
rect 15936 24692 15988 24744
rect 16120 24624 16172 24676
rect 16948 24692 17000 24744
rect 17592 24803 17644 24812
rect 17592 24769 17601 24803
rect 17601 24769 17635 24803
rect 17635 24769 17644 24803
rect 17592 24760 17644 24769
rect 19892 24760 19944 24812
rect 22008 24803 22060 24812
rect 22008 24769 22017 24803
rect 22017 24769 22051 24803
rect 22051 24769 22060 24803
rect 22008 24760 22060 24769
rect 23756 24828 23808 24880
rect 11704 24556 11756 24608
rect 12992 24556 13044 24608
rect 15844 24556 15896 24608
rect 18052 24624 18104 24676
rect 21456 24624 21508 24676
rect 22928 24803 22980 24812
rect 22928 24769 22937 24803
rect 22937 24769 22971 24803
rect 22971 24769 22980 24803
rect 22928 24760 22980 24769
rect 23112 24803 23164 24812
rect 23112 24769 23121 24803
rect 23121 24769 23155 24803
rect 23155 24769 23164 24803
rect 23112 24760 23164 24769
rect 17224 24556 17276 24608
rect 17868 24556 17920 24608
rect 21364 24556 21416 24608
rect 22192 24599 22244 24608
rect 22192 24565 22201 24599
rect 22201 24565 22235 24599
rect 22235 24565 22244 24599
rect 22192 24556 22244 24565
rect 22376 24599 22428 24608
rect 22376 24565 22385 24599
rect 22385 24565 22419 24599
rect 22419 24565 22428 24599
rect 22376 24556 22428 24565
rect 25228 24760 25280 24812
rect 25780 24803 25832 24812
rect 25780 24769 25789 24803
rect 25789 24769 25823 24803
rect 25823 24769 25832 24803
rect 25780 24760 25832 24769
rect 25872 24803 25924 24812
rect 25872 24769 25881 24803
rect 25881 24769 25915 24803
rect 25915 24769 25924 24803
rect 25872 24760 25924 24769
rect 26240 24828 26292 24880
rect 25044 24692 25096 24744
rect 25596 24735 25648 24744
rect 25596 24701 25605 24735
rect 25605 24701 25639 24735
rect 25639 24701 25648 24735
rect 25596 24692 25648 24701
rect 23480 24556 23532 24608
rect 25872 24556 25924 24608
rect 26884 24556 26936 24608
rect 27160 24599 27212 24608
rect 27160 24565 27169 24599
rect 27169 24565 27203 24599
rect 27203 24565 27212 24599
rect 27160 24556 27212 24565
rect 27712 24599 27764 24608
rect 27712 24565 27721 24599
rect 27721 24565 27755 24599
rect 27755 24565 27764 24599
rect 27712 24556 27764 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 2780 24352 2832 24404
rect 3424 24395 3476 24404
rect 3424 24361 3433 24395
rect 3433 24361 3467 24395
rect 3467 24361 3476 24395
rect 3424 24352 3476 24361
rect 8392 24352 8444 24404
rect 14832 24352 14884 24404
rect 2504 24191 2556 24200
rect 2504 24157 2513 24191
rect 2513 24157 2547 24191
rect 2547 24157 2556 24191
rect 2504 24148 2556 24157
rect 2596 24148 2648 24200
rect 4068 24284 4120 24336
rect 2964 24216 3016 24268
rect 4804 24216 4856 24268
rect 5080 24259 5132 24268
rect 5080 24225 5089 24259
rect 5089 24225 5123 24259
rect 5123 24225 5132 24259
rect 5080 24216 5132 24225
rect 10876 24284 10928 24336
rect 12716 24284 12768 24336
rect 14188 24284 14240 24336
rect 11704 24259 11756 24268
rect 11704 24225 11713 24259
rect 11713 24225 11747 24259
rect 11747 24225 11756 24259
rect 11704 24216 11756 24225
rect 848 24080 900 24132
rect 2136 24080 2188 24132
rect 4712 24148 4764 24200
rect 5264 24148 5316 24200
rect 7472 24191 7524 24200
rect 7472 24157 7481 24191
rect 7481 24157 7515 24191
rect 7515 24157 7524 24191
rect 7472 24148 7524 24157
rect 7564 24148 7616 24200
rect 9404 24191 9456 24200
rect 9404 24157 9413 24191
rect 9413 24157 9447 24191
rect 9447 24157 9456 24191
rect 9404 24148 9456 24157
rect 9864 24148 9916 24200
rect 9956 24191 10008 24200
rect 9956 24157 9965 24191
rect 9965 24157 9999 24191
rect 9999 24157 10008 24191
rect 9956 24148 10008 24157
rect 2228 24012 2280 24064
rect 3148 24012 3200 24064
rect 4436 24080 4488 24132
rect 4896 24080 4948 24132
rect 5632 24123 5684 24132
rect 5632 24089 5641 24123
rect 5641 24089 5675 24123
rect 5675 24089 5684 24123
rect 5632 24080 5684 24089
rect 9220 24123 9272 24132
rect 9220 24089 9229 24123
rect 9229 24089 9263 24123
rect 9263 24089 9272 24123
rect 10140 24148 10192 24200
rect 10876 24148 10928 24200
rect 11980 24191 12032 24200
rect 11980 24157 11989 24191
rect 11989 24157 12023 24191
rect 12023 24157 12032 24191
rect 11980 24148 12032 24157
rect 12072 24148 12124 24200
rect 15660 24352 15712 24404
rect 22008 24352 22060 24404
rect 23112 24352 23164 24404
rect 17040 24284 17092 24336
rect 17592 24284 17644 24336
rect 18052 24259 18104 24268
rect 18052 24225 18061 24259
rect 18061 24225 18095 24259
rect 18095 24225 18104 24259
rect 18052 24216 18104 24225
rect 18512 24216 18564 24268
rect 22376 24216 22428 24268
rect 23480 24395 23532 24404
rect 23480 24361 23489 24395
rect 23489 24361 23523 24395
rect 23523 24361 23532 24395
rect 23480 24352 23532 24361
rect 25872 24395 25924 24404
rect 25872 24361 25881 24395
rect 25881 24361 25915 24395
rect 25915 24361 25924 24395
rect 25872 24352 25924 24361
rect 27528 24352 27580 24404
rect 24676 24284 24728 24336
rect 25044 24216 25096 24268
rect 12992 24191 13044 24200
rect 12992 24157 13001 24191
rect 13001 24157 13035 24191
rect 13035 24157 13044 24191
rect 12992 24148 13044 24157
rect 14372 24148 14424 24200
rect 9220 24080 9272 24089
rect 10600 24080 10652 24132
rect 15660 24191 15712 24200
rect 15660 24157 15669 24191
rect 15669 24157 15703 24191
rect 15703 24157 15712 24191
rect 15660 24148 15712 24157
rect 15936 24123 15988 24132
rect 15936 24089 15945 24123
rect 15945 24089 15979 24123
rect 15979 24089 15988 24123
rect 15936 24080 15988 24089
rect 16396 24080 16448 24132
rect 21272 24191 21324 24200
rect 21272 24157 21281 24191
rect 21281 24157 21315 24191
rect 21315 24157 21324 24191
rect 21272 24148 21324 24157
rect 21456 24191 21508 24200
rect 21456 24157 21465 24191
rect 21465 24157 21499 24191
rect 21499 24157 21508 24191
rect 21456 24148 21508 24157
rect 21548 24191 21600 24200
rect 21548 24157 21557 24191
rect 21557 24157 21591 24191
rect 21591 24157 21600 24191
rect 21548 24148 21600 24157
rect 20352 24080 20404 24132
rect 12440 24012 12492 24064
rect 13544 24012 13596 24064
rect 17500 24012 17552 24064
rect 19064 24012 19116 24064
rect 20536 24080 20588 24132
rect 22008 24012 22060 24064
rect 22192 24012 22244 24064
rect 23756 24191 23808 24200
rect 23756 24157 23765 24191
rect 23765 24157 23799 24191
rect 23799 24157 23808 24191
rect 23756 24148 23808 24157
rect 24952 24148 25004 24200
rect 25136 24191 25188 24200
rect 25136 24157 25145 24191
rect 25145 24157 25179 24191
rect 25179 24157 25188 24191
rect 25136 24148 25188 24157
rect 26332 24284 26384 24336
rect 25596 24216 25648 24268
rect 25964 24216 26016 24268
rect 27160 24216 27212 24268
rect 26884 24191 26936 24200
rect 26884 24157 26893 24191
rect 26893 24157 26927 24191
rect 26927 24157 26936 24191
rect 26884 24148 26936 24157
rect 27068 24191 27120 24200
rect 27068 24157 27077 24191
rect 27077 24157 27111 24191
rect 27111 24157 27120 24191
rect 27068 24148 27120 24157
rect 27344 24148 27396 24200
rect 25872 24080 25924 24132
rect 24492 24055 24544 24064
rect 24492 24021 24501 24055
rect 24501 24021 24535 24055
rect 24535 24021 24544 24055
rect 24492 24012 24544 24021
rect 24768 24012 24820 24064
rect 24860 24055 24912 24064
rect 24860 24021 24869 24055
rect 24869 24021 24903 24055
rect 24903 24021 24912 24055
rect 24860 24012 24912 24021
rect 26056 24055 26108 24064
rect 26056 24021 26065 24055
rect 26065 24021 26099 24055
rect 26099 24021 26108 24055
rect 26056 24012 26108 24021
rect 27068 24012 27120 24064
rect 27712 24055 27764 24064
rect 27712 24021 27721 24055
rect 27721 24021 27755 24055
rect 27755 24021 27764 24055
rect 27712 24012 27764 24021
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 4804 23808 4856 23860
rect 2504 23783 2556 23792
rect 2504 23749 2513 23783
rect 2513 23749 2547 23783
rect 2547 23749 2556 23783
rect 2504 23740 2556 23749
rect 2596 23672 2648 23724
rect 4620 23740 4672 23792
rect 5632 23740 5684 23792
rect 4712 23715 4764 23724
rect 4712 23681 4721 23715
rect 4721 23681 4755 23715
rect 4755 23681 4764 23715
rect 4712 23672 4764 23681
rect 5908 23715 5960 23724
rect 5908 23681 5951 23715
rect 5951 23681 5960 23715
rect 9220 23851 9272 23860
rect 9220 23817 9229 23851
rect 9229 23817 9263 23851
rect 9263 23817 9272 23851
rect 9220 23808 9272 23817
rect 9404 23783 9456 23792
rect 9404 23749 9413 23783
rect 9413 23749 9447 23783
rect 9447 23749 9456 23783
rect 9404 23740 9456 23749
rect 10876 23740 10928 23792
rect 15660 23808 15712 23860
rect 18236 23808 18288 23860
rect 20536 23808 20588 23860
rect 21548 23808 21600 23860
rect 23480 23808 23532 23860
rect 5908 23672 5960 23681
rect 7472 23672 7524 23724
rect 9036 23672 9088 23724
rect 9312 23715 9364 23724
rect 9312 23681 9321 23715
rect 9321 23681 9355 23715
rect 9355 23681 9364 23715
rect 9312 23672 9364 23681
rect 10232 23715 10284 23724
rect 10232 23681 10241 23715
rect 10241 23681 10275 23715
rect 10275 23681 10284 23715
rect 10232 23672 10284 23681
rect 12716 23672 12768 23724
rect 12900 23715 12952 23724
rect 12900 23681 12909 23715
rect 12909 23681 12943 23715
rect 12943 23681 12952 23715
rect 12900 23672 12952 23681
rect 13544 23783 13596 23792
rect 13544 23749 13553 23783
rect 13553 23749 13587 23783
rect 13587 23749 13596 23783
rect 13544 23740 13596 23749
rect 1952 23647 2004 23656
rect 1952 23613 1961 23647
rect 1961 23613 1995 23647
rect 1995 23613 2004 23647
rect 1952 23604 2004 23613
rect 5264 23604 5316 23656
rect 2780 23536 2832 23588
rect 5540 23536 5592 23588
rect 7564 23604 7616 23656
rect 9864 23604 9916 23656
rect 12348 23604 12400 23656
rect 12808 23604 12860 23656
rect 13544 23604 13596 23656
rect 16396 23740 16448 23792
rect 17500 23783 17552 23792
rect 17500 23749 17509 23783
rect 17509 23749 17543 23783
rect 17543 23749 17552 23783
rect 17500 23740 17552 23749
rect 15844 23672 15896 23724
rect 16120 23715 16172 23724
rect 16120 23681 16129 23715
rect 16129 23681 16163 23715
rect 16163 23681 16172 23715
rect 16120 23672 16172 23681
rect 17040 23672 17092 23724
rect 17132 23715 17184 23724
rect 17132 23681 17141 23715
rect 17141 23681 17175 23715
rect 17175 23681 17184 23715
rect 17132 23672 17184 23681
rect 17224 23715 17276 23724
rect 17224 23681 17233 23715
rect 17233 23681 17267 23715
rect 17267 23681 17276 23715
rect 17224 23672 17276 23681
rect 18052 23672 18104 23724
rect 18604 23672 18656 23724
rect 17868 23647 17920 23656
rect 17868 23613 17877 23647
rect 17877 23613 17911 23647
rect 17911 23613 17920 23647
rect 19156 23783 19208 23792
rect 19156 23749 19165 23783
rect 19165 23749 19199 23783
rect 19199 23749 19208 23783
rect 19156 23740 19208 23749
rect 20352 23740 20404 23792
rect 21364 23783 21416 23792
rect 21364 23749 21373 23783
rect 21373 23749 21407 23783
rect 21407 23749 21416 23783
rect 21364 23740 21416 23749
rect 22008 23740 22060 23792
rect 18788 23715 18840 23724
rect 18788 23681 18797 23715
rect 18797 23681 18831 23715
rect 18831 23681 18840 23715
rect 18788 23672 18840 23681
rect 19064 23715 19116 23724
rect 19064 23681 19073 23715
rect 19073 23681 19107 23715
rect 19107 23681 19116 23715
rect 19064 23672 19116 23681
rect 17868 23604 17920 23613
rect 19892 23647 19944 23656
rect 19892 23613 19901 23647
rect 19901 23613 19935 23647
rect 19935 23613 19944 23647
rect 19892 23604 19944 23613
rect 21640 23647 21692 23656
rect 21640 23613 21649 23647
rect 21649 23613 21683 23647
rect 21683 23613 21692 23647
rect 21640 23604 21692 23613
rect 25504 23740 25556 23792
rect 25596 23715 25648 23724
rect 25596 23681 25605 23715
rect 25605 23681 25639 23715
rect 25639 23681 25648 23715
rect 25596 23672 25648 23681
rect 26148 23808 26200 23860
rect 26424 23808 26476 23860
rect 25872 23783 25924 23792
rect 25872 23749 25881 23783
rect 25881 23749 25915 23783
rect 25915 23749 25924 23783
rect 25872 23740 25924 23749
rect 25964 23783 26016 23792
rect 25964 23749 25973 23783
rect 25973 23749 26007 23783
rect 26007 23749 26016 23783
rect 25964 23740 26016 23749
rect 22560 23604 22612 23656
rect 23296 23647 23348 23656
rect 23296 23613 23305 23647
rect 23305 23613 23339 23647
rect 23339 23613 23348 23647
rect 23296 23604 23348 23613
rect 23572 23647 23624 23656
rect 23572 23613 23581 23647
rect 23581 23613 23615 23647
rect 23615 23613 23624 23647
rect 23572 23604 23624 23613
rect 24032 23647 24084 23656
rect 24032 23613 24041 23647
rect 24041 23613 24075 23647
rect 24075 23613 24084 23647
rect 24032 23604 24084 23613
rect 25044 23604 25096 23656
rect 25412 23604 25464 23656
rect 26056 23715 26108 23724
rect 26056 23681 26070 23715
rect 26070 23681 26104 23715
rect 26104 23681 26108 23715
rect 26056 23672 26108 23681
rect 26976 23672 27028 23724
rect 6920 23536 6972 23588
rect 8116 23536 8168 23588
rect 13176 23579 13228 23588
rect 13176 23545 13185 23579
rect 13185 23545 13219 23579
rect 13219 23545 13228 23579
rect 13176 23536 13228 23545
rect 16856 23579 16908 23588
rect 16856 23545 16865 23579
rect 16865 23545 16899 23579
rect 16899 23545 16908 23579
rect 16856 23536 16908 23545
rect 17408 23536 17460 23588
rect 18236 23536 18288 23588
rect 10508 23468 10560 23520
rect 15016 23511 15068 23520
rect 15016 23477 15025 23511
rect 15025 23477 15059 23511
rect 15059 23477 15068 23511
rect 15016 23468 15068 23477
rect 15752 23468 15804 23520
rect 17132 23468 17184 23520
rect 17960 23511 18012 23520
rect 17960 23477 17969 23511
rect 17969 23477 18003 23511
rect 18003 23477 18012 23511
rect 17960 23468 18012 23477
rect 18328 23511 18380 23520
rect 18328 23477 18337 23511
rect 18337 23477 18371 23511
rect 18371 23477 18380 23511
rect 18328 23468 18380 23477
rect 21916 23468 21968 23520
rect 27528 23468 27580 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 7840 23264 7892 23316
rect 9864 23264 9916 23316
rect 11980 23264 12032 23316
rect 12716 23264 12768 23316
rect 18052 23264 18104 23316
rect 848 23060 900 23112
rect 2688 23128 2740 23180
rect 2136 22992 2188 23044
rect 3148 23060 3200 23112
rect 2320 22967 2372 22976
rect 2320 22933 2329 22967
rect 2329 22933 2363 22967
rect 2363 22933 2372 22967
rect 2320 22924 2372 22933
rect 2688 22924 2740 22976
rect 2964 22924 3016 22976
rect 3792 22924 3844 22976
rect 4620 23128 4672 23180
rect 5540 23128 5592 23180
rect 9312 23128 9364 23180
rect 16856 23196 16908 23248
rect 18236 23196 18288 23248
rect 22284 23264 22336 23316
rect 4252 22992 4304 23044
rect 4620 22992 4672 23044
rect 5632 23060 5684 23112
rect 6092 23060 6144 23112
rect 6920 23060 6972 23112
rect 6276 23035 6328 23044
rect 6276 23001 6285 23035
rect 6285 23001 6319 23035
rect 6319 23001 6328 23035
rect 6276 22992 6328 23001
rect 6736 22992 6788 23044
rect 9036 23060 9088 23112
rect 7656 22992 7708 23044
rect 8392 23035 8444 23044
rect 8392 23001 8401 23035
rect 8401 23001 8435 23035
rect 8435 23001 8444 23035
rect 8392 22992 8444 23001
rect 10416 23103 10468 23112
rect 10416 23069 10425 23103
rect 10425 23069 10459 23103
rect 10459 23069 10468 23103
rect 10416 23060 10468 23069
rect 10508 23103 10560 23112
rect 10508 23069 10517 23103
rect 10517 23069 10551 23103
rect 10551 23069 10560 23103
rect 10508 23060 10560 23069
rect 10600 23103 10652 23112
rect 10600 23069 10609 23103
rect 10609 23069 10643 23103
rect 10643 23069 10652 23103
rect 10600 23060 10652 23069
rect 10876 23103 10928 23112
rect 10876 23069 10885 23103
rect 10885 23069 10919 23103
rect 10919 23069 10928 23103
rect 12164 23171 12216 23180
rect 12164 23137 12173 23171
rect 12173 23137 12207 23171
rect 12207 23137 12216 23171
rect 12164 23128 12216 23137
rect 12900 23128 12952 23180
rect 14188 23171 14240 23180
rect 14188 23137 14197 23171
rect 14197 23137 14231 23171
rect 14231 23137 14240 23171
rect 14188 23128 14240 23137
rect 14556 23128 14608 23180
rect 22284 23128 22336 23180
rect 10876 23060 10928 23069
rect 15016 23060 15068 23112
rect 15752 23060 15804 23112
rect 17040 23103 17092 23112
rect 17040 23069 17049 23103
rect 17049 23069 17083 23103
rect 17083 23069 17092 23103
rect 17040 23060 17092 23069
rect 19432 23103 19484 23112
rect 19432 23069 19441 23103
rect 19441 23069 19475 23103
rect 19475 23069 19484 23103
rect 19432 23060 19484 23069
rect 21180 23060 21232 23112
rect 21916 23103 21968 23112
rect 21916 23069 21925 23103
rect 21925 23069 21959 23103
rect 21959 23069 21968 23103
rect 21916 23060 21968 23069
rect 23296 23264 23348 23316
rect 24032 23264 24084 23316
rect 25780 23264 25832 23316
rect 22928 23128 22980 23180
rect 23112 23103 23164 23112
rect 23112 23069 23121 23103
rect 23121 23069 23155 23103
rect 23155 23069 23164 23103
rect 23112 23060 23164 23069
rect 24492 23128 24544 23180
rect 24768 23171 24820 23180
rect 24768 23137 24777 23171
rect 24777 23137 24811 23171
rect 24811 23137 24820 23171
rect 24768 23128 24820 23137
rect 25596 23196 25648 23248
rect 26976 23307 27028 23316
rect 26976 23273 26985 23307
rect 26985 23273 27019 23307
rect 27019 23273 27028 23307
rect 26976 23264 27028 23273
rect 26240 23128 26292 23180
rect 26608 23128 26660 23180
rect 22008 23035 22060 23044
rect 22008 23001 22017 23035
rect 22017 23001 22051 23035
rect 22051 23001 22060 23035
rect 22008 22992 22060 23001
rect 22652 22992 22704 23044
rect 6368 22924 6420 22976
rect 8116 22924 8168 22976
rect 8852 22924 8904 22976
rect 9588 22924 9640 22976
rect 11060 22967 11112 22976
rect 11060 22933 11069 22967
rect 11069 22933 11103 22967
rect 11103 22933 11112 22967
rect 11060 22924 11112 22933
rect 12624 22967 12676 22976
rect 12624 22933 12633 22967
rect 12633 22933 12667 22967
rect 12667 22933 12676 22967
rect 12624 22924 12676 22933
rect 12716 22924 12768 22976
rect 14648 22967 14700 22976
rect 14648 22933 14657 22967
rect 14657 22933 14691 22967
rect 14691 22933 14700 22967
rect 14648 22924 14700 22933
rect 18420 22924 18472 22976
rect 18880 22924 18932 22976
rect 19340 22924 19392 22976
rect 22100 22924 22152 22976
rect 23020 22967 23072 22976
rect 23020 22933 23029 22967
rect 23029 22933 23063 22967
rect 23063 22933 23072 22967
rect 23020 22924 23072 22933
rect 24216 23060 24268 23112
rect 25412 23103 25464 23112
rect 25412 23069 25421 23103
rect 25421 23069 25455 23103
rect 25455 23069 25464 23103
rect 25412 23060 25464 23069
rect 26056 23060 26108 23112
rect 26608 23035 26660 23044
rect 26608 23001 26617 23035
rect 26617 23001 26651 23035
rect 26651 23001 26660 23035
rect 26608 22992 26660 23001
rect 27160 22992 27212 23044
rect 27436 23060 27488 23112
rect 24860 22924 24912 22976
rect 25412 22967 25464 22976
rect 25412 22933 25421 22967
rect 25421 22933 25455 22967
rect 25455 22933 25464 22967
rect 25412 22924 25464 22933
rect 26148 22924 26200 22976
rect 27344 22967 27396 22976
rect 27344 22933 27353 22967
rect 27353 22933 27387 22967
rect 27387 22933 27396 22967
rect 27344 22924 27396 22933
rect 27528 22924 27580 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 2872 22720 2924 22772
rect 3792 22695 3844 22704
rect 3792 22661 3801 22695
rect 3801 22661 3835 22695
rect 3835 22661 3844 22695
rect 3792 22652 3844 22661
rect 4068 22763 4120 22772
rect 4068 22729 4077 22763
rect 4077 22729 4111 22763
rect 4111 22729 4120 22763
rect 4068 22720 4120 22729
rect 4252 22652 4304 22704
rect 8392 22720 8444 22772
rect 9588 22720 9640 22772
rect 10600 22720 10652 22772
rect 18420 22720 18472 22772
rect 18880 22763 18932 22772
rect 18880 22729 18889 22763
rect 18889 22729 18923 22763
rect 18923 22729 18932 22763
rect 18880 22720 18932 22729
rect 22284 22720 22336 22772
rect 23020 22720 23072 22772
rect 25136 22720 25188 22772
rect 8116 22695 8168 22704
rect 8116 22661 8125 22695
rect 8125 22661 8159 22695
rect 8159 22661 8168 22695
rect 8116 22652 8168 22661
rect 8852 22695 8904 22704
rect 8852 22661 8861 22695
rect 8861 22661 8895 22695
rect 8895 22661 8904 22695
rect 8852 22652 8904 22661
rect 2320 22584 2372 22636
rect 3148 22584 3200 22636
rect 6736 22627 6788 22636
rect 6736 22593 6745 22627
rect 6745 22593 6779 22627
rect 6779 22593 6788 22627
rect 6736 22584 6788 22593
rect 6920 22627 6972 22636
rect 6920 22593 6929 22627
rect 6929 22593 6963 22627
rect 6963 22593 6972 22627
rect 6920 22584 6972 22593
rect 7472 22627 7524 22636
rect 7472 22593 7481 22627
rect 7481 22593 7515 22627
rect 7515 22593 7524 22627
rect 7472 22584 7524 22593
rect 7656 22627 7708 22636
rect 7656 22593 7665 22627
rect 7665 22593 7699 22627
rect 7699 22593 7708 22627
rect 7656 22584 7708 22593
rect 7840 22627 7892 22636
rect 7840 22593 7849 22627
rect 7849 22593 7883 22627
rect 7883 22593 7892 22627
rect 7840 22584 7892 22593
rect 9036 22627 9088 22636
rect 2136 22516 2188 22568
rect 2964 22516 3016 22568
rect 3608 22559 3660 22568
rect 3608 22525 3617 22559
rect 3617 22525 3651 22559
rect 3651 22525 3660 22559
rect 3608 22516 3660 22525
rect 4804 22448 4856 22500
rect 9036 22593 9045 22627
rect 9045 22593 9079 22627
rect 9079 22593 9088 22627
rect 9036 22584 9088 22593
rect 9312 22584 9364 22636
rect 11060 22652 11112 22704
rect 10232 22584 10284 22636
rect 12624 22627 12676 22636
rect 12624 22593 12633 22627
rect 12633 22593 12667 22627
rect 12667 22593 12676 22627
rect 12624 22584 12676 22593
rect 13176 22584 13228 22636
rect 18696 22652 18748 22704
rect 22008 22652 22060 22704
rect 22376 22695 22428 22704
rect 22376 22661 22385 22695
rect 22385 22661 22419 22695
rect 22419 22661 22428 22695
rect 22376 22652 22428 22661
rect 25596 22720 25648 22772
rect 26148 22720 26200 22772
rect 27160 22720 27212 22772
rect 3884 22380 3936 22432
rect 16856 22516 16908 22568
rect 18880 22584 18932 22636
rect 18972 22584 19024 22636
rect 19524 22584 19576 22636
rect 20720 22584 20772 22636
rect 25688 22695 25740 22704
rect 25688 22661 25697 22695
rect 25697 22661 25731 22695
rect 25731 22661 25740 22695
rect 25688 22652 25740 22661
rect 26056 22652 26108 22704
rect 25964 22584 26016 22636
rect 27068 22584 27120 22636
rect 21180 22516 21232 22568
rect 23112 22516 23164 22568
rect 25596 22516 25648 22568
rect 26148 22516 26200 22568
rect 27528 22720 27580 22772
rect 27344 22584 27396 22636
rect 18880 22448 18932 22500
rect 19432 22448 19484 22500
rect 24676 22448 24728 22500
rect 14188 22380 14240 22432
rect 18236 22423 18288 22432
rect 18236 22389 18245 22423
rect 18245 22389 18279 22423
rect 18279 22389 18288 22423
rect 18236 22380 18288 22389
rect 18420 22380 18472 22432
rect 18604 22380 18656 22432
rect 19340 22423 19392 22432
rect 19340 22389 19349 22423
rect 19349 22389 19383 22423
rect 19383 22389 19392 22423
rect 19340 22380 19392 22389
rect 24952 22491 25004 22500
rect 24952 22457 24961 22491
rect 24961 22457 24995 22491
rect 24995 22457 25004 22491
rect 24952 22448 25004 22457
rect 25228 22448 25280 22500
rect 25688 22448 25740 22500
rect 27712 22491 27764 22500
rect 27712 22457 27721 22491
rect 27721 22457 27755 22491
rect 27755 22457 27764 22491
rect 27712 22448 27764 22457
rect 25780 22380 25832 22432
rect 26056 22380 26108 22432
rect 27528 22380 27580 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 12624 22219 12676 22228
rect 12624 22185 12633 22219
rect 12633 22185 12667 22219
rect 12667 22185 12676 22219
rect 12624 22176 12676 22185
rect 14280 22176 14332 22228
rect 17224 22176 17276 22228
rect 21180 22219 21232 22228
rect 21180 22185 21189 22219
rect 21189 22185 21223 22219
rect 21223 22185 21232 22219
rect 21180 22176 21232 22185
rect 24216 22176 24268 22228
rect 2320 22040 2372 22092
rect 4068 22108 4120 22160
rect 1400 22015 1452 22024
rect 1400 21981 1409 22015
rect 1409 21981 1443 22015
rect 1443 21981 1452 22015
rect 1400 21972 1452 21981
rect 2688 22015 2740 22024
rect 2688 21981 2697 22015
rect 2697 21981 2731 22015
rect 2731 21981 2740 22015
rect 2688 21972 2740 21981
rect 2872 22015 2924 22024
rect 2872 21981 2881 22015
rect 2881 21981 2915 22015
rect 2915 21981 2924 22015
rect 2872 21972 2924 21981
rect 2136 21904 2188 21956
rect 4068 21972 4120 22024
rect 4804 22015 4856 22024
rect 4804 21981 4813 22015
rect 4813 21981 4847 22015
rect 4847 21981 4856 22015
rect 4804 21972 4856 21981
rect 5264 22015 5316 22024
rect 5264 21981 5273 22015
rect 5273 21981 5307 22015
rect 5307 21981 5316 22015
rect 5264 21972 5316 21981
rect 9312 21972 9364 22024
rect 9588 22015 9640 22024
rect 9588 21981 9597 22015
rect 9597 21981 9631 22015
rect 9631 21981 9640 22015
rect 9588 21972 9640 21981
rect 10232 21972 10284 22024
rect 11888 22015 11940 22024
rect 3056 21836 3108 21888
rect 3884 21836 3936 21888
rect 3976 21879 4028 21888
rect 3976 21845 3985 21879
rect 3985 21845 4019 21879
rect 4019 21845 4028 21879
rect 3976 21836 4028 21845
rect 6092 21904 6144 21956
rect 11888 21981 11897 22015
rect 11897 21981 11931 22015
rect 11931 21981 11940 22015
rect 11888 21972 11940 21981
rect 12164 22015 12216 22024
rect 12164 21981 12173 22015
rect 12173 21981 12207 22015
rect 12207 21981 12216 22015
rect 12164 21972 12216 21981
rect 14372 22040 14424 22092
rect 14740 22040 14792 22092
rect 16212 22040 16264 22092
rect 12532 21972 12584 22024
rect 15016 21972 15068 22024
rect 15292 21972 15344 22024
rect 4620 21836 4672 21888
rect 11704 21879 11756 21888
rect 11704 21845 11713 21879
rect 11713 21845 11747 21879
rect 11747 21845 11756 21879
rect 11704 21836 11756 21845
rect 14280 21904 14332 21956
rect 12716 21836 12768 21888
rect 14096 21836 14148 21888
rect 14648 21947 14700 21956
rect 14648 21913 14673 21947
rect 14673 21913 14700 21947
rect 14648 21904 14700 21913
rect 14556 21836 14608 21888
rect 14832 21879 14884 21888
rect 14832 21845 14841 21879
rect 14841 21845 14875 21879
rect 14875 21845 14884 21879
rect 14832 21836 14884 21845
rect 17224 22040 17276 22092
rect 19064 22040 19116 22092
rect 20720 22083 20772 22092
rect 20720 22049 20729 22083
rect 20729 22049 20763 22083
rect 20763 22049 20772 22083
rect 20720 22040 20772 22049
rect 25228 22176 25280 22228
rect 25320 22176 25372 22228
rect 22192 21972 22244 22024
rect 16948 21879 17000 21888
rect 16948 21845 16957 21879
rect 16957 21845 16991 21879
rect 16991 21845 17000 21879
rect 16948 21836 17000 21845
rect 17316 21947 17368 21956
rect 17316 21913 17325 21947
rect 17325 21913 17359 21947
rect 17359 21913 17368 21947
rect 17316 21904 17368 21913
rect 21088 21904 21140 21956
rect 25412 22108 25464 22160
rect 24584 22015 24636 22024
rect 24584 21981 24593 22015
rect 24593 21981 24627 22015
rect 24627 21981 24636 22015
rect 24584 21972 24636 21981
rect 24676 22015 24728 22024
rect 24676 21981 24685 22015
rect 24685 21981 24719 22015
rect 24719 21981 24728 22015
rect 24676 21972 24728 21981
rect 24860 22015 24912 22024
rect 24860 21981 24869 22015
rect 24869 21981 24903 22015
rect 24903 21981 24912 22015
rect 25688 22040 25740 22092
rect 24860 21972 24912 21981
rect 25596 21972 25648 22024
rect 25872 21972 25924 22024
rect 26240 21972 26292 22024
rect 27528 22015 27580 22024
rect 27528 21981 27537 22015
rect 27537 21981 27571 22015
rect 27571 21981 27580 22015
rect 27528 21972 27580 21981
rect 19432 21836 19484 21888
rect 25964 21904 26016 21956
rect 24584 21836 24636 21888
rect 24768 21836 24820 21888
rect 25136 21836 25188 21888
rect 25688 21879 25740 21888
rect 25688 21845 25697 21879
rect 25697 21845 25731 21879
rect 25731 21845 25740 21879
rect 25688 21836 25740 21845
rect 25872 21836 25924 21888
rect 27712 21879 27764 21888
rect 27712 21845 27721 21879
rect 27721 21845 27755 21879
rect 27755 21845 27764 21879
rect 27712 21836 27764 21845
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 14280 21675 14332 21684
rect 14280 21641 14289 21675
rect 14289 21641 14323 21675
rect 14323 21641 14332 21675
rect 14280 21632 14332 21641
rect 1308 21564 1360 21616
rect 2964 21564 3016 21616
rect 7472 21564 7524 21616
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 2320 21496 2372 21548
rect 3608 21539 3660 21548
rect 3608 21505 3617 21539
rect 3617 21505 3651 21539
rect 3651 21505 3660 21539
rect 3608 21496 3660 21505
rect 3976 21539 4028 21548
rect 3976 21505 3985 21539
rect 3985 21505 4019 21539
rect 4019 21505 4028 21539
rect 3976 21496 4028 21505
rect 4804 21496 4856 21548
rect 5264 21496 5316 21548
rect 7656 21496 7708 21548
rect 14096 21564 14148 21616
rect 12072 21496 12124 21548
rect 15016 21632 15068 21684
rect 17224 21632 17276 21684
rect 25136 21632 25188 21684
rect 25228 21632 25280 21684
rect 4712 21428 4764 21480
rect 5724 21471 5776 21480
rect 5724 21437 5733 21471
rect 5733 21437 5767 21471
rect 5767 21437 5776 21471
rect 5724 21428 5776 21437
rect 6092 21428 6144 21480
rect 14004 21471 14056 21480
rect 14004 21437 14013 21471
rect 14013 21437 14047 21471
rect 14047 21437 14056 21471
rect 14004 21428 14056 21437
rect 8576 21403 8628 21412
rect 8576 21369 8585 21403
rect 8585 21369 8619 21403
rect 8619 21369 8628 21403
rect 8576 21360 8628 21369
rect 13820 21360 13872 21412
rect 15292 21539 15344 21548
rect 15292 21505 15301 21539
rect 15301 21505 15335 21539
rect 15335 21505 15344 21539
rect 15292 21496 15344 21505
rect 17040 21564 17092 21616
rect 17316 21564 17368 21616
rect 18880 21564 18932 21616
rect 16212 21539 16264 21548
rect 16212 21505 16221 21539
rect 16221 21505 16255 21539
rect 16255 21505 16264 21539
rect 16212 21496 16264 21505
rect 16396 21496 16448 21548
rect 14372 21428 14424 21480
rect 14648 21428 14700 21480
rect 14832 21428 14884 21480
rect 16764 21471 16816 21480
rect 16764 21437 16773 21471
rect 16773 21437 16807 21471
rect 16807 21437 16816 21471
rect 16764 21428 16816 21437
rect 17592 21496 17644 21548
rect 18144 21496 18196 21548
rect 18328 21496 18380 21548
rect 18420 21496 18472 21548
rect 18604 21539 18656 21548
rect 18604 21505 18613 21539
rect 18613 21505 18647 21539
rect 18647 21505 18656 21539
rect 18604 21496 18656 21505
rect 19616 21564 19668 21616
rect 6920 21292 6972 21344
rect 13912 21335 13964 21344
rect 13912 21301 13921 21335
rect 13921 21301 13955 21335
rect 13955 21301 13964 21335
rect 13912 21292 13964 21301
rect 14464 21292 14516 21344
rect 14740 21292 14792 21344
rect 14832 21292 14884 21344
rect 15384 21360 15436 21412
rect 16580 21360 16632 21412
rect 18052 21428 18104 21480
rect 19064 21496 19116 21548
rect 24676 21564 24728 21616
rect 25320 21607 25372 21616
rect 25320 21573 25329 21607
rect 25329 21573 25363 21607
rect 25363 21573 25372 21607
rect 25320 21564 25372 21573
rect 25412 21564 25464 21616
rect 27436 21632 27488 21684
rect 19432 21471 19484 21480
rect 19432 21437 19441 21471
rect 19441 21437 19475 21471
rect 19475 21437 19484 21471
rect 19432 21428 19484 21437
rect 17224 21360 17276 21412
rect 19984 21360 20036 21412
rect 24584 21496 24636 21548
rect 24768 21539 24820 21548
rect 24768 21505 24777 21539
rect 24777 21505 24811 21539
rect 24811 21505 24820 21539
rect 24768 21496 24820 21505
rect 27804 21539 27856 21548
rect 27804 21505 27813 21539
rect 27813 21505 27847 21539
rect 27847 21505 27856 21539
rect 27804 21496 27856 21505
rect 24676 21428 24728 21480
rect 26056 21428 26108 21480
rect 24952 21360 25004 21412
rect 15016 21292 15068 21344
rect 17040 21292 17092 21344
rect 24216 21292 24268 21344
rect 25872 21292 25924 21344
rect 27620 21335 27672 21344
rect 27620 21301 27629 21335
rect 27629 21301 27663 21335
rect 27663 21301 27672 21335
rect 27620 21292 27672 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 12164 21088 12216 21140
rect 15108 21088 15160 21140
rect 15200 21088 15252 21140
rect 2320 20952 2372 21004
rect 2596 20884 2648 20936
rect 4620 20884 4672 20936
rect 5264 20927 5316 20936
rect 5264 20893 5273 20927
rect 5273 20893 5307 20927
rect 5307 20893 5316 20927
rect 5264 20884 5316 20893
rect 5724 20884 5776 20936
rect 6092 20927 6144 20936
rect 6092 20893 6101 20927
rect 6101 20893 6135 20927
rect 6135 20893 6144 20927
rect 6092 20884 6144 20893
rect 7104 20884 7156 20936
rect 6552 20816 6604 20868
rect 11152 20927 11204 20936
rect 11152 20893 11161 20927
rect 11161 20893 11195 20927
rect 11195 20893 11204 20927
rect 11152 20884 11204 20893
rect 11520 20995 11572 21004
rect 11520 20961 11529 20995
rect 11529 20961 11563 20995
rect 11563 20961 11572 20995
rect 11520 20952 11572 20961
rect 12072 20995 12124 21004
rect 12072 20961 12081 20995
rect 12081 20961 12115 20995
rect 12115 20961 12124 20995
rect 12072 20952 12124 20961
rect 12808 20952 12860 21004
rect 14740 20952 14792 21004
rect 15844 21020 15896 21072
rect 11336 20884 11388 20936
rect 11612 20927 11664 20936
rect 11612 20893 11621 20927
rect 11621 20893 11655 20927
rect 11655 20893 11664 20927
rect 11612 20884 11664 20893
rect 12532 20884 12584 20936
rect 13176 20884 13228 20936
rect 13544 20884 13596 20936
rect 14096 20884 14148 20936
rect 14372 20884 14424 20936
rect 14556 20927 14608 20936
rect 14556 20893 14565 20927
rect 14565 20893 14599 20927
rect 14599 20893 14608 20927
rect 14556 20884 14608 20893
rect 14924 20927 14976 20936
rect 14924 20893 14933 20927
rect 14933 20893 14967 20927
rect 14967 20893 14976 20927
rect 14924 20884 14976 20893
rect 17224 21131 17276 21140
rect 17224 21097 17233 21131
rect 17233 21097 17267 21131
rect 17267 21097 17276 21131
rect 17224 21088 17276 21097
rect 18328 21088 18380 21140
rect 18788 21088 18840 21140
rect 19064 21088 19116 21140
rect 21456 21088 21508 21140
rect 16580 21020 16632 21072
rect 16764 20952 16816 21004
rect 17132 20952 17184 21004
rect 17592 20995 17644 21004
rect 17592 20961 17601 20995
rect 17601 20961 17635 20995
rect 17635 20961 17644 20995
rect 17592 20952 17644 20961
rect 18420 20952 18472 21004
rect 2044 20748 2096 20800
rect 6276 20748 6328 20800
rect 8300 20859 8352 20868
rect 8300 20825 8309 20859
rect 8309 20825 8343 20859
rect 8343 20825 8352 20859
rect 8300 20816 8352 20825
rect 11888 20859 11940 20868
rect 11888 20825 11897 20859
rect 11897 20825 11931 20859
rect 11931 20825 11940 20859
rect 11888 20816 11940 20825
rect 14740 20816 14792 20868
rect 16212 20884 16264 20936
rect 17776 20884 17828 20936
rect 18052 20884 18104 20936
rect 19892 21063 19944 21072
rect 19892 21029 19901 21063
rect 19901 21029 19935 21063
rect 19935 21029 19944 21063
rect 19892 21020 19944 21029
rect 20444 21063 20496 21072
rect 20444 21029 20453 21063
rect 20453 21029 20487 21063
rect 20487 21029 20496 21063
rect 22652 21088 22704 21140
rect 20444 21020 20496 21029
rect 22192 21020 22244 21072
rect 16488 20859 16540 20868
rect 16488 20825 16497 20859
rect 16497 20825 16531 20859
rect 16531 20825 16540 20859
rect 16488 20816 16540 20825
rect 13544 20791 13596 20800
rect 13544 20757 13553 20791
rect 13553 20757 13587 20791
rect 13587 20757 13596 20791
rect 13544 20748 13596 20757
rect 14280 20748 14332 20800
rect 14464 20748 14516 20800
rect 15200 20748 15252 20800
rect 15476 20748 15528 20800
rect 18144 20816 18196 20868
rect 18788 20927 18840 20936
rect 18788 20893 18797 20927
rect 18797 20893 18831 20927
rect 18831 20893 18840 20927
rect 18788 20884 18840 20893
rect 19064 20927 19116 20936
rect 18696 20816 18748 20868
rect 19064 20893 19073 20927
rect 19073 20893 19107 20927
rect 19107 20893 19116 20927
rect 19064 20884 19116 20893
rect 19156 20884 19208 20936
rect 19708 20884 19760 20936
rect 19892 20884 19944 20936
rect 19984 20927 20036 20936
rect 19984 20893 19993 20927
rect 19993 20893 20027 20927
rect 20027 20893 20036 20927
rect 19984 20884 20036 20893
rect 20076 20927 20128 20936
rect 20076 20893 20085 20927
rect 20085 20893 20119 20927
rect 20119 20893 20128 20927
rect 20076 20884 20128 20893
rect 18328 20748 18380 20800
rect 18420 20791 18472 20800
rect 18420 20757 18429 20791
rect 18429 20757 18463 20791
rect 18463 20757 18472 20791
rect 18420 20748 18472 20757
rect 18788 20748 18840 20800
rect 19800 20748 19852 20800
rect 21548 20952 21600 21004
rect 21456 20884 21508 20936
rect 25044 20952 25096 21004
rect 21824 20884 21876 20936
rect 21548 20816 21600 20868
rect 22376 20927 22428 20936
rect 22376 20893 22385 20927
rect 22385 20893 22419 20927
rect 22419 20893 22428 20927
rect 22376 20884 22428 20893
rect 22468 20884 22520 20936
rect 23572 20884 23624 20936
rect 24676 20927 24728 20936
rect 24676 20893 24685 20927
rect 24685 20893 24719 20927
rect 24719 20893 24728 20927
rect 24676 20884 24728 20893
rect 24032 20816 24084 20868
rect 25412 20816 25464 20868
rect 21916 20748 21968 20800
rect 22100 20748 22152 20800
rect 26424 20791 26476 20800
rect 26424 20757 26433 20791
rect 26433 20757 26467 20791
rect 26467 20757 26476 20791
rect 26424 20748 26476 20757
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 11612 20544 11664 20596
rect 13820 20544 13872 20596
rect 2044 20451 2096 20460
rect 2044 20417 2053 20451
rect 2053 20417 2087 20451
rect 2087 20417 2096 20451
rect 2044 20408 2096 20417
rect 2228 20451 2280 20460
rect 2228 20417 2237 20451
rect 2237 20417 2271 20451
rect 2271 20417 2280 20451
rect 2228 20408 2280 20417
rect 2780 20408 2832 20460
rect 11152 20476 11204 20528
rect 3424 20383 3476 20392
rect 3424 20349 3433 20383
rect 3433 20349 3467 20383
rect 3467 20349 3476 20383
rect 3424 20340 3476 20349
rect 6276 20408 6328 20460
rect 6920 20451 6972 20460
rect 6920 20417 6929 20451
rect 6929 20417 6963 20451
rect 6963 20417 6972 20451
rect 6920 20408 6972 20417
rect 7932 20451 7984 20460
rect 7932 20417 7941 20451
rect 7941 20417 7975 20451
rect 7975 20417 7984 20451
rect 7932 20408 7984 20417
rect 8300 20408 8352 20460
rect 11060 20451 11112 20460
rect 11060 20417 11069 20451
rect 11069 20417 11103 20451
rect 11103 20417 11112 20451
rect 11060 20408 11112 20417
rect 11244 20451 11296 20460
rect 11244 20417 11253 20451
rect 11253 20417 11287 20451
rect 11287 20417 11296 20451
rect 11244 20408 11296 20417
rect 11336 20451 11388 20460
rect 11336 20417 11345 20451
rect 11345 20417 11379 20451
rect 11379 20417 11388 20451
rect 11336 20408 11388 20417
rect 11520 20519 11572 20528
rect 11520 20485 11529 20519
rect 11529 20485 11563 20519
rect 11563 20485 11572 20519
rect 11520 20476 11572 20485
rect 11796 20408 11848 20460
rect 12256 20476 12308 20528
rect 13544 20476 13596 20528
rect 14924 20544 14976 20596
rect 15108 20544 15160 20596
rect 16948 20544 17000 20596
rect 12348 20451 12400 20460
rect 12348 20417 12357 20451
rect 12357 20417 12391 20451
rect 12391 20417 12400 20451
rect 12348 20408 12400 20417
rect 12440 20451 12492 20460
rect 12440 20417 12449 20451
rect 12449 20417 12483 20451
rect 12483 20417 12492 20451
rect 12440 20408 12492 20417
rect 13268 20451 13320 20460
rect 13268 20417 13277 20451
rect 13277 20417 13311 20451
rect 13311 20417 13320 20451
rect 13268 20408 13320 20417
rect 12624 20340 12676 20392
rect 13820 20408 13872 20460
rect 16580 20476 16632 20528
rect 15016 20451 15068 20460
rect 15016 20417 15025 20451
rect 15025 20417 15059 20451
rect 15059 20417 15068 20451
rect 15016 20408 15068 20417
rect 15200 20408 15252 20460
rect 15292 20451 15344 20460
rect 15292 20417 15301 20451
rect 15301 20417 15335 20451
rect 15335 20417 15344 20451
rect 15292 20408 15344 20417
rect 15384 20451 15436 20460
rect 15384 20417 15393 20451
rect 15393 20417 15427 20451
rect 15427 20417 15436 20451
rect 15384 20408 15436 20417
rect 15476 20451 15528 20460
rect 15476 20417 15485 20451
rect 15485 20417 15519 20451
rect 15519 20417 15528 20451
rect 15476 20408 15528 20417
rect 16764 20408 16816 20460
rect 17040 20476 17092 20528
rect 18420 20544 18472 20596
rect 18880 20544 18932 20596
rect 8392 20272 8444 20324
rect 11244 20272 11296 20324
rect 12164 20272 12216 20324
rect 13728 20272 13780 20324
rect 3148 20204 3200 20256
rect 11060 20204 11112 20256
rect 12256 20204 12308 20256
rect 13544 20247 13596 20256
rect 13544 20213 13553 20247
rect 13553 20213 13587 20247
rect 13587 20213 13596 20247
rect 13544 20204 13596 20213
rect 14556 20340 14608 20392
rect 14740 20340 14792 20392
rect 16488 20340 16540 20392
rect 17960 20451 18012 20460
rect 17960 20417 17969 20451
rect 17969 20417 18003 20451
rect 18003 20417 18012 20451
rect 17960 20408 18012 20417
rect 18604 20408 18656 20460
rect 18972 20451 19024 20460
rect 18972 20417 18981 20451
rect 18981 20417 19015 20451
rect 19015 20417 19024 20451
rect 18972 20408 19024 20417
rect 19800 20476 19852 20528
rect 19248 20451 19300 20460
rect 19248 20417 19257 20451
rect 19257 20417 19291 20451
rect 19291 20417 19300 20451
rect 19248 20408 19300 20417
rect 19340 20451 19392 20460
rect 19340 20417 19349 20451
rect 19349 20417 19383 20451
rect 19383 20417 19392 20451
rect 19340 20408 19392 20417
rect 22376 20544 22428 20596
rect 23572 20587 23624 20596
rect 23572 20553 23581 20587
rect 23581 20553 23615 20587
rect 23615 20553 23624 20587
rect 23572 20544 23624 20553
rect 20076 20476 20128 20528
rect 20536 20519 20588 20528
rect 20536 20485 20545 20519
rect 20545 20485 20579 20519
rect 20579 20485 20588 20519
rect 20536 20476 20588 20485
rect 22100 20519 22152 20528
rect 22100 20485 22109 20519
rect 22109 20485 22143 20519
rect 22143 20485 22152 20519
rect 22100 20476 22152 20485
rect 22560 20476 22612 20528
rect 25228 20476 25280 20528
rect 26424 20476 26476 20528
rect 21180 20451 21232 20460
rect 21180 20417 21189 20451
rect 21189 20417 21223 20451
rect 21223 20417 21232 20451
rect 21180 20408 21232 20417
rect 20996 20340 21048 20392
rect 21364 20451 21416 20460
rect 21364 20417 21373 20451
rect 21373 20417 21407 20451
rect 21407 20417 21416 20451
rect 21364 20408 21416 20417
rect 21548 20451 21600 20460
rect 21548 20417 21557 20451
rect 21557 20417 21591 20451
rect 21591 20417 21600 20451
rect 21548 20408 21600 20417
rect 19708 20272 19760 20324
rect 21456 20340 21508 20392
rect 16396 20204 16448 20256
rect 17500 20204 17552 20256
rect 18972 20204 19024 20256
rect 20628 20204 20680 20256
rect 20904 20204 20956 20256
rect 21088 20204 21140 20256
rect 21824 20383 21876 20392
rect 21824 20349 21833 20383
rect 21833 20349 21867 20383
rect 21867 20349 21876 20383
rect 21824 20340 21876 20349
rect 22560 20340 22612 20392
rect 24032 20340 24084 20392
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 12440 20000 12492 20052
rect 13268 20000 13320 20052
rect 13728 20000 13780 20052
rect 15292 20000 15344 20052
rect 19340 20000 19392 20052
rect 19432 20000 19484 20052
rect 19708 20000 19760 20052
rect 20628 20000 20680 20052
rect 21180 20000 21232 20052
rect 22652 20043 22704 20052
rect 22652 20009 22661 20043
rect 22661 20009 22695 20043
rect 22695 20009 22704 20043
rect 22652 20000 22704 20009
rect 23296 20000 23348 20052
rect 27804 20043 27856 20052
rect 27804 20009 27813 20043
rect 27813 20009 27847 20043
rect 27847 20009 27856 20043
rect 27804 20000 27856 20009
rect 2596 19932 2648 19984
rect 2044 19907 2096 19916
rect 2044 19873 2053 19907
rect 2053 19873 2087 19907
rect 2087 19873 2096 19907
rect 2044 19864 2096 19873
rect 2688 19907 2740 19916
rect 2688 19873 2697 19907
rect 2697 19873 2731 19907
rect 2731 19873 2740 19907
rect 2688 19864 2740 19873
rect 3148 19907 3200 19916
rect 3148 19873 3157 19907
rect 3157 19873 3191 19907
rect 3191 19873 3200 19907
rect 3148 19864 3200 19873
rect 3424 19907 3476 19916
rect 3424 19873 3433 19907
rect 3433 19873 3467 19907
rect 3467 19873 3476 19907
rect 3424 19864 3476 19873
rect 848 19796 900 19848
rect 2228 19796 2280 19848
rect 2964 19728 3016 19780
rect 4712 19839 4764 19848
rect 4712 19805 4721 19839
rect 4721 19805 4755 19839
rect 4755 19805 4764 19839
rect 4712 19796 4764 19805
rect 12348 19932 12400 19984
rect 14004 19932 14056 19984
rect 15016 19932 15068 19984
rect 18972 19932 19024 19984
rect 8300 19864 8352 19916
rect 11612 19864 11664 19916
rect 6368 19796 6420 19848
rect 7932 19796 7984 19848
rect 12532 19864 12584 19916
rect 14188 19864 14240 19916
rect 14740 19864 14792 19916
rect 17960 19864 18012 19916
rect 12808 19839 12860 19848
rect 12808 19805 12817 19839
rect 12817 19805 12851 19839
rect 12851 19805 12860 19839
rect 12808 19796 12860 19805
rect 13636 19839 13688 19848
rect 13636 19805 13645 19839
rect 13645 19805 13679 19839
rect 13679 19805 13688 19839
rect 13636 19796 13688 19805
rect 4528 19728 4580 19780
rect 2320 19660 2372 19712
rect 9496 19728 9548 19780
rect 5356 19660 5408 19712
rect 6000 19660 6052 19712
rect 8760 19660 8812 19712
rect 12440 19728 12492 19780
rect 13912 19796 13964 19848
rect 14004 19728 14056 19780
rect 15108 19728 15160 19780
rect 20720 19796 20772 19848
rect 21088 19864 21140 19916
rect 22284 19932 22336 19984
rect 21456 19864 21508 19916
rect 11888 19660 11940 19712
rect 12256 19660 12308 19712
rect 15200 19660 15252 19712
rect 16488 19660 16540 19712
rect 20812 19728 20864 19780
rect 19800 19660 19852 19712
rect 19892 19660 19944 19712
rect 21364 19796 21416 19848
rect 21548 19728 21600 19780
rect 21640 19728 21692 19780
rect 22192 19864 22244 19916
rect 22560 19907 22612 19916
rect 22560 19873 22569 19907
rect 22569 19873 22603 19907
rect 22603 19873 22612 19907
rect 22560 19864 22612 19873
rect 23480 19864 23532 19916
rect 24676 19864 24728 19916
rect 22008 19839 22060 19848
rect 22008 19805 22017 19839
rect 22017 19805 22051 19839
rect 22051 19805 22060 19839
rect 22008 19796 22060 19805
rect 22100 19839 22152 19848
rect 22100 19805 22109 19839
rect 22109 19805 22143 19839
rect 22143 19805 22152 19839
rect 22100 19796 22152 19805
rect 22376 19839 22428 19848
rect 22376 19805 22385 19839
rect 22385 19805 22419 19839
rect 22419 19805 22428 19839
rect 22376 19796 22428 19805
rect 22284 19728 22336 19780
rect 25688 19728 25740 19780
rect 22008 19660 22060 19712
rect 22100 19660 22152 19712
rect 22928 19660 22980 19712
rect 24860 19660 24912 19712
rect 25504 19660 25556 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 1584 19320 1636 19372
rect 2596 19320 2648 19372
rect 2964 19363 3016 19372
rect 2964 19329 2973 19363
rect 2973 19329 3007 19363
rect 3007 19329 3016 19363
rect 2964 19320 3016 19329
rect 4068 19388 4120 19440
rect 5448 19456 5500 19508
rect 8392 19456 8444 19508
rect 12624 19456 12676 19508
rect 15016 19456 15068 19508
rect 4528 19431 4580 19440
rect 4528 19397 4537 19431
rect 4537 19397 4571 19431
rect 4571 19397 4580 19431
rect 4528 19388 4580 19397
rect 5264 19388 5316 19440
rect 3424 19295 3476 19304
rect 3424 19261 3433 19295
rect 3433 19261 3467 19295
rect 3467 19261 3476 19295
rect 3424 19252 3476 19261
rect 4068 19295 4120 19304
rect 4068 19261 4077 19295
rect 4077 19261 4111 19295
rect 4111 19261 4120 19295
rect 4068 19252 4120 19261
rect 4712 19252 4764 19304
rect 5356 19320 5408 19372
rect 6000 19363 6052 19372
rect 6000 19329 6009 19363
rect 6009 19329 6043 19363
rect 6043 19329 6052 19363
rect 6000 19320 6052 19329
rect 6092 19116 6144 19168
rect 6552 19363 6604 19372
rect 6552 19329 6561 19363
rect 6561 19329 6595 19363
rect 6595 19329 6604 19363
rect 6552 19320 6604 19329
rect 8208 19363 8260 19372
rect 8208 19329 8217 19363
rect 8217 19329 8251 19363
rect 8251 19329 8260 19363
rect 8208 19320 8260 19329
rect 8576 19363 8628 19372
rect 8576 19329 8585 19363
rect 8585 19329 8619 19363
rect 8619 19329 8628 19363
rect 8576 19320 8628 19329
rect 12440 19388 12492 19440
rect 13268 19388 13320 19440
rect 14096 19388 14148 19440
rect 14372 19388 14424 19440
rect 15108 19388 15160 19440
rect 16304 19388 16356 19440
rect 18788 19456 18840 19508
rect 20812 19456 20864 19508
rect 21640 19456 21692 19508
rect 12532 19320 12584 19372
rect 18052 19320 18104 19372
rect 18696 19363 18748 19372
rect 18696 19329 18705 19363
rect 18705 19329 18739 19363
rect 18739 19329 18748 19363
rect 18696 19320 18748 19329
rect 18972 19363 19024 19372
rect 18972 19329 18981 19363
rect 18981 19329 19015 19363
rect 19015 19329 19024 19363
rect 18972 19320 19024 19329
rect 19524 19388 19576 19440
rect 12716 19295 12768 19304
rect 12716 19261 12725 19295
rect 12725 19261 12759 19295
rect 12759 19261 12768 19295
rect 12716 19252 12768 19261
rect 9772 19227 9824 19236
rect 9772 19193 9781 19227
rect 9781 19193 9815 19227
rect 9815 19193 9824 19227
rect 9772 19184 9824 19193
rect 12992 19295 13044 19304
rect 12992 19261 13001 19295
rect 13001 19261 13035 19295
rect 13035 19261 13044 19295
rect 12992 19252 13044 19261
rect 14004 19252 14056 19304
rect 14372 19252 14424 19304
rect 19432 19363 19484 19372
rect 19432 19329 19441 19363
rect 19441 19329 19475 19363
rect 19475 19329 19484 19363
rect 19432 19320 19484 19329
rect 19800 19363 19852 19372
rect 19800 19329 19809 19363
rect 19809 19329 19843 19363
rect 19843 19329 19852 19363
rect 19800 19320 19852 19329
rect 19524 19295 19576 19304
rect 19524 19261 19533 19295
rect 19533 19261 19567 19295
rect 19567 19261 19576 19295
rect 19524 19252 19576 19261
rect 13728 19184 13780 19236
rect 21732 19388 21784 19440
rect 22376 19388 22428 19440
rect 20444 19320 20496 19372
rect 20720 19320 20772 19372
rect 20812 19363 20864 19372
rect 20812 19329 20821 19363
rect 20821 19329 20855 19363
rect 20855 19329 20864 19363
rect 20812 19320 20864 19329
rect 6460 19159 6512 19168
rect 6460 19125 6469 19159
rect 6469 19125 6503 19159
rect 6503 19125 6512 19159
rect 6460 19116 6512 19125
rect 8392 19116 8444 19168
rect 12532 19159 12584 19168
rect 12532 19125 12541 19159
rect 12541 19125 12575 19159
rect 12575 19125 12584 19159
rect 12532 19116 12584 19125
rect 13636 19116 13688 19168
rect 14464 19116 14516 19168
rect 18696 19116 18748 19168
rect 18972 19116 19024 19168
rect 22284 19227 22336 19236
rect 22284 19193 22293 19227
rect 22293 19193 22327 19227
rect 22327 19193 22336 19227
rect 22284 19184 22336 19193
rect 21640 19116 21692 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 8208 18955 8260 18964
rect 8208 18921 8217 18955
rect 8217 18921 8251 18955
rect 8251 18921 8260 18955
rect 8208 18912 8260 18921
rect 8668 18819 8720 18828
rect 8668 18785 8677 18819
rect 8677 18785 8711 18819
rect 8711 18785 8720 18819
rect 8668 18776 8720 18785
rect 4804 18708 4856 18760
rect 5356 18751 5408 18760
rect 5356 18717 5365 18751
rect 5365 18717 5399 18751
rect 5399 18717 5408 18751
rect 5356 18708 5408 18717
rect 6092 18751 6144 18760
rect 6092 18717 6101 18751
rect 6101 18717 6135 18751
rect 6135 18717 6144 18751
rect 6092 18708 6144 18717
rect 6552 18751 6604 18760
rect 6552 18717 6561 18751
rect 6561 18717 6595 18751
rect 6595 18717 6604 18751
rect 6552 18708 6604 18717
rect 8300 18708 8352 18760
rect 8576 18708 8628 18760
rect 8760 18751 8812 18760
rect 8760 18717 8769 18751
rect 8769 18717 8803 18751
rect 8803 18717 8812 18751
rect 8760 18708 8812 18717
rect 12348 18844 12400 18896
rect 13820 18912 13872 18964
rect 24216 18955 24268 18964
rect 24216 18921 24225 18955
rect 24225 18921 24259 18955
rect 24259 18921 24268 18955
rect 24216 18912 24268 18921
rect 13912 18776 13964 18828
rect 12900 18751 12952 18760
rect 12900 18717 12909 18751
rect 12909 18717 12943 18751
rect 12943 18717 12952 18751
rect 12900 18708 12952 18717
rect 13728 18751 13780 18760
rect 13728 18717 13737 18751
rect 13737 18717 13771 18751
rect 13771 18717 13780 18751
rect 13728 18708 13780 18717
rect 14372 18751 14424 18760
rect 14372 18717 14381 18751
rect 14381 18717 14415 18751
rect 14415 18717 14424 18751
rect 14372 18708 14424 18717
rect 14464 18751 14516 18760
rect 14464 18717 14473 18751
rect 14473 18717 14507 18751
rect 14507 18717 14516 18751
rect 14464 18708 14516 18717
rect 7656 18640 7708 18692
rect 14096 18640 14148 18692
rect 15384 18708 15436 18760
rect 21824 18819 21876 18828
rect 21824 18785 21833 18819
rect 21833 18785 21867 18819
rect 21867 18785 21876 18819
rect 21824 18776 21876 18785
rect 23388 18776 23440 18828
rect 18144 18751 18196 18760
rect 18144 18717 18153 18751
rect 18153 18717 18187 18751
rect 18187 18717 18196 18751
rect 18144 18708 18196 18717
rect 18420 18751 18472 18760
rect 18420 18717 18429 18751
rect 18429 18717 18463 18751
rect 18463 18717 18472 18751
rect 18420 18708 18472 18717
rect 5724 18615 5776 18624
rect 5724 18581 5733 18615
rect 5733 18581 5767 18615
rect 5767 18581 5776 18615
rect 5724 18572 5776 18581
rect 9220 18572 9272 18624
rect 9680 18615 9732 18624
rect 9680 18581 9689 18615
rect 9689 18581 9723 18615
rect 9723 18581 9732 18615
rect 9680 18572 9732 18581
rect 12716 18615 12768 18624
rect 12716 18581 12725 18615
rect 12725 18581 12759 18615
rect 12759 18581 12768 18615
rect 12716 18572 12768 18581
rect 13176 18615 13228 18624
rect 13176 18581 13185 18615
rect 13185 18581 13219 18615
rect 13219 18581 13228 18615
rect 13176 18572 13228 18581
rect 17316 18572 17368 18624
rect 18328 18640 18380 18692
rect 18512 18640 18564 18692
rect 18696 18751 18748 18760
rect 18696 18717 18705 18751
rect 18705 18717 18739 18751
rect 18739 18717 18748 18751
rect 18696 18708 18748 18717
rect 18972 18640 19024 18692
rect 19708 18640 19760 18692
rect 22744 18683 22796 18692
rect 22744 18649 22753 18683
rect 22753 18649 22787 18683
rect 22787 18649 22796 18683
rect 22744 18640 22796 18649
rect 24032 18640 24084 18692
rect 19248 18572 19300 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 4804 18368 4856 18420
rect 1952 18343 2004 18352
rect 1952 18309 1961 18343
rect 1961 18309 1995 18343
rect 1995 18309 2004 18343
rect 1952 18300 2004 18309
rect 2320 18343 2372 18352
rect 2320 18309 2329 18343
rect 2329 18309 2363 18343
rect 2363 18309 2372 18343
rect 2320 18300 2372 18309
rect 1492 18275 1544 18284
rect 1492 18241 1501 18275
rect 1501 18241 1535 18275
rect 1535 18241 1544 18275
rect 1492 18232 1544 18241
rect 2872 18232 2924 18284
rect 2964 18207 3016 18216
rect 2964 18173 2973 18207
rect 2973 18173 3007 18207
rect 3007 18173 3016 18207
rect 2964 18164 3016 18173
rect 3148 18207 3200 18216
rect 3148 18173 3157 18207
rect 3157 18173 3191 18207
rect 3191 18173 3200 18207
rect 6460 18300 6512 18352
rect 3148 18164 3200 18173
rect 3884 18164 3936 18216
rect 4712 18164 4764 18216
rect 5264 18232 5316 18284
rect 6368 18275 6420 18284
rect 6368 18241 6377 18275
rect 6377 18241 6411 18275
rect 6411 18241 6420 18275
rect 6368 18232 6420 18241
rect 8668 18368 8720 18420
rect 12440 18411 12492 18420
rect 12440 18377 12449 18411
rect 12449 18377 12483 18411
rect 12483 18377 12492 18411
rect 12440 18368 12492 18377
rect 12532 18411 12584 18420
rect 12532 18377 12541 18411
rect 12541 18377 12575 18411
rect 12575 18377 12584 18411
rect 12532 18368 12584 18377
rect 12716 18368 12768 18420
rect 7564 18232 7616 18284
rect 9220 18275 9272 18284
rect 9220 18241 9229 18275
rect 9229 18241 9263 18275
rect 9263 18241 9272 18275
rect 9220 18232 9272 18241
rect 9772 18300 9824 18352
rect 9680 18232 9732 18284
rect 9864 18275 9916 18284
rect 9864 18241 9873 18275
rect 9873 18241 9907 18275
rect 9907 18241 9916 18275
rect 9864 18232 9916 18241
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 3424 18071 3476 18080
rect 3424 18037 3433 18071
rect 3433 18037 3467 18071
rect 3467 18037 3476 18071
rect 3424 18028 3476 18037
rect 7656 18164 7708 18216
rect 11796 18232 11848 18284
rect 12532 18232 12584 18284
rect 13176 18300 13228 18352
rect 13912 18300 13964 18352
rect 12716 18275 12768 18284
rect 12716 18241 12725 18275
rect 12725 18241 12759 18275
rect 12759 18241 12768 18275
rect 12716 18232 12768 18241
rect 12992 18232 13044 18284
rect 14188 18232 14240 18284
rect 15936 18411 15988 18420
rect 15936 18377 15945 18411
rect 15945 18377 15979 18411
rect 15979 18377 15988 18411
rect 15936 18368 15988 18377
rect 15660 18300 15712 18352
rect 17040 18368 17092 18420
rect 15108 18232 15160 18284
rect 15844 18232 15896 18284
rect 16120 18275 16172 18284
rect 16120 18241 16129 18275
rect 16129 18241 16163 18275
rect 16163 18241 16172 18275
rect 16120 18232 16172 18241
rect 10048 18207 10100 18216
rect 10048 18173 10057 18207
rect 10057 18173 10091 18207
rect 10091 18173 10100 18207
rect 10048 18164 10100 18173
rect 12256 18207 12308 18216
rect 12256 18173 12265 18207
rect 12265 18173 12299 18207
rect 12299 18173 12308 18207
rect 12256 18164 12308 18173
rect 12900 18164 12952 18216
rect 9680 18096 9732 18148
rect 11796 18096 11848 18148
rect 7012 18028 7064 18080
rect 9496 18028 9548 18080
rect 11980 18071 12032 18080
rect 11980 18037 11989 18071
rect 11989 18037 12023 18071
rect 12023 18037 12032 18071
rect 11980 18028 12032 18037
rect 14096 18071 14148 18080
rect 14096 18037 14105 18071
rect 14105 18037 14139 18071
rect 14139 18037 14148 18071
rect 14096 18028 14148 18037
rect 14464 18071 14516 18080
rect 14464 18037 14473 18071
rect 14473 18037 14507 18071
rect 14507 18037 14516 18071
rect 14464 18028 14516 18037
rect 16396 18164 16448 18216
rect 17684 18164 17736 18216
rect 18144 18164 18196 18216
rect 17592 18096 17644 18148
rect 16856 18028 16908 18080
rect 20352 18232 20404 18284
rect 19248 18207 19300 18216
rect 19248 18173 19257 18207
rect 19257 18173 19291 18207
rect 19291 18173 19300 18207
rect 19248 18164 19300 18173
rect 20720 18411 20772 18420
rect 20720 18377 20729 18411
rect 20729 18377 20763 18411
rect 20763 18377 20772 18411
rect 20720 18368 20772 18377
rect 21364 18368 21416 18420
rect 22560 18368 22612 18420
rect 20628 18300 20680 18352
rect 22008 18232 22060 18284
rect 22468 18096 22520 18148
rect 19708 18028 19760 18080
rect 22284 18071 22336 18080
rect 22284 18037 22293 18071
rect 22293 18037 22327 18071
rect 22327 18037 22336 18071
rect 22284 18028 22336 18037
rect 23020 18028 23072 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 2964 17824 3016 17876
rect 9588 17824 9640 17876
rect 12164 17867 12216 17876
rect 12164 17833 12173 17867
rect 12173 17833 12207 17867
rect 12207 17833 12216 17867
rect 12164 17824 12216 17833
rect 12256 17867 12308 17876
rect 12256 17833 12265 17867
rect 12265 17833 12299 17867
rect 12299 17833 12308 17867
rect 12256 17824 12308 17833
rect 12532 17824 12584 17876
rect 13452 17824 13504 17876
rect 16580 17824 16632 17876
rect 18052 17824 18104 17876
rect 3148 17756 3200 17808
rect 14464 17756 14516 17808
rect 1952 17731 2004 17740
rect 1952 17697 1961 17731
rect 1961 17697 1995 17731
rect 1995 17697 2004 17731
rect 1952 17688 2004 17697
rect 2412 17688 2464 17740
rect 1584 17663 1636 17672
rect 1584 17629 1593 17663
rect 1593 17629 1627 17663
rect 1627 17629 1636 17663
rect 1584 17620 1636 17629
rect 2596 17620 2648 17672
rect 8300 17731 8352 17740
rect 8300 17697 8309 17731
rect 8309 17697 8343 17731
rect 8343 17697 8352 17731
rect 8300 17688 8352 17697
rect 10048 17731 10100 17740
rect 10048 17697 10057 17731
rect 10057 17697 10091 17731
rect 10091 17697 10100 17731
rect 10048 17688 10100 17697
rect 12808 17688 12860 17740
rect 14648 17731 14700 17740
rect 14648 17697 14657 17731
rect 14657 17697 14691 17731
rect 14691 17697 14700 17731
rect 15200 17756 15252 17808
rect 14648 17688 14700 17697
rect 7564 17663 7616 17672
rect 7564 17629 7573 17663
rect 7573 17629 7607 17663
rect 7607 17629 7616 17663
rect 7564 17620 7616 17629
rect 7656 17663 7708 17672
rect 7656 17629 7665 17663
rect 7665 17629 7699 17663
rect 7699 17629 7708 17663
rect 7656 17620 7708 17629
rect 8852 17620 8904 17672
rect 9496 17620 9548 17672
rect 9864 17663 9916 17672
rect 9864 17629 9873 17663
rect 9873 17629 9907 17663
rect 9907 17629 9916 17663
rect 9864 17620 9916 17629
rect 14188 17620 14240 17672
rect 14832 17663 14884 17672
rect 14832 17629 14841 17663
rect 14841 17629 14875 17663
rect 14875 17629 14884 17663
rect 14832 17620 14884 17629
rect 15108 17663 15160 17672
rect 15108 17629 15117 17663
rect 15117 17629 15151 17663
rect 15151 17629 15160 17663
rect 15108 17620 15160 17629
rect 15384 17620 15436 17672
rect 15752 17663 15804 17672
rect 15752 17629 15761 17663
rect 15761 17629 15795 17663
rect 15795 17629 15804 17663
rect 15752 17620 15804 17629
rect 16120 17756 16172 17808
rect 16396 17756 16448 17808
rect 2964 17552 3016 17604
rect 10600 17527 10652 17536
rect 10600 17493 10609 17527
rect 10609 17493 10643 17527
rect 10643 17493 10652 17527
rect 10600 17484 10652 17493
rect 11796 17484 11848 17536
rect 12072 17484 12124 17536
rect 12532 17552 12584 17604
rect 15660 17552 15712 17604
rect 16304 17663 16356 17672
rect 16304 17629 16313 17663
rect 16313 17629 16347 17663
rect 16347 17629 16356 17663
rect 16304 17620 16356 17629
rect 16580 17663 16632 17672
rect 16580 17629 16589 17663
rect 16589 17629 16623 17663
rect 16623 17629 16632 17663
rect 16580 17620 16632 17629
rect 17408 17688 17460 17740
rect 17500 17731 17552 17740
rect 17500 17697 17509 17731
rect 17509 17697 17543 17731
rect 17543 17697 17552 17731
rect 17500 17688 17552 17697
rect 19800 17756 19852 17808
rect 20996 17756 21048 17808
rect 17960 17688 18012 17740
rect 16856 17663 16908 17672
rect 16856 17629 16865 17663
rect 16865 17629 16899 17663
rect 16899 17629 16908 17663
rect 16856 17620 16908 17629
rect 17592 17620 17644 17672
rect 17684 17663 17736 17672
rect 17684 17629 17693 17663
rect 17693 17629 17727 17663
rect 17727 17629 17736 17663
rect 17684 17620 17736 17629
rect 18052 17663 18104 17672
rect 18052 17629 18061 17663
rect 18061 17629 18095 17663
rect 18095 17629 18104 17663
rect 18052 17620 18104 17629
rect 18236 17688 18288 17740
rect 18328 17663 18380 17672
rect 18328 17629 18337 17663
rect 18337 17629 18371 17663
rect 18371 17629 18380 17663
rect 18328 17620 18380 17629
rect 18696 17620 18748 17672
rect 19156 17688 19208 17740
rect 19340 17620 19392 17672
rect 20720 17663 20772 17672
rect 20720 17629 20729 17663
rect 20729 17629 20763 17663
rect 20763 17629 20772 17663
rect 20720 17620 20772 17629
rect 20904 17663 20956 17672
rect 20904 17629 20913 17663
rect 20913 17629 20947 17663
rect 20947 17629 20956 17663
rect 20904 17620 20956 17629
rect 20996 17663 21048 17672
rect 20996 17629 21005 17663
rect 21005 17629 21039 17663
rect 21039 17629 21048 17663
rect 20996 17620 21048 17629
rect 12348 17484 12400 17536
rect 15016 17527 15068 17536
rect 15016 17493 15025 17527
rect 15025 17493 15059 17527
rect 15059 17493 15068 17527
rect 15016 17484 15068 17493
rect 15844 17484 15896 17536
rect 16396 17484 16448 17536
rect 17684 17484 17736 17536
rect 18972 17484 19024 17536
rect 19340 17484 19392 17536
rect 21272 17663 21324 17672
rect 21272 17629 21281 17663
rect 21281 17629 21315 17663
rect 21315 17629 21324 17663
rect 21272 17620 21324 17629
rect 21916 17620 21968 17672
rect 22468 17731 22520 17740
rect 22468 17697 22477 17731
rect 22477 17697 22511 17731
rect 22511 17697 22520 17731
rect 22468 17688 22520 17697
rect 24492 17688 24544 17740
rect 24032 17552 24084 17604
rect 22284 17484 22336 17536
rect 22468 17484 22520 17536
rect 24216 17527 24268 17536
rect 24216 17493 24225 17527
rect 24225 17493 24259 17527
rect 24259 17493 24268 17527
rect 24216 17484 24268 17493
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 2412 17323 2464 17332
rect 2412 17289 2421 17323
rect 2421 17289 2455 17323
rect 2455 17289 2464 17323
rect 2412 17280 2464 17289
rect 4068 17280 4120 17332
rect 1860 17187 1912 17196
rect 1860 17153 1869 17187
rect 1869 17153 1903 17187
rect 1903 17153 1912 17187
rect 1860 17144 1912 17153
rect 3424 17144 3476 17196
rect 4068 17144 4120 17196
rect 8300 17280 8352 17332
rect 10048 17280 10100 17332
rect 13268 17212 13320 17264
rect 15476 17212 15528 17264
rect 7564 17187 7616 17196
rect 7564 17153 7573 17187
rect 7573 17153 7607 17187
rect 7607 17153 7616 17187
rect 7564 17144 7616 17153
rect 7840 17187 7892 17196
rect 7840 17153 7849 17187
rect 7849 17153 7883 17187
rect 7883 17153 7892 17187
rect 7840 17144 7892 17153
rect 8668 17144 8720 17196
rect 9680 17187 9732 17196
rect 9680 17153 9689 17187
rect 9689 17153 9723 17187
rect 9723 17153 9732 17187
rect 9680 17144 9732 17153
rect 9772 17144 9824 17196
rect 11612 17144 11664 17196
rect 1952 17119 2004 17128
rect 1952 17085 1961 17119
rect 1961 17085 1995 17119
rect 1995 17085 2004 17119
rect 1952 17076 2004 17085
rect 2688 17008 2740 17060
rect 8852 17119 8904 17128
rect 8852 17085 8861 17119
rect 8861 17085 8895 17119
rect 8895 17085 8904 17119
rect 8852 17076 8904 17085
rect 8944 17119 8996 17128
rect 8944 17085 8953 17119
rect 8953 17085 8987 17119
rect 8987 17085 8996 17119
rect 8944 17076 8996 17085
rect 4620 17008 4672 17060
rect 12716 17076 12768 17128
rect 13820 17187 13872 17196
rect 13820 17153 13829 17187
rect 13829 17153 13863 17187
rect 13863 17153 13872 17187
rect 13820 17144 13872 17153
rect 14372 17144 14424 17196
rect 14464 17187 14516 17196
rect 14464 17153 14473 17187
rect 14473 17153 14507 17187
rect 14507 17153 14516 17187
rect 14464 17144 14516 17153
rect 14648 17144 14700 17196
rect 10232 17008 10284 17060
rect 13268 17008 13320 17060
rect 4712 16983 4764 16992
rect 4712 16949 4721 16983
rect 4721 16949 4755 16983
rect 4755 16949 4764 16983
rect 4712 16940 4764 16949
rect 12624 16940 12676 16992
rect 14004 16940 14056 16992
rect 14372 16983 14424 16992
rect 14372 16949 14381 16983
rect 14381 16949 14415 16983
rect 14415 16949 14424 16983
rect 14372 16940 14424 16949
rect 14556 17008 14608 17060
rect 15752 17280 15804 17332
rect 18052 17280 18104 17332
rect 18696 17280 18748 17332
rect 20812 17280 20864 17332
rect 20904 17280 20956 17332
rect 15660 17187 15712 17196
rect 15660 17153 15669 17187
rect 15669 17153 15703 17187
rect 15703 17153 15712 17187
rect 15660 17144 15712 17153
rect 15752 17187 15804 17196
rect 15752 17153 15761 17187
rect 15761 17153 15795 17187
rect 15795 17153 15804 17187
rect 15752 17144 15804 17153
rect 16028 17144 16080 17196
rect 20996 17212 21048 17264
rect 16856 17187 16908 17196
rect 16856 17153 16865 17187
rect 16865 17153 16899 17187
rect 16899 17153 16908 17187
rect 16856 17144 16908 17153
rect 17132 17144 17184 17196
rect 18328 17144 18380 17196
rect 19064 17144 19116 17196
rect 19340 17187 19392 17196
rect 19340 17153 19349 17187
rect 19349 17153 19383 17187
rect 19383 17153 19392 17187
rect 19340 17144 19392 17153
rect 19892 17144 19944 17196
rect 21272 17187 21324 17196
rect 21272 17153 21281 17187
rect 21281 17153 21315 17187
rect 21315 17153 21324 17187
rect 21272 17144 21324 17153
rect 17408 17008 17460 17060
rect 17960 17008 18012 17060
rect 19800 17119 19852 17128
rect 19800 17085 19809 17119
rect 19809 17085 19843 17119
rect 19843 17085 19852 17119
rect 19800 17076 19852 17085
rect 20168 17076 20220 17128
rect 21732 17144 21784 17196
rect 23480 17187 23532 17196
rect 23480 17153 23489 17187
rect 23489 17153 23523 17187
rect 23523 17153 23532 17187
rect 23480 17144 23532 17153
rect 24216 17144 24268 17196
rect 25228 17187 25280 17196
rect 25228 17153 25237 17187
rect 25237 17153 25271 17187
rect 25271 17153 25280 17187
rect 25228 17144 25280 17153
rect 24860 17076 24912 17128
rect 22744 17008 22796 17060
rect 14832 16940 14884 16992
rect 16304 16940 16356 16992
rect 18052 16940 18104 16992
rect 19156 16940 19208 16992
rect 20904 16940 20956 16992
rect 20996 16940 21048 16992
rect 23112 16940 23164 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 8668 16736 8720 16788
rect 8392 16668 8444 16720
rect 2964 16643 3016 16652
rect 2964 16609 2973 16643
rect 2973 16609 3007 16643
rect 3007 16609 3016 16643
rect 2964 16600 3016 16609
rect 3516 16643 3568 16652
rect 3516 16609 3525 16643
rect 3525 16609 3559 16643
rect 3559 16609 3568 16643
rect 3516 16600 3568 16609
rect 8116 16643 8168 16652
rect 8116 16609 8125 16643
rect 8125 16609 8159 16643
rect 8159 16609 8168 16643
rect 8116 16600 8168 16609
rect 9312 16643 9364 16652
rect 9312 16609 9321 16643
rect 9321 16609 9355 16643
rect 9355 16609 9364 16643
rect 9312 16600 9364 16609
rect 2872 16575 2924 16584
rect 2872 16541 2881 16575
rect 2881 16541 2915 16575
rect 2915 16541 2924 16575
rect 2872 16532 2924 16541
rect 5724 16532 5776 16584
rect 7380 16575 7432 16584
rect 7380 16541 7389 16575
rect 7389 16541 7423 16575
rect 7423 16541 7432 16575
rect 7380 16532 7432 16541
rect 7472 16532 7524 16584
rect 8576 16532 8628 16584
rect 8944 16532 8996 16584
rect 12348 16736 12400 16788
rect 15384 16736 15436 16788
rect 16028 16779 16080 16788
rect 16028 16745 16037 16779
rect 16037 16745 16071 16779
rect 16071 16745 16080 16779
rect 16028 16736 16080 16745
rect 16120 16736 16172 16788
rect 20720 16736 20772 16788
rect 20812 16736 20864 16788
rect 23112 16779 23164 16788
rect 23112 16745 23121 16779
rect 23121 16745 23155 16779
rect 23155 16745 23164 16779
rect 23112 16736 23164 16745
rect 11612 16668 11664 16720
rect 11980 16600 12032 16652
rect 12716 16600 12768 16652
rect 10232 16575 10284 16584
rect 10232 16541 10241 16575
rect 10241 16541 10275 16575
rect 10275 16541 10284 16575
rect 10232 16532 10284 16541
rect 4804 16464 4856 16516
rect 9496 16464 9548 16516
rect 11888 16532 11940 16584
rect 12256 16575 12308 16584
rect 12256 16541 12265 16575
rect 12265 16541 12299 16575
rect 12299 16541 12308 16575
rect 12256 16532 12308 16541
rect 12532 16532 12584 16584
rect 12624 16575 12676 16584
rect 12624 16541 12633 16575
rect 12633 16541 12667 16575
rect 12667 16541 12676 16575
rect 12624 16532 12676 16541
rect 12164 16464 12216 16516
rect 13176 16575 13228 16584
rect 13176 16541 13185 16575
rect 13185 16541 13219 16575
rect 13219 16541 13228 16575
rect 13176 16532 13228 16541
rect 16028 16532 16080 16584
rect 17040 16532 17092 16584
rect 20168 16600 20220 16652
rect 20904 16643 20956 16652
rect 20904 16609 20909 16643
rect 20909 16609 20943 16643
rect 20943 16609 20956 16643
rect 20904 16600 20956 16609
rect 21088 16643 21140 16652
rect 21088 16609 21097 16643
rect 21097 16609 21131 16643
rect 21131 16609 21140 16643
rect 21088 16600 21140 16609
rect 21732 16643 21784 16652
rect 21732 16609 21741 16643
rect 21741 16609 21775 16643
rect 21775 16609 21784 16643
rect 21732 16600 21784 16609
rect 20444 16532 20496 16584
rect 21640 16575 21692 16584
rect 13360 16439 13412 16448
rect 13360 16405 13369 16439
rect 13369 16405 13403 16439
rect 13403 16405 13412 16439
rect 13360 16396 13412 16405
rect 14372 16507 14424 16516
rect 14372 16473 14381 16507
rect 14381 16473 14415 16507
rect 14415 16473 14424 16507
rect 14372 16464 14424 16473
rect 15660 16464 15712 16516
rect 19524 16464 19576 16516
rect 14556 16396 14608 16448
rect 15108 16396 15160 16448
rect 19800 16396 19852 16448
rect 20168 16507 20220 16516
rect 20168 16473 20177 16507
rect 20177 16473 20211 16507
rect 20211 16473 20220 16507
rect 21640 16541 21649 16575
rect 21649 16541 21683 16575
rect 21683 16541 21692 16575
rect 21640 16532 21692 16541
rect 24032 16668 24084 16720
rect 20168 16464 20220 16473
rect 21456 16464 21508 16516
rect 22652 16532 22704 16584
rect 22836 16575 22888 16584
rect 22836 16541 22845 16575
rect 22845 16541 22879 16575
rect 22879 16541 22888 16575
rect 22836 16532 22888 16541
rect 22928 16532 22980 16584
rect 23572 16575 23624 16584
rect 23572 16541 23581 16575
rect 23581 16541 23615 16575
rect 23615 16541 23624 16575
rect 23572 16532 23624 16541
rect 23848 16575 23900 16584
rect 23848 16541 23857 16575
rect 23857 16541 23891 16575
rect 23891 16541 23900 16575
rect 23848 16532 23900 16541
rect 24492 16532 24544 16584
rect 24860 16464 24912 16516
rect 19984 16396 20036 16448
rect 20904 16439 20956 16448
rect 20904 16405 20913 16439
rect 20913 16405 20947 16439
rect 20947 16405 20956 16439
rect 20904 16396 20956 16405
rect 20996 16396 21048 16448
rect 22284 16439 22336 16448
rect 22284 16405 22293 16439
rect 22293 16405 22327 16439
rect 22327 16405 22336 16439
rect 22284 16396 22336 16405
rect 23204 16396 23256 16448
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 2872 16192 2924 16244
rect 7564 16192 7616 16244
rect 10232 16192 10284 16244
rect 13176 16192 13228 16244
rect 14096 16192 14148 16244
rect 848 16056 900 16108
rect 1860 15988 1912 16040
rect 3148 16099 3200 16108
rect 3148 16065 3157 16099
rect 3157 16065 3191 16099
rect 3191 16065 3200 16099
rect 3148 16056 3200 16065
rect 3884 16099 3936 16108
rect 3884 16065 3893 16099
rect 3893 16065 3927 16099
rect 3927 16065 3936 16099
rect 3884 16056 3936 16065
rect 3976 15988 4028 16040
rect 4620 16099 4672 16108
rect 4620 16065 4629 16099
rect 4629 16065 4663 16099
rect 4663 16065 4672 16099
rect 4620 16056 4672 16065
rect 4712 16056 4764 16108
rect 5724 16056 5776 16108
rect 4804 16031 4856 16040
rect 4804 15997 4813 16031
rect 4813 15997 4847 16031
rect 4847 15997 4856 16031
rect 4804 15988 4856 15997
rect 7196 16099 7248 16108
rect 7196 16065 7205 16099
rect 7205 16065 7239 16099
rect 7239 16065 7248 16099
rect 7196 16056 7248 16065
rect 7840 16056 7892 16108
rect 8300 16099 8352 16108
rect 8300 16065 8309 16099
rect 8309 16065 8343 16099
rect 8343 16065 8352 16099
rect 8300 16056 8352 16065
rect 9588 16099 9640 16108
rect 9588 16065 9597 16099
rect 9597 16065 9631 16099
rect 9631 16065 9640 16099
rect 9588 16056 9640 16065
rect 9864 16056 9916 16108
rect 11796 16124 11848 16176
rect 10048 16031 10100 16040
rect 10048 15997 10057 16031
rect 10057 15997 10091 16031
rect 10091 15997 10100 16031
rect 10048 15988 10100 15997
rect 7288 15920 7340 15972
rect 11704 16056 11756 16108
rect 12716 16124 12768 16176
rect 15108 16192 15160 16244
rect 17132 16235 17184 16244
rect 17132 16201 17141 16235
rect 17141 16201 17175 16235
rect 17175 16201 17184 16235
rect 17132 16192 17184 16201
rect 17224 16192 17276 16244
rect 17868 16192 17920 16244
rect 18052 16192 18104 16244
rect 18880 16192 18932 16244
rect 19616 16235 19668 16244
rect 19616 16201 19625 16235
rect 19625 16201 19659 16235
rect 19659 16201 19668 16235
rect 19616 16192 19668 16201
rect 20168 16192 20220 16244
rect 23204 16235 23256 16244
rect 23204 16201 23213 16235
rect 23213 16201 23247 16235
rect 23247 16201 23256 16235
rect 23204 16192 23256 16201
rect 24032 16192 24084 16244
rect 13820 16056 13872 16108
rect 10600 15988 10652 16040
rect 14464 16056 14516 16108
rect 15016 16056 15068 16108
rect 17224 16056 17276 16108
rect 17408 16099 17460 16108
rect 17408 16065 17417 16099
rect 17417 16065 17451 16099
rect 17451 16065 17460 16099
rect 17408 16056 17460 16065
rect 15200 15988 15252 16040
rect 17776 15988 17828 16040
rect 14004 15920 14056 15972
rect 16948 15920 17000 15972
rect 17132 15920 17184 15972
rect 18052 16099 18104 16108
rect 18052 16065 18061 16099
rect 18061 16065 18095 16099
rect 18095 16065 18104 16099
rect 18052 16056 18104 16065
rect 18880 16099 18932 16108
rect 18880 16065 18889 16099
rect 18889 16065 18923 16099
rect 18923 16065 18932 16099
rect 18880 16056 18932 16065
rect 19892 16124 19944 16176
rect 22284 16124 22336 16176
rect 20904 16056 20956 16108
rect 19340 15920 19392 15972
rect 3792 15895 3844 15904
rect 3792 15861 3801 15895
rect 3801 15861 3835 15895
rect 3835 15861 3844 15895
rect 3792 15852 3844 15861
rect 4620 15852 4672 15904
rect 5724 15895 5776 15904
rect 5724 15861 5733 15895
rect 5733 15861 5767 15895
rect 5767 15861 5776 15895
rect 5724 15852 5776 15861
rect 8116 15852 8168 15904
rect 9312 15895 9364 15904
rect 9312 15861 9321 15895
rect 9321 15861 9355 15895
rect 9355 15861 9364 15895
rect 9312 15852 9364 15861
rect 9680 15895 9732 15904
rect 9680 15861 9689 15895
rect 9689 15861 9723 15895
rect 9723 15861 9732 15895
rect 9680 15852 9732 15861
rect 13820 15895 13872 15904
rect 13820 15861 13829 15895
rect 13829 15861 13863 15895
rect 13863 15861 13872 15895
rect 13820 15852 13872 15861
rect 14096 15895 14148 15904
rect 14096 15861 14105 15895
rect 14105 15861 14139 15895
rect 14139 15861 14148 15895
rect 14096 15852 14148 15861
rect 14280 15895 14332 15904
rect 14280 15861 14289 15895
rect 14289 15861 14323 15895
rect 14323 15861 14332 15895
rect 14280 15852 14332 15861
rect 15108 15895 15160 15904
rect 15108 15861 15117 15895
rect 15117 15861 15151 15895
rect 15151 15861 15160 15895
rect 15108 15852 15160 15861
rect 16672 15895 16724 15904
rect 16672 15861 16681 15895
rect 16681 15861 16715 15895
rect 16715 15861 16724 15895
rect 16672 15852 16724 15861
rect 17224 15852 17276 15904
rect 17408 15852 17460 15904
rect 20444 15988 20496 16040
rect 21088 15988 21140 16040
rect 21640 15988 21692 16040
rect 23388 16099 23440 16108
rect 23388 16065 23397 16099
rect 23397 16065 23431 16099
rect 23431 16065 23440 16099
rect 23388 16056 23440 16065
rect 23756 15988 23808 16040
rect 20260 15852 20312 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 12164 15691 12216 15700
rect 12164 15657 12173 15691
rect 12173 15657 12207 15691
rect 12207 15657 12216 15691
rect 12164 15648 12216 15657
rect 13820 15648 13872 15700
rect 16856 15648 16908 15700
rect 18696 15648 18748 15700
rect 22836 15648 22888 15700
rect 23572 15648 23624 15700
rect 24768 15648 24820 15700
rect 16948 15580 17000 15632
rect 4620 15512 4672 15564
rect 13360 15512 13412 15564
rect 3792 15444 3844 15496
rect 7288 15487 7340 15496
rect 7288 15453 7297 15487
rect 7297 15453 7331 15487
rect 7331 15453 7340 15487
rect 7288 15444 7340 15453
rect 8116 15487 8168 15496
rect 8116 15453 8125 15487
rect 8125 15453 8159 15487
rect 8159 15453 8168 15487
rect 8116 15444 8168 15453
rect 9312 15487 9364 15496
rect 9312 15453 9321 15487
rect 9321 15453 9355 15487
rect 9355 15453 9364 15487
rect 9312 15444 9364 15453
rect 9680 15444 9732 15496
rect 10508 15444 10560 15496
rect 9864 15376 9916 15428
rect 11704 15444 11756 15496
rect 11796 15487 11848 15496
rect 11796 15453 11805 15487
rect 11805 15453 11839 15487
rect 11839 15453 11848 15487
rect 11796 15444 11848 15453
rect 11980 15487 12032 15496
rect 11980 15453 11989 15487
rect 11989 15453 12023 15487
rect 12023 15453 12032 15487
rect 11980 15444 12032 15453
rect 16580 15444 16632 15496
rect 16764 15487 16816 15496
rect 16764 15453 16773 15487
rect 16773 15453 16807 15487
rect 16807 15453 16816 15487
rect 16764 15444 16816 15453
rect 17040 15555 17092 15564
rect 17040 15521 17049 15555
rect 17049 15521 17083 15555
rect 17083 15521 17092 15555
rect 17040 15512 17092 15521
rect 19616 15580 19668 15632
rect 23204 15580 23256 15632
rect 23480 15623 23532 15632
rect 23480 15589 23489 15623
rect 23489 15589 23523 15623
rect 23523 15589 23532 15623
rect 23480 15580 23532 15589
rect 20260 15555 20312 15564
rect 20260 15521 20269 15555
rect 20269 15521 20303 15555
rect 20303 15521 20312 15555
rect 20260 15512 20312 15521
rect 20720 15512 20772 15564
rect 19984 15487 20036 15496
rect 19984 15453 19993 15487
rect 19993 15453 20027 15487
rect 20027 15453 20036 15487
rect 19984 15444 20036 15453
rect 20812 15444 20864 15496
rect 21456 15512 21508 15564
rect 21640 15444 21692 15496
rect 4712 15351 4764 15360
rect 4712 15317 4721 15351
rect 4721 15317 4755 15351
rect 4755 15317 4764 15351
rect 4712 15308 4764 15317
rect 19524 15376 19576 15428
rect 20352 15376 20404 15428
rect 24860 15512 24912 15564
rect 23112 15444 23164 15496
rect 23572 15487 23624 15496
rect 23572 15453 23581 15487
rect 23581 15453 23615 15487
rect 23615 15453 23624 15487
rect 23572 15444 23624 15453
rect 24216 15444 24268 15496
rect 23756 15376 23808 15428
rect 16028 15308 16080 15360
rect 16764 15308 16816 15360
rect 19800 15351 19852 15360
rect 19800 15317 19809 15351
rect 19809 15317 19843 15351
rect 19843 15317 19852 15351
rect 19800 15308 19852 15317
rect 21088 15351 21140 15360
rect 21088 15317 21097 15351
rect 21097 15317 21131 15351
rect 21131 15317 21140 15351
rect 21088 15308 21140 15317
rect 24032 15308 24084 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 7288 15104 7340 15156
rect 2412 14968 2464 15020
rect 2688 15011 2740 15020
rect 2688 14977 2697 15011
rect 2697 14977 2731 15011
rect 2731 14977 2740 15011
rect 2688 14968 2740 14977
rect 3332 14968 3384 15020
rect 3516 15011 3568 15020
rect 3516 14977 3525 15011
rect 3525 14977 3559 15011
rect 3559 14977 3568 15011
rect 8116 15036 8168 15088
rect 9588 15104 9640 15156
rect 12072 15104 12124 15156
rect 12348 15147 12400 15156
rect 12348 15113 12357 15147
rect 12357 15113 12391 15147
rect 12391 15113 12400 15147
rect 12348 15104 12400 15113
rect 14280 15104 14332 15156
rect 16764 15104 16816 15156
rect 16948 15104 17000 15156
rect 20812 15147 20864 15156
rect 20812 15113 20821 15147
rect 20821 15113 20855 15147
rect 20855 15113 20864 15147
rect 20812 15104 20864 15113
rect 23388 15147 23440 15156
rect 23388 15113 23397 15147
rect 23397 15113 23431 15147
rect 23431 15113 23440 15147
rect 23388 15104 23440 15113
rect 23848 15104 23900 15156
rect 10692 15036 10744 15088
rect 3516 14968 3568 14977
rect 4712 14968 4764 15020
rect 5264 15011 5316 15020
rect 5264 14977 5273 15011
rect 5273 14977 5307 15011
rect 5307 14977 5316 15011
rect 5264 14968 5316 14977
rect 5724 14968 5776 15020
rect 7380 14968 7432 15020
rect 7472 15011 7524 15020
rect 7472 14977 7481 15011
rect 7481 14977 7515 15011
rect 7515 14977 7524 15011
rect 7472 14968 7524 14977
rect 8668 15011 8720 15020
rect 8668 14977 8677 15011
rect 8677 14977 8711 15011
rect 8711 14977 8720 15011
rect 8668 14968 8720 14977
rect 4068 14943 4120 14952
rect 4068 14909 4077 14943
rect 4077 14909 4111 14943
rect 4111 14909 4120 14943
rect 4068 14900 4120 14909
rect 6828 14900 6880 14952
rect 7196 14832 7248 14884
rect 8576 14900 8628 14952
rect 9864 15011 9916 15020
rect 9864 14977 9873 15011
rect 9873 14977 9907 15011
rect 9907 14977 9916 15011
rect 9864 14968 9916 14977
rect 10048 14968 10100 15020
rect 11796 15011 11848 15020
rect 11796 14977 11805 15011
rect 11805 14977 11839 15011
rect 11839 14977 11848 15011
rect 11796 14968 11848 14977
rect 7932 14832 7984 14884
rect 10508 14832 10560 14884
rect 12072 15011 12124 15020
rect 12072 14977 12081 15011
rect 12081 14977 12115 15011
rect 12115 14977 12124 15011
rect 12072 14968 12124 14977
rect 12072 14832 12124 14884
rect 2872 14764 2924 14816
rect 3884 14764 3936 14816
rect 11336 14764 11388 14816
rect 12440 14968 12492 15020
rect 14372 15036 14424 15088
rect 12900 15011 12952 15020
rect 12900 14977 12909 15011
rect 12909 14977 12943 15011
rect 12943 14977 12952 15011
rect 12900 14968 12952 14977
rect 13360 14968 13412 15020
rect 14280 15011 14332 15020
rect 14280 14977 14289 15011
rect 14289 14977 14323 15011
rect 14323 14977 14332 15011
rect 14280 14968 14332 14977
rect 14832 14968 14884 15020
rect 17040 15011 17092 15020
rect 17040 14977 17049 15011
rect 17049 14977 17083 15011
rect 17083 14977 17092 15011
rect 17040 14968 17092 14977
rect 18052 15036 18104 15088
rect 20628 15036 20680 15088
rect 22192 15036 22244 15088
rect 23756 15079 23808 15088
rect 23756 15045 23765 15079
rect 23765 15045 23799 15079
rect 23799 15045 23808 15079
rect 23756 15036 23808 15045
rect 14188 14943 14240 14952
rect 14188 14909 14197 14943
rect 14197 14909 14231 14943
rect 14231 14909 14240 14943
rect 14188 14900 14240 14909
rect 14464 14900 14516 14952
rect 14740 14900 14792 14952
rect 15016 14900 15068 14952
rect 15292 14900 15344 14952
rect 17408 14900 17460 14952
rect 17776 14943 17828 14952
rect 17776 14909 17785 14943
rect 17785 14909 17819 14943
rect 17819 14909 17828 14943
rect 17776 14900 17828 14909
rect 18144 15011 18196 15020
rect 18144 14977 18153 15011
rect 18153 14977 18187 15011
rect 18187 14977 18196 15011
rect 18144 14968 18196 14977
rect 19984 15011 20036 15020
rect 19984 14977 19993 15011
rect 19993 14977 20027 15011
rect 20027 14977 20036 15011
rect 19984 14968 20036 14977
rect 20260 15011 20312 15020
rect 20260 14977 20269 15011
rect 20269 14977 20303 15011
rect 20303 14977 20312 15011
rect 20260 14968 20312 14977
rect 20904 14968 20956 15020
rect 20996 15011 21048 15020
rect 20996 14977 21005 15011
rect 21005 14977 21039 15011
rect 21039 14977 21048 15011
rect 20996 14968 21048 14977
rect 21088 14968 21140 15020
rect 21456 15011 21508 15020
rect 21456 14977 21465 15011
rect 21465 14977 21499 15011
rect 21499 14977 21508 15011
rect 21456 14968 21508 14977
rect 21640 15011 21692 15020
rect 21640 14977 21649 15011
rect 21649 14977 21683 15011
rect 21683 14977 21692 15011
rect 21640 14968 21692 14977
rect 22376 14968 22428 15020
rect 23940 15011 23992 15020
rect 23940 14977 23949 15011
rect 23949 14977 23983 15011
rect 23983 14977 23992 15011
rect 23940 14968 23992 14977
rect 24032 15011 24084 15020
rect 24032 14977 24041 15011
rect 24041 14977 24075 15011
rect 24075 14977 24084 15011
rect 24032 14968 24084 14977
rect 17592 14832 17644 14884
rect 20628 14900 20680 14952
rect 20720 14900 20772 14952
rect 24216 14900 24268 14952
rect 18788 14832 18840 14884
rect 12256 14764 12308 14816
rect 14924 14764 14976 14816
rect 16948 14764 17000 14816
rect 17316 14807 17368 14816
rect 17316 14773 17325 14807
rect 17325 14773 17359 14807
rect 17359 14773 17368 14807
rect 17316 14764 17368 14773
rect 19708 14764 19760 14816
rect 20076 14807 20128 14816
rect 20076 14773 20085 14807
rect 20085 14773 20119 14807
rect 20119 14773 20128 14807
rect 20076 14764 20128 14773
rect 21180 14875 21232 14884
rect 21180 14841 21189 14875
rect 21189 14841 21223 14875
rect 21223 14841 21232 14875
rect 21180 14832 21232 14841
rect 21824 14832 21876 14884
rect 23296 14832 23348 14884
rect 23572 14832 23624 14884
rect 22008 14764 22060 14816
rect 23388 14764 23440 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 3332 14603 3384 14612
rect 3332 14569 3341 14603
rect 3341 14569 3375 14603
rect 3375 14569 3384 14603
rect 3332 14560 3384 14569
rect 3792 14560 3844 14612
rect 2780 14492 2832 14544
rect 2688 14424 2740 14476
rect 2872 14467 2924 14476
rect 2872 14433 2881 14467
rect 2881 14433 2915 14467
rect 2915 14433 2924 14467
rect 2872 14424 2924 14433
rect 3976 14492 4028 14544
rect 12072 14560 12124 14612
rect 14924 14560 14976 14612
rect 15292 14560 15344 14612
rect 17040 14560 17092 14612
rect 4712 14492 4764 14544
rect 7288 14492 7340 14544
rect 16856 14492 16908 14544
rect 18604 14603 18656 14612
rect 18604 14569 18613 14603
rect 18613 14569 18647 14603
rect 18647 14569 18656 14603
rect 18604 14560 18656 14569
rect 21364 14560 21416 14612
rect 22560 14560 22612 14612
rect 23112 14560 23164 14612
rect 23756 14560 23808 14612
rect 19248 14492 19300 14544
rect 19432 14535 19484 14544
rect 19432 14501 19441 14535
rect 19441 14501 19475 14535
rect 19475 14501 19484 14535
rect 19432 14492 19484 14501
rect 20628 14535 20680 14544
rect 20628 14501 20637 14535
rect 20637 14501 20671 14535
rect 20671 14501 20680 14535
rect 20628 14492 20680 14501
rect 2412 14356 2464 14408
rect 3332 14356 3384 14408
rect 3884 14399 3936 14408
rect 3884 14365 3893 14399
rect 3893 14365 3927 14399
rect 3927 14365 3936 14399
rect 3884 14356 3936 14365
rect 5264 14467 5316 14476
rect 5264 14433 5273 14467
rect 5273 14433 5307 14467
rect 5307 14433 5316 14467
rect 5264 14424 5316 14433
rect 6828 14424 6880 14476
rect 14004 14424 14056 14476
rect 14648 14424 14700 14476
rect 15384 14424 15436 14476
rect 17040 14424 17092 14476
rect 3148 14288 3200 14340
rect 3608 14288 3660 14340
rect 6736 14399 6788 14408
rect 6736 14365 6745 14399
rect 6745 14365 6779 14399
rect 6779 14365 6788 14399
rect 6736 14356 6788 14365
rect 13268 14356 13320 14408
rect 13452 14399 13504 14408
rect 13452 14365 13461 14399
rect 13461 14365 13495 14399
rect 13495 14365 13504 14399
rect 13452 14356 13504 14365
rect 11336 14331 11388 14340
rect 11336 14297 11345 14331
rect 11345 14297 11379 14331
rect 11379 14297 11388 14331
rect 11336 14288 11388 14297
rect 14556 14288 14608 14340
rect 15200 14399 15252 14408
rect 15200 14365 15209 14399
rect 15209 14365 15243 14399
rect 15243 14365 15252 14399
rect 15200 14356 15252 14365
rect 16856 14399 16908 14408
rect 16856 14365 16865 14399
rect 16865 14365 16899 14399
rect 16899 14365 16908 14399
rect 16856 14356 16908 14365
rect 17960 14424 18012 14476
rect 17224 14399 17276 14408
rect 17224 14365 17233 14399
rect 17233 14365 17267 14399
rect 17267 14365 17276 14399
rect 17224 14356 17276 14365
rect 17684 14399 17736 14408
rect 17684 14365 17693 14399
rect 17693 14365 17727 14399
rect 17727 14365 17736 14399
rect 17684 14356 17736 14365
rect 20076 14424 20128 14476
rect 20904 14467 20956 14476
rect 20904 14433 20913 14467
rect 20913 14433 20947 14467
rect 20947 14433 20956 14467
rect 20904 14424 20956 14433
rect 21180 14424 21232 14476
rect 19432 14399 19484 14408
rect 19432 14365 19441 14399
rect 19441 14365 19475 14399
rect 19475 14365 19484 14399
rect 19432 14356 19484 14365
rect 19800 14399 19852 14408
rect 19800 14365 19809 14399
rect 19809 14365 19843 14399
rect 19843 14365 19852 14399
rect 19800 14356 19852 14365
rect 20996 14399 21048 14408
rect 20996 14365 21005 14399
rect 21005 14365 21039 14399
rect 21039 14365 21048 14399
rect 23296 14492 23348 14544
rect 22100 14424 22152 14476
rect 20996 14356 21048 14365
rect 22652 14356 22704 14408
rect 23940 14492 23992 14544
rect 24768 14492 24820 14544
rect 23664 14424 23716 14476
rect 18144 14331 18196 14340
rect 18144 14297 18153 14331
rect 18153 14297 18187 14331
rect 18187 14297 18196 14331
rect 18144 14288 18196 14297
rect 19340 14288 19392 14340
rect 21824 14288 21876 14340
rect 22008 14331 22060 14340
rect 22008 14297 22017 14331
rect 22017 14297 22051 14331
rect 22051 14297 22060 14331
rect 22008 14288 22060 14297
rect 23756 14399 23808 14408
rect 23756 14365 23765 14399
rect 23765 14365 23799 14399
rect 23799 14365 23808 14399
rect 23756 14356 23808 14365
rect 23940 14399 23992 14408
rect 23940 14365 23949 14399
rect 23949 14365 23983 14399
rect 23983 14365 23992 14399
rect 23940 14356 23992 14365
rect 24216 14356 24268 14408
rect 4160 14220 4212 14272
rect 12808 14263 12860 14272
rect 12808 14229 12817 14263
rect 12817 14229 12851 14263
rect 12851 14229 12860 14263
rect 12808 14220 12860 14229
rect 12992 14263 13044 14272
rect 12992 14229 13001 14263
rect 13001 14229 13035 14263
rect 13035 14229 13044 14263
rect 12992 14220 13044 14229
rect 13360 14263 13412 14272
rect 13360 14229 13369 14263
rect 13369 14229 13403 14263
rect 13403 14229 13412 14263
rect 13360 14220 13412 14229
rect 14924 14220 14976 14272
rect 17132 14263 17184 14272
rect 17132 14229 17141 14263
rect 17141 14229 17175 14263
rect 17175 14229 17184 14263
rect 17132 14220 17184 14229
rect 19064 14220 19116 14272
rect 23388 14288 23440 14340
rect 22928 14220 22980 14272
rect 23572 14263 23624 14272
rect 23572 14229 23581 14263
rect 23581 14229 23615 14263
rect 23615 14229 23624 14263
rect 23572 14220 23624 14229
rect 24492 14331 24544 14340
rect 24492 14297 24501 14331
rect 24501 14297 24535 14331
rect 24535 14297 24544 14331
rect 24492 14288 24544 14297
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 1952 13812 2004 13864
rect 3332 14016 3384 14068
rect 3792 14016 3844 14068
rect 4068 14016 4120 14068
rect 3148 13923 3200 13932
rect 3148 13889 3157 13923
rect 3157 13889 3191 13923
rect 3191 13889 3200 13923
rect 3148 13880 3200 13889
rect 3608 13948 3660 14000
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 2780 13812 2832 13821
rect 4068 13880 4120 13932
rect 4160 13923 4212 13932
rect 4160 13889 4169 13923
rect 4169 13889 4203 13923
rect 4203 13889 4212 13923
rect 4160 13880 4212 13889
rect 7932 13948 7984 14000
rect 6736 13880 6788 13932
rect 10508 13880 10560 13932
rect 5540 13812 5592 13864
rect 6828 13812 6880 13864
rect 8300 13812 8352 13864
rect 11336 14016 11388 14068
rect 11980 14016 12032 14068
rect 12256 14016 12308 14068
rect 15660 14016 15712 14068
rect 20812 14016 20864 14068
rect 12992 13948 13044 14000
rect 11060 13812 11112 13864
rect 11980 13812 12032 13864
rect 12072 13855 12124 13864
rect 12072 13821 12081 13855
rect 12081 13821 12115 13855
rect 12115 13821 12124 13855
rect 12072 13812 12124 13821
rect 12440 13812 12492 13864
rect 3056 13787 3108 13796
rect 3056 13753 3065 13787
rect 3065 13753 3099 13787
rect 3099 13753 3108 13787
rect 3056 13744 3108 13753
rect 8576 13744 8628 13796
rect 12348 13744 12400 13796
rect 12808 13880 12860 13932
rect 14648 13855 14700 13864
rect 14648 13821 14657 13855
rect 14657 13821 14691 13855
rect 14691 13821 14700 13855
rect 14648 13812 14700 13821
rect 14832 13948 14884 14000
rect 14924 13923 14976 13932
rect 14924 13889 14933 13923
rect 14933 13889 14967 13923
rect 14967 13889 14976 13923
rect 14924 13880 14976 13889
rect 15016 13880 15068 13932
rect 15384 13812 15436 13864
rect 15936 13812 15988 13864
rect 18236 13880 18288 13932
rect 18328 13923 18380 13932
rect 18328 13889 18337 13923
rect 18337 13889 18371 13923
rect 18371 13889 18380 13923
rect 18328 13880 18380 13889
rect 18512 13880 18564 13932
rect 19616 13880 19668 13932
rect 15108 13787 15160 13796
rect 15108 13753 15117 13787
rect 15117 13753 15151 13787
rect 15151 13753 15160 13787
rect 15108 13744 15160 13753
rect 16120 13744 16172 13796
rect 18880 13744 18932 13796
rect 20904 13744 20956 13796
rect 21456 13744 21508 13796
rect 22376 14059 22428 14068
rect 22376 14025 22385 14059
rect 22385 14025 22419 14059
rect 22419 14025 22428 14059
rect 22376 14016 22428 14025
rect 23480 14016 23532 14068
rect 22100 13923 22152 13932
rect 22100 13889 22109 13923
rect 22109 13889 22143 13923
rect 22143 13889 22152 13923
rect 22100 13880 22152 13889
rect 22928 13923 22980 13932
rect 22928 13889 22937 13923
rect 22937 13889 22971 13923
rect 22971 13889 22980 13923
rect 22928 13880 22980 13889
rect 22008 13744 22060 13796
rect 22284 13812 22336 13864
rect 22560 13812 22612 13864
rect 23572 13948 23624 14000
rect 24768 14016 24820 14068
rect 25780 14016 25832 14068
rect 25136 13948 25188 14000
rect 23296 13923 23348 13932
rect 23296 13889 23305 13923
rect 23305 13889 23339 13923
rect 23339 13889 23348 13923
rect 23296 13880 23348 13889
rect 23388 13923 23440 13932
rect 23388 13889 23397 13923
rect 23397 13889 23431 13923
rect 23431 13889 23440 13923
rect 23388 13880 23440 13889
rect 24952 13880 25004 13932
rect 27528 13880 27580 13932
rect 23112 13812 23164 13864
rect 23572 13855 23624 13864
rect 23572 13821 23581 13855
rect 23581 13821 23615 13855
rect 23615 13821 23624 13855
rect 23572 13812 23624 13821
rect 24216 13812 24268 13864
rect 22376 13744 22428 13796
rect 23388 13744 23440 13796
rect 6828 13719 6880 13728
rect 6828 13685 6837 13719
rect 6837 13685 6871 13719
rect 6871 13685 6880 13719
rect 6828 13676 6880 13685
rect 8944 13719 8996 13728
rect 8944 13685 8953 13719
rect 8953 13685 8987 13719
rect 8987 13685 8996 13719
rect 8944 13676 8996 13685
rect 12164 13676 12216 13728
rect 13360 13676 13412 13728
rect 14372 13719 14424 13728
rect 14372 13685 14381 13719
rect 14381 13685 14415 13719
rect 14415 13685 14424 13719
rect 14372 13676 14424 13685
rect 15292 13676 15344 13728
rect 17776 13676 17828 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 2412 13515 2464 13524
rect 2412 13481 2421 13515
rect 2421 13481 2455 13515
rect 2455 13481 2464 13515
rect 2412 13472 2464 13481
rect 8576 13472 8628 13524
rect 8668 13515 8720 13524
rect 8668 13481 8677 13515
rect 8677 13481 8711 13515
rect 8711 13481 8720 13515
rect 8668 13472 8720 13481
rect 12072 13472 12124 13524
rect 12440 13515 12492 13524
rect 12440 13481 12449 13515
rect 12449 13481 12483 13515
rect 12483 13481 12492 13515
rect 12440 13472 12492 13481
rect 1952 13379 2004 13388
rect 1952 13345 1961 13379
rect 1961 13345 1995 13379
rect 1995 13345 2004 13379
rect 1952 13336 2004 13345
rect 2228 13379 2280 13388
rect 2228 13345 2237 13379
rect 2237 13345 2271 13379
rect 2271 13345 2280 13379
rect 2228 13336 2280 13345
rect 11888 13404 11940 13456
rect 22744 13472 22796 13524
rect 15936 13447 15988 13456
rect 15936 13413 15945 13447
rect 15945 13413 15979 13447
rect 15979 13413 15988 13447
rect 15936 13404 15988 13413
rect 17408 13447 17460 13456
rect 17408 13413 17417 13447
rect 17417 13413 17451 13447
rect 17451 13413 17460 13447
rect 17408 13404 17460 13413
rect 17868 13404 17920 13456
rect 1860 13311 1912 13320
rect 1860 13277 1869 13311
rect 1869 13277 1903 13311
rect 1903 13277 1912 13311
rect 1860 13268 1912 13277
rect 2964 13268 3016 13320
rect 6828 13311 6880 13320
rect 6828 13277 6837 13311
rect 6837 13277 6871 13311
rect 6871 13277 6880 13311
rect 6828 13268 6880 13277
rect 7104 13311 7156 13320
rect 7104 13277 7113 13311
rect 7113 13277 7147 13311
rect 7147 13277 7156 13311
rect 7104 13268 7156 13277
rect 7472 13311 7524 13320
rect 7472 13277 7481 13311
rect 7481 13277 7515 13311
rect 7515 13277 7524 13311
rect 7472 13268 7524 13277
rect 8116 13311 8168 13320
rect 8116 13277 8125 13311
rect 8125 13277 8159 13311
rect 8159 13277 8168 13311
rect 8116 13268 8168 13277
rect 8300 13336 8352 13388
rect 8300 13200 8352 13252
rect 8024 13132 8076 13184
rect 8944 13268 8996 13320
rect 9220 13311 9272 13320
rect 9220 13277 9229 13311
rect 9229 13277 9263 13311
rect 9263 13277 9272 13311
rect 9220 13268 9272 13277
rect 12256 13268 12308 13320
rect 12808 13336 12860 13388
rect 14004 13336 14056 13388
rect 16672 13336 16724 13388
rect 18052 13336 18104 13388
rect 19340 13336 19392 13388
rect 19984 13336 20036 13388
rect 13912 13268 13964 13320
rect 16212 13268 16264 13320
rect 12624 13243 12676 13252
rect 12624 13209 12633 13243
rect 12633 13209 12667 13243
rect 12667 13209 12676 13243
rect 12624 13200 12676 13209
rect 14372 13243 14424 13252
rect 14372 13209 14381 13243
rect 14381 13209 14415 13243
rect 14415 13209 14424 13243
rect 14372 13200 14424 13209
rect 14832 13200 14884 13252
rect 16948 13268 17000 13320
rect 17500 13311 17552 13320
rect 17500 13277 17509 13311
rect 17509 13277 17543 13311
rect 17543 13277 17552 13311
rect 17500 13268 17552 13277
rect 17040 13200 17092 13252
rect 17868 13311 17920 13320
rect 17868 13277 17877 13311
rect 17877 13277 17911 13311
rect 17911 13277 17920 13311
rect 17868 13268 17920 13277
rect 21272 13268 21324 13320
rect 19340 13200 19392 13252
rect 12716 13132 12768 13184
rect 12808 13175 12860 13184
rect 12808 13141 12817 13175
rect 12817 13141 12851 13175
rect 12851 13141 12860 13175
rect 12808 13132 12860 13141
rect 14556 13132 14608 13184
rect 15752 13132 15804 13184
rect 16120 13132 16172 13184
rect 16304 13175 16356 13184
rect 16304 13141 16313 13175
rect 16313 13141 16347 13175
rect 16347 13141 16356 13175
rect 16304 13132 16356 13141
rect 20076 13175 20128 13184
rect 20076 13141 20085 13175
rect 20085 13141 20119 13175
rect 20119 13141 20128 13175
rect 20076 13132 20128 13141
rect 20260 13132 20312 13184
rect 22008 13404 22060 13456
rect 21456 13336 21508 13388
rect 21548 13268 21600 13320
rect 22100 13311 22152 13320
rect 22100 13277 22109 13311
rect 22109 13277 22143 13311
rect 22143 13277 22152 13311
rect 22100 13268 22152 13277
rect 22284 13268 22336 13320
rect 22836 13311 22888 13320
rect 22836 13277 22845 13311
rect 22845 13277 22879 13311
rect 22879 13277 22888 13311
rect 22836 13268 22888 13277
rect 22928 13311 22980 13320
rect 22928 13277 22937 13311
rect 22937 13277 22971 13311
rect 22971 13277 22980 13311
rect 22928 13268 22980 13277
rect 23480 13379 23532 13388
rect 23480 13345 23489 13379
rect 23489 13345 23523 13379
rect 23523 13345 23532 13379
rect 23480 13336 23532 13345
rect 23940 13404 23992 13456
rect 24032 13336 24084 13388
rect 24768 13311 24820 13320
rect 24768 13277 24777 13311
rect 24777 13277 24811 13311
rect 24811 13277 24820 13311
rect 24768 13268 24820 13277
rect 22284 13175 22336 13184
rect 22284 13141 22293 13175
rect 22293 13141 22327 13175
rect 22327 13141 22336 13175
rect 22284 13132 22336 13141
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 7104 12928 7156 12980
rect 8300 12928 8352 12980
rect 9220 12928 9272 12980
rect 12256 12971 12308 12980
rect 12256 12937 12265 12971
rect 12265 12937 12299 12971
rect 12299 12937 12308 12971
rect 12256 12928 12308 12937
rect 12624 12928 12676 12980
rect 14648 12928 14700 12980
rect 2964 12792 3016 12844
rect 5540 12792 5592 12844
rect 6184 12835 6236 12844
rect 6184 12801 6193 12835
rect 6193 12801 6227 12835
rect 6227 12801 6236 12835
rect 6184 12792 6236 12801
rect 6644 12835 6696 12844
rect 6644 12801 6653 12835
rect 6653 12801 6687 12835
rect 6687 12801 6696 12835
rect 6644 12792 6696 12801
rect 8024 12835 8076 12844
rect 8024 12801 8033 12835
rect 8033 12801 8067 12835
rect 8067 12801 8076 12835
rect 8024 12792 8076 12801
rect 8208 12792 8260 12844
rect 11428 12792 11480 12844
rect 12072 12903 12124 12912
rect 12072 12869 12097 12903
rect 12097 12869 12124 12903
rect 12072 12860 12124 12869
rect 12716 12860 12768 12912
rect 12348 12835 12400 12844
rect 12348 12801 12357 12835
rect 12357 12801 12391 12835
rect 12391 12801 12400 12835
rect 12348 12792 12400 12801
rect 12624 12792 12676 12844
rect 14556 12792 14608 12844
rect 16304 12860 16356 12912
rect 15292 12835 15344 12844
rect 15292 12801 15301 12835
rect 15301 12801 15335 12835
rect 15335 12801 15344 12835
rect 15292 12792 15344 12801
rect 15476 12835 15528 12844
rect 15476 12801 15485 12835
rect 15485 12801 15519 12835
rect 15519 12801 15528 12835
rect 15476 12792 15528 12801
rect 15568 12792 15620 12844
rect 15752 12835 15804 12844
rect 15752 12801 15761 12835
rect 15761 12801 15795 12835
rect 15795 12801 15804 12835
rect 15752 12792 15804 12801
rect 18052 12835 18104 12844
rect 18052 12801 18061 12835
rect 18061 12801 18095 12835
rect 18095 12801 18104 12835
rect 18052 12792 18104 12801
rect 20628 12928 20680 12980
rect 18236 12860 18288 12912
rect 18420 12835 18472 12844
rect 18420 12801 18429 12835
rect 18429 12801 18463 12835
rect 18463 12801 18472 12835
rect 18420 12792 18472 12801
rect 18512 12792 18564 12844
rect 20076 12860 20128 12912
rect 21272 12971 21324 12980
rect 21272 12937 21281 12971
rect 21281 12937 21315 12971
rect 21315 12937 21324 12971
rect 21272 12928 21324 12937
rect 22744 12928 22796 12980
rect 23296 12928 23348 12980
rect 22376 12860 22428 12912
rect 20904 12792 20956 12844
rect 21824 12835 21876 12844
rect 21824 12801 21833 12835
rect 21833 12801 21867 12835
rect 21867 12801 21876 12835
rect 21824 12792 21876 12801
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 22008 12792 22060 12801
rect 2228 12724 2280 12776
rect 5356 12767 5408 12776
rect 5356 12733 5365 12767
rect 5365 12733 5399 12767
rect 5399 12733 5408 12767
rect 5356 12724 5408 12733
rect 9772 12724 9824 12776
rect 15200 12724 15252 12776
rect 17868 12724 17920 12776
rect 19156 12724 19208 12776
rect 19524 12767 19576 12776
rect 19524 12733 19533 12767
rect 19533 12733 19567 12767
rect 19567 12733 19576 12767
rect 19524 12724 19576 12733
rect 19800 12767 19852 12776
rect 19800 12733 19809 12767
rect 19809 12733 19843 12767
rect 19843 12733 19852 12767
rect 19800 12724 19852 12733
rect 20812 12724 20864 12776
rect 25780 12792 25832 12844
rect 11796 12656 11848 12708
rect 2228 12631 2280 12640
rect 2228 12597 2237 12631
rect 2237 12597 2271 12631
rect 2271 12597 2280 12631
rect 2228 12588 2280 12597
rect 12072 12631 12124 12640
rect 12072 12597 12081 12631
rect 12081 12597 12115 12631
rect 12115 12597 12124 12631
rect 12072 12588 12124 12597
rect 17040 12656 17092 12708
rect 18880 12699 18932 12708
rect 18880 12665 18889 12699
rect 18889 12665 18923 12699
rect 18923 12665 18932 12699
rect 18880 12656 18932 12665
rect 16856 12588 16908 12640
rect 19340 12656 19392 12708
rect 22284 12656 22336 12708
rect 23480 12656 23532 12708
rect 19156 12588 19208 12640
rect 22100 12588 22152 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 16212 12384 16264 12436
rect 3240 12316 3292 12368
rect 3056 12248 3108 12300
rect 3240 12223 3292 12232
rect 3240 12189 3249 12223
rect 3249 12189 3283 12223
rect 3283 12189 3292 12223
rect 3240 12180 3292 12189
rect 7380 12316 7432 12368
rect 5356 12248 5408 12300
rect 4712 12223 4764 12232
rect 4712 12189 4721 12223
rect 4721 12189 4755 12223
rect 4755 12189 4764 12223
rect 4712 12180 4764 12189
rect 4804 12180 4856 12232
rect 8300 12291 8352 12300
rect 8300 12257 8309 12291
rect 8309 12257 8343 12291
rect 8343 12257 8352 12291
rect 8300 12248 8352 12257
rect 5540 12180 5592 12232
rect 6184 12223 6236 12232
rect 6184 12189 6193 12223
rect 6193 12189 6227 12223
rect 6227 12189 6236 12223
rect 6184 12180 6236 12189
rect 6644 12180 6696 12232
rect 7104 12180 7156 12232
rect 11336 12223 11388 12232
rect 11336 12189 11345 12223
rect 11345 12189 11379 12223
rect 11379 12189 11388 12223
rect 11336 12180 11388 12189
rect 15568 12316 15620 12368
rect 16488 12316 16540 12368
rect 16580 12359 16632 12368
rect 16580 12325 16589 12359
rect 16589 12325 16623 12359
rect 16623 12325 16632 12359
rect 16580 12316 16632 12325
rect 12256 12291 12308 12300
rect 12256 12257 12265 12291
rect 12265 12257 12299 12291
rect 12299 12257 12308 12291
rect 12256 12248 12308 12257
rect 12440 12291 12492 12300
rect 12440 12257 12449 12291
rect 12449 12257 12483 12291
rect 12483 12257 12492 12291
rect 12440 12248 12492 12257
rect 12532 12248 12584 12300
rect 12808 12248 12860 12300
rect 16856 12248 16908 12300
rect 18788 12384 18840 12436
rect 18052 12316 18104 12368
rect 19156 12316 19208 12368
rect 19340 12384 19392 12436
rect 7748 12112 7800 12164
rect 4528 12044 4580 12096
rect 11152 12087 11204 12096
rect 11152 12053 11161 12087
rect 11161 12053 11195 12087
rect 11195 12053 11204 12087
rect 11152 12044 11204 12053
rect 11520 12087 11572 12096
rect 11520 12053 11529 12087
rect 11529 12053 11563 12087
rect 11563 12053 11572 12087
rect 11520 12044 11572 12053
rect 16028 12180 16080 12232
rect 16304 12223 16356 12232
rect 16304 12189 16313 12223
rect 16313 12189 16347 12223
rect 16347 12189 16356 12223
rect 16304 12180 16356 12189
rect 18512 12248 18564 12300
rect 19340 12248 19392 12300
rect 12808 12112 12860 12164
rect 13268 12112 13320 12164
rect 17132 12180 17184 12232
rect 17224 12223 17276 12232
rect 17224 12189 17233 12223
rect 17233 12189 17267 12223
rect 17267 12189 17276 12223
rect 17224 12180 17276 12189
rect 18052 12180 18104 12232
rect 18420 12180 18472 12232
rect 18788 12223 18840 12232
rect 18788 12189 18797 12223
rect 18797 12189 18831 12223
rect 18831 12189 18840 12223
rect 18788 12180 18840 12189
rect 19156 12180 19208 12232
rect 19892 12384 19944 12436
rect 21088 12384 21140 12436
rect 22008 12384 22060 12436
rect 19892 12248 19944 12300
rect 21824 12316 21876 12368
rect 20536 12291 20588 12300
rect 20536 12257 20545 12291
rect 20545 12257 20579 12291
rect 20579 12257 20588 12291
rect 20536 12248 20588 12257
rect 20720 12248 20772 12300
rect 21272 12291 21324 12300
rect 12624 12044 12676 12096
rect 12900 12044 12952 12096
rect 13176 12044 13228 12096
rect 16580 12044 16632 12096
rect 17040 12044 17092 12096
rect 18236 12087 18288 12096
rect 18236 12053 18245 12087
rect 18245 12053 18279 12087
rect 18279 12053 18288 12087
rect 18236 12044 18288 12053
rect 18696 12087 18748 12096
rect 18696 12053 18705 12087
rect 18705 12053 18739 12087
rect 18739 12053 18748 12087
rect 18696 12044 18748 12053
rect 19064 12044 19116 12096
rect 20260 12223 20312 12232
rect 20260 12189 20269 12223
rect 20269 12189 20303 12223
rect 20303 12189 20312 12223
rect 20260 12180 20312 12189
rect 19800 12112 19852 12164
rect 20628 12223 20680 12232
rect 20628 12189 20637 12223
rect 20637 12189 20671 12223
rect 20671 12189 20680 12223
rect 20628 12180 20680 12189
rect 20812 12223 20864 12232
rect 20812 12189 20821 12223
rect 20821 12189 20855 12223
rect 20855 12189 20864 12223
rect 20812 12180 20864 12189
rect 21272 12257 21281 12291
rect 21281 12257 21315 12291
rect 21315 12257 21324 12291
rect 21272 12248 21324 12257
rect 21088 12180 21140 12232
rect 21548 12112 21600 12164
rect 23204 12112 23256 12164
rect 22468 12044 22520 12096
rect 23112 12044 23164 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 3240 11840 3292 11892
rect 8208 11840 8260 11892
rect 11336 11883 11388 11892
rect 11336 11849 11345 11883
rect 11345 11849 11379 11883
rect 11379 11849 11388 11883
rect 11336 11840 11388 11849
rect 11520 11883 11572 11892
rect 11520 11849 11529 11883
rect 11529 11849 11563 11883
rect 11563 11849 11572 11883
rect 11520 11840 11572 11849
rect 2228 11772 2280 11824
rect 848 11704 900 11756
rect 2320 11704 2372 11756
rect 4804 11772 4856 11824
rect 4068 11704 4120 11756
rect 3332 11679 3384 11688
rect 3332 11645 3341 11679
rect 3341 11645 3375 11679
rect 3375 11645 3384 11679
rect 3332 11636 3384 11645
rect 2780 11568 2832 11620
rect 3516 11679 3568 11688
rect 3516 11645 3525 11679
rect 3525 11645 3559 11679
rect 3559 11645 3568 11679
rect 3516 11636 3568 11645
rect 4528 11679 4580 11688
rect 4528 11645 4537 11679
rect 4537 11645 4571 11679
rect 4571 11645 4580 11679
rect 4528 11636 4580 11645
rect 4712 11704 4764 11756
rect 5080 11747 5132 11756
rect 5080 11713 5089 11747
rect 5089 11713 5123 11747
rect 5123 11713 5132 11747
rect 5080 11704 5132 11713
rect 10508 11772 10560 11824
rect 7104 11704 7156 11756
rect 7748 11747 7800 11756
rect 7748 11713 7757 11747
rect 7757 11713 7791 11747
rect 7791 11713 7800 11747
rect 7748 11704 7800 11713
rect 10876 11747 10928 11756
rect 10876 11713 10885 11747
rect 10885 11713 10919 11747
rect 10919 11713 10928 11747
rect 10876 11704 10928 11713
rect 5540 11568 5592 11620
rect 6736 11500 6788 11552
rect 11704 11747 11756 11756
rect 11704 11713 11713 11747
rect 11713 11713 11747 11747
rect 11747 11713 11756 11747
rect 11704 11704 11756 11713
rect 12532 11815 12584 11824
rect 11980 11747 12032 11756
rect 11980 11713 11989 11747
rect 11989 11713 12023 11747
rect 12023 11713 12032 11747
rect 11980 11704 12032 11713
rect 12532 11781 12541 11815
rect 12541 11781 12575 11815
rect 12575 11781 12584 11815
rect 12532 11772 12584 11781
rect 12164 11747 12216 11756
rect 12164 11713 12173 11747
rect 12173 11713 12207 11747
rect 12207 11713 12216 11747
rect 12164 11704 12216 11713
rect 12256 11747 12308 11756
rect 12256 11713 12265 11747
rect 12265 11713 12299 11747
rect 12299 11713 12308 11747
rect 12256 11704 12308 11713
rect 12440 11704 12492 11756
rect 13820 11840 13872 11892
rect 16212 11840 16264 11892
rect 16304 11840 16356 11892
rect 19432 11840 19484 11892
rect 19524 11840 19576 11892
rect 20168 11840 20220 11892
rect 22836 11840 22888 11892
rect 23296 11840 23348 11892
rect 23480 11840 23532 11892
rect 14740 11704 14792 11756
rect 17040 11772 17092 11824
rect 17776 11772 17828 11824
rect 15568 11747 15620 11756
rect 15568 11713 15577 11747
rect 15577 11713 15611 11747
rect 15611 11713 15620 11747
rect 15568 11704 15620 11713
rect 15844 11747 15896 11756
rect 15844 11713 15853 11747
rect 15853 11713 15887 11747
rect 15887 11713 15896 11747
rect 15844 11704 15896 11713
rect 15936 11704 15988 11756
rect 12164 11568 12216 11620
rect 12716 11568 12768 11620
rect 13820 11500 13872 11552
rect 16120 11568 16172 11620
rect 16580 11704 16632 11756
rect 16672 11747 16724 11756
rect 16672 11713 16681 11747
rect 16681 11713 16715 11747
rect 16715 11713 16724 11747
rect 16672 11704 16724 11713
rect 18696 11747 18748 11756
rect 18696 11713 18705 11747
rect 18705 11713 18739 11747
rect 18739 11713 18748 11747
rect 18696 11704 18748 11713
rect 18880 11747 18932 11756
rect 18880 11713 18889 11747
rect 18889 11713 18923 11747
rect 18923 11713 18932 11747
rect 18880 11704 18932 11713
rect 19064 11747 19116 11756
rect 19064 11713 19073 11747
rect 19073 11713 19107 11747
rect 19107 11713 19116 11747
rect 19064 11704 19116 11713
rect 18236 11636 18288 11688
rect 19524 11747 19576 11756
rect 19524 11713 19533 11747
rect 19533 11713 19567 11747
rect 19567 11713 19576 11747
rect 19524 11704 19576 11713
rect 19708 11704 19760 11756
rect 20996 11636 21048 11688
rect 22836 11704 22888 11756
rect 23204 11747 23256 11756
rect 23204 11713 23213 11747
rect 23213 11713 23247 11747
rect 23247 11713 23256 11747
rect 23204 11704 23256 11713
rect 23296 11747 23348 11756
rect 23296 11713 23305 11747
rect 23305 11713 23339 11747
rect 23339 11713 23348 11747
rect 23296 11704 23348 11713
rect 23480 11704 23532 11756
rect 24032 11636 24084 11688
rect 16488 11568 16540 11620
rect 18328 11568 18380 11620
rect 22744 11568 22796 11620
rect 23664 11568 23716 11620
rect 17316 11500 17368 11552
rect 18788 11500 18840 11552
rect 20720 11500 20772 11552
rect 21272 11500 21324 11552
rect 23020 11500 23072 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 2964 11296 3016 11348
rect 3516 11296 3568 11348
rect 10048 11339 10100 11348
rect 10048 11305 10057 11339
rect 10057 11305 10091 11339
rect 10091 11305 10100 11339
rect 10048 11296 10100 11305
rect 10232 11339 10284 11348
rect 10232 11305 10241 11339
rect 10241 11305 10275 11339
rect 10275 11305 10284 11339
rect 10232 11296 10284 11305
rect 10784 11296 10836 11348
rect 12072 11296 12124 11348
rect 12440 11296 12492 11348
rect 12532 11339 12584 11348
rect 12532 11305 12541 11339
rect 12541 11305 12575 11339
rect 12575 11305 12584 11339
rect 12532 11296 12584 11305
rect 13176 11296 13228 11348
rect 14464 11296 14516 11348
rect 6736 11228 6788 11280
rect 2228 11203 2280 11212
rect 2228 11169 2237 11203
rect 2237 11169 2271 11203
rect 2271 11169 2280 11203
rect 2228 11160 2280 11169
rect 7196 11203 7248 11212
rect 7196 11169 7205 11203
rect 7205 11169 7239 11203
rect 7239 11169 7248 11203
rect 7196 11160 7248 11169
rect 10140 11160 10192 11212
rect 11520 11228 11572 11280
rect 11612 11271 11664 11280
rect 11612 11237 11621 11271
rect 11621 11237 11655 11271
rect 11655 11237 11664 11271
rect 11612 11228 11664 11237
rect 2320 11135 2372 11144
rect 2320 11101 2329 11135
rect 2329 11101 2363 11135
rect 2363 11101 2372 11135
rect 2320 11092 2372 11101
rect 7380 11092 7432 11144
rect 10508 11135 10560 11144
rect 10508 11101 10517 11135
rect 10517 11101 10551 11135
rect 10551 11101 10560 11135
rect 10508 11092 10560 11101
rect 11152 11160 11204 11212
rect 11980 11160 12032 11212
rect 10784 11135 10836 11144
rect 10784 11101 10793 11135
rect 10793 11101 10827 11135
rect 10827 11101 10836 11135
rect 10784 11092 10836 11101
rect 10876 11135 10928 11144
rect 10876 11101 10885 11135
rect 10885 11101 10919 11135
rect 10919 11101 10928 11135
rect 10876 11092 10928 11101
rect 11336 11135 11388 11144
rect 11336 11101 11345 11135
rect 11345 11101 11379 11135
rect 11379 11101 11388 11135
rect 11336 11092 11388 11101
rect 12256 11135 12308 11144
rect 12256 11101 12265 11135
rect 12265 11101 12299 11135
rect 12299 11101 12308 11135
rect 12256 11092 12308 11101
rect 6552 11067 6604 11076
rect 6552 11033 6561 11067
rect 6561 11033 6595 11067
rect 6595 11033 6604 11067
rect 6552 11024 6604 11033
rect 9772 11024 9824 11076
rect 7104 10999 7156 11008
rect 7104 10965 7113 10999
rect 7113 10965 7147 10999
rect 7147 10965 7156 10999
rect 7104 10956 7156 10965
rect 9956 10956 10008 11008
rect 11060 11024 11112 11076
rect 12072 11067 12124 11076
rect 12072 11033 12081 11067
rect 12081 11033 12115 11067
rect 12115 11033 12124 11067
rect 12072 11024 12124 11033
rect 12164 11024 12216 11076
rect 11796 10956 11848 11008
rect 11888 10956 11940 11008
rect 13084 11135 13136 11144
rect 13084 11101 13093 11135
rect 13093 11101 13127 11135
rect 13127 11101 13136 11135
rect 13084 11092 13136 11101
rect 14556 11092 14608 11144
rect 14924 11160 14976 11212
rect 15384 11160 15436 11212
rect 16580 11296 16632 11348
rect 16764 11296 16816 11348
rect 18328 11296 18380 11348
rect 19248 11296 19300 11348
rect 20260 11296 20312 11348
rect 18052 11228 18104 11280
rect 14740 11135 14792 11144
rect 14740 11101 14749 11135
rect 14749 11101 14783 11135
rect 14783 11101 14792 11135
rect 14740 11092 14792 11101
rect 13176 11024 13228 11076
rect 15292 11135 15344 11144
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 15568 11092 15620 11144
rect 16856 11160 16908 11212
rect 19064 11160 19116 11212
rect 12532 10956 12584 11008
rect 13268 10956 13320 11008
rect 15016 10956 15068 11008
rect 15476 11067 15528 11076
rect 15476 11033 15485 11067
rect 15485 11033 15519 11067
rect 15519 11033 15528 11067
rect 15476 11024 15528 11033
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16028 11092 16080 11101
rect 18052 11135 18104 11144
rect 18052 11101 18061 11135
rect 18061 11101 18095 11135
rect 18095 11101 18104 11135
rect 18052 11092 18104 11101
rect 18696 11092 18748 11144
rect 22008 11160 22060 11212
rect 16304 11024 16356 11076
rect 16856 11024 16908 11076
rect 20996 11092 21048 11144
rect 21180 11135 21232 11144
rect 21180 11101 21189 11135
rect 21189 11101 21223 11135
rect 21223 11101 21232 11135
rect 21180 11092 21232 11101
rect 21732 11092 21784 11144
rect 23020 11228 23072 11280
rect 23112 11228 23164 11280
rect 23480 11296 23532 11348
rect 23664 11296 23716 11348
rect 24492 11228 24544 11280
rect 21456 11024 21508 11076
rect 22192 11024 22244 11076
rect 23020 11092 23072 11144
rect 23940 11160 23992 11212
rect 24032 11160 24084 11212
rect 23756 11024 23808 11076
rect 23848 11067 23900 11076
rect 23848 11033 23857 11067
rect 23857 11033 23891 11067
rect 23891 11033 23900 11067
rect 23848 11024 23900 11033
rect 23940 11024 23992 11076
rect 16120 10956 16172 11008
rect 18420 10956 18472 11008
rect 20720 10999 20772 11008
rect 20720 10965 20729 10999
rect 20729 10965 20763 10999
rect 20763 10965 20772 10999
rect 20720 10956 20772 10965
rect 22468 10956 22520 11008
rect 23020 10956 23072 11008
rect 23296 10956 23348 11008
rect 25228 11024 25280 11076
rect 25320 10956 25372 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 2320 10752 2372 10804
rect 1952 10684 2004 10736
rect 2688 10752 2740 10804
rect 2780 10752 2832 10804
rect 6552 10752 6604 10804
rect 8116 10795 8168 10804
rect 8116 10761 8125 10795
rect 8125 10761 8159 10795
rect 8159 10761 8168 10795
rect 8116 10752 8168 10761
rect 2136 10412 2188 10464
rect 2596 10616 2648 10668
rect 2964 10591 3016 10600
rect 2964 10557 2973 10591
rect 2973 10557 3007 10591
rect 3007 10557 3016 10591
rect 2964 10548 3016 10557
rect 3332 10616 3384 10668
rect 7656 10684 7708 10736
rect 10876 10752 10928 10804
rect 12164 10752 12216 10804
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 5540 10591 5592 10600
rect 5540 10557 5549 10591
rect 5549 10557 5583 10591
rect 5583 10557 5592 10591
rect 7380 10616 7432 10668
rect 8392 10659 8444 10668
rect 8392 10625 8401 10659
rect 8401 10625 8435 10659
rect 8435 10625 8444 10659
rect 8392 10616 8444 10625
rect 12348 10752 12400 10804
rect 12440 10752 12492 10804
rect 12900 10795 12952 10804
rect 12900 10761 12930 10795
rect 12930 10761 12952 10795
rect 12900 10752 12952 10761
rect 14004 10752 14056 10804
rect 8852 10659 8904 10668
rect 8852 10625 8861 10659
rect 8861 10625 8895 10659
rect 8895 10625 8904 10659
rect 8852 10616 8904 10625
rect 5540 10548 5592 10557
rect 3976 10480 4028 10532
rect 7196 10548 7248 10600
rect 8300 10548 8352 10600
rect 9128 10548 9180 10600
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 11060 10616 11112 10668
rect 11428 10616 11480 10668
rect 10048 10548 10100 10600
rect 11612 10548 11664 10600
rect 11336 10480 11388 10532
rect 11888 10659 11940 10668
rect 11888 10625 11897 10659
rect 11897 10625 11931 10659
rect 11931 10625 11940 10659
rect 11888 10616 11940 10625
rect 12532 10684 12584 10736
rect 12624 10684 12676 10736
rect 14096 10684 14148 10736
rect 14924 10752 14976 10804
rect 15108 10795 15160 10804
rect 15108 10761 15117 10795
rect 15117 10761 15151 10795
rect 15151 10761 15160 10795
rect 15108 10752 15160 10761
rect 15292 10752 15344 10804
rect 15936 10752 15988 10804
rect 18880 10752 18932 10804
rect 12256 10659 12308 10668
rect 12256 10625 12265 10659
rect 12265 10625 12299 10659
rect 12299 10625 12308 10659
rect 12256 10616 12308 10625
rect 11796 10548 11848 10600
rect 14372 10616 14424 10668
rect 14832 10684 14884 10736
rect 15384 10684 15436 10736
rect 15568 10684 15620 10736
rect 12532 10548 12584 10600
rect 12716 10548 12768 10600
rect 14924 10659 14976 10668
rect 14924 10625 14933 10659
rect 14933 10625 14967 10659
rect 14967 10625 14976 10659
rect 14924 10616 14976 10625
rect 15016 10616 15068 10668
rect 15844 10616 15896 10668
rect 16764 10727 16816 10736
rect 16764 10693 16773 10727
rect 16773 10693 16807 10727
rect 16807 10693 16816 10727
rect 16764 10684 16816 10693
rect 17224 10684 17276 10736
rect 19708 10684 19760 10736
rect 16120 10659 16172 10668
rect 16120 10625 16129 10659
rect 16129 10625 16163 10659
rect 16163 10625 16172 10659
rect 16120 10616 16172 10625
rect 17040 10616 17092 10668
rect 18512 10616 18564 10668
rect 19248 10616 19300 10668
rect 19616 10616 19668 10668
rect 20720 10752 20772 10804
rect 20536 10659 20588 10668
rect 20536 10625 20545 10659
rect 20545 10625 20579 10659
rect 20579 10625 20588 10659
rect 20536 10616 20588 10625
rect 12348 10480 12400 10532
rect 8208 10412 8260 10464
rect 10600 10412 10652 10464
rect 12808 10412 12860 10464
rect 12992 10480 13044 10532
rect 15384 10591 15436 10600
rect 15384 10557 15393 10591
rect 15393 10557 15427 10591
rect 15427 10557 15436 10591
rect 15384 10548 15436 10557
rect 13912 10480 13964 10532
rect 18696 10591 18748 10600
rect 18696 10557 18705 10591
rect 18705 10557 18739 10591
rect 18739 10557 18748 10591
rect 18696 10548 18748 10557
rect 18788 10591 18840 10600
rect 18788 10557 18797 10591
rect 18797 10557 18831 10591
rect 18831 10557 18840 10591
rect 18788 10548 18840 10557
rect 18880 10591 18932 10600
rect 18880 10557 18889 10591
rect 18889 10557 18923 10591
rect 18923 10557 18932 10591
rect 18880 10548 18932 10557
rect 16672 10480 16724 10532
rect 17316 10480 17368 10532
rect 19984 10548 20036 10600
rect 20168 10548 20220 10600
rect 20996 10684 21048 10736
rect 22836 10727 22888 10736
rect 22836 10693 22845 10727
rect 22845 10693 22879 10727
rect 22879 10693 22888 10727
rect 22836 10684 22888 10693
rect 23112 10684 23164 10736
rect 19248 10480 19300 10532
rect 16856 10412 16908 10464
rect 18052 10412 18104 10464
rect 18972 10412 19024 10464
rect 19892 10455 19944 10464
rect 19892 10421 19901 10455
rect 19901 10421 19935 10455
rect 19935 10421 19944 10455
rect 19892 10412 19944 10421
rect 19984 10412 20036 10464
rect 21456 10659 21508 10668
rect 21456 10625 21465 10659
rect 21465 10625 21499 10659
rect 21499 10625 21508 10659
rect 21456 10616 21508 10625
rect 21272 10548 21324 10600
rect 23480 10684 23532 10736
rect 23664 10752 23716 10804
rect 23848 10752 23900 10804
rect 24032 10684 24084 10736
rect 25320 10659 25372 10668
rect 25320 10625 25329 10659
rect 25329 10625 25363 10659
rect 25363 10625 25372 10659
rect 25320 10616 25372 10625
rect 24584 10480 24636 10532
rect 24768 10480 24820 10532
rect 23020 10455 23072 10464
rect 23020 10421 23029 10455
rect 23029 10421 23063 10455
rect 23063 10421 23072 10455
rect 23020 10412 23072 10421
rect 24676 10412 24728 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 8116 10208 8168 10260
rect 8852 10208 8904 10260
rect 8208 10183 8260 10192
rect 8208 10149 8217 10183
rect 8217 10149 8251 10183
rect 8251 10149 8260 10183
rect 8208 10140 8260 10149
rect 8392 10140 8444 10192
rect 9312 10251 9364 10260
rect 9312 10217 9321 10251
rect 9321 10217 9355 10251
rect 9355 10217 9364 10251
rect 9312 10208 9364 10217
rect 9956 10251 10008 10260
rect 9956 10217 9965 10251
rect 9965 10217 9999 10251
rect 9999 10217 10008 10251
rect 9956 10208 10008 10217
rect 10600 10208 10652 10260
rect 13912 10251 13964 10260
rect 13912 10217 13921 10251
rect 13921 10217 13955 10251
rect 13955 10217 13964 10251
rect 13912 10208 13964 10217
rect 14004 10208 14056 10260
rect 12900 10140 12952 10192
rect 13084 10140 13136 10192
rect 2136 10115 2188 10124
rect 2136 10081 2145 10115
rect 2145 10081 2179 10115
rect 2179 10081 2188 10115
rect 2136 10072 2188 10081
rect 7932 10072 7984 10124
rect 2596 10004 2648 10056
rect 7380 10004 7432 10056
rect 7656 10004 7708 10056
rect 12256 10072 12308 10124
rect 12808 10072 12860 10124
rect 7472 9936 7524 9988
rect 10140 10004 10192 10056
rect 11152 10047 11204 10056
rect 11152 10013 11161 10047
rect 11161 10013 11195 10047
rect 11195 10013 11204 10047
rect 11152 10004 11204 10013
rect 12440 10047 12492 10056
rect 12440 10013 12449 10047
rect 12449 10013 12483 10047
rect 12483 10013 12492 10047
rect 12440 10004 12492 10013
rect 8300 9936 8352 9988
rect 9128 9979 9180 9988
rect 9128 9945 9153 9979
rect 9153 9945 9180 9979
rect 9128 9936 9180 9945
rect 11428 9936 11480 9988
rect 11980 9936 12032 9988
rect 12348 9936 12400 9988
rect 12624 9936 12676 9988
rect 13084 10047 13136 10056
rect 13084 10013 13093 10047
rect 13093 10013 13127 10047
rect 13127 10013 13136 10047
rect 13084 10004 13136 10013
rect 2964 9868 3016 9920
rect 8760 9868 8812 9920
rect 9588 9911 9640 9920
rect 9588 9877 9597 9911
rect 9597 9877 9631 9911
rect 9631 9877 9640 9911
rect 9588 9868 9640 9877
rect 9680 9911 9732 9920
rect 9680 9877 9689 9911
rect 9689 9877 9723 9911
rect 9723 9877 9732 9911
rect 9680 9868 9732 9877
rect 9772 9868 9824 9920
rect 11060 9911 11112 9920
rect 11060 9877 11069 9911
rect 11069 9877 11103 9911
rect 11103 9877 11112 9911
rect 11060 9868 11112 9877
rect 12808 9868 12860 9920
rect 14096 10047 14148 10056
rect 14096 10013 14105 10047
rect 14105 10013 14139 10047
rect 14139 10013 14148 10047
rect 14096 10004 14148 10013
rect 14832 10251 14884 10260
rect 14832 10217 14841 10251
rect 14841 10217 14875 10251
rect 14875 10217 14884 10251
rect 14832 10208 14884 10217
rect 15292 10251 15344 10260
rect 15292 10217 15326 10251
rect 15326 10217 15344 10251
rect 15292 10208 15344 10217
rect 15752 10208 15804 10260
rect 16212 10208 16264 10260
rect 18144 10208 18196 10260
rect 18788 10208 18840 10260
rect 20996 10208 21048 10260
rect 21456 10208 21508 10260
rect 22560 10208 22612 10260
rect 23664 10208 23716 10260
rect 23940 10208 23992 10260
rect 15292 10072 15344 10124
rect 14464 10047 14516 10056
rect 14464 10013 14473 10047
rect 14473 10013 14507 10047
rect 14507 10013 14516 10047
rect 14464 10004 14516 10013
rect 14924 10004 14976 10056
rect 15384 10004 15436 10056
rect 18604 10140 18656 10192
rect 19892 10140 19944 10192
rect 16856 10072 16908 10124
rect 16488 10047 16540 10056
rect 16488 10013 16497 10047
rect 16497 10013 16531 10047
rect 16531 10013 16540 10047
rect 16488 10004 16540 10013
rect 16948 10047 17000 10056
rect 16948 10013 16962 10047
rect 16962 10013 16996 10047
rect 16996 10013 17000 10047
rect 16948 10004 17000 10013
rect 17316 10004 17368 10056
rect 17684 10004 17736 10056
rect 17960 10047 18012 10056
rect 17960 10013 17969 10047
rect 17969 10013 18003 10047
rect 18003 10013 18012 10047
rect 17960 10004 18012 10013
rect 18512 10115 18564 10124
rect 18512 10081 18521 10115
rect 18521 10081 18555 10115
rect 18555 10081 18564 10115
rect 18512 10072 18564 10081
rect 20168 10115 20220 10124
rect 20168 10081 20177 10115
rect 20177 10081 20211 10115
rect 20211 10081 20220 10115
rect 20168 10072 20220 10081
rect 22468 10140 22520 10192
rect 21640 10072 21692 10124
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 22744 10004 22796 10056
rect 23572 10140 23624 10192
rect 23756 10072 23808 10124
rect 24308 10072 24360 10124
rect 24400 10115 24452 10124
rect 24400 10081 24409 10115
rect 24409 10081 24443 10115
rect 24443 10081 24452 10115
rect 24400 10072 24452 10081
rect 24676 10115 24728 10124
rect 24676 10081 24685 10115
rect 24685 10081 24719 10115
rect 24719 10081 24728 10115
rect 24676 10072 24728 10081
rect 15016 9868 15068 9920
rect 15200 9868 15252 9920
rect 16764 9979 16816 9988
rect 16764 9945 16773 9979
rect 16773 9945 16807 9979
rect 16807 9945 16816 9979
rect 16764 9936 16816 9945
rect 16856 9979 16908 9988
rect 16856 9945 16865 9979
rect 16865 9945 16899 9979
rect 16899 9945 16908 9979
rect 16856 9936 16908 9945
rect 18052 9936 18104 9988
rect 17132 9868 17184 9920
rect 20904 9936 20956 9988
rect 24952 9936 25004 9988
rect 25136 9936 25188 9988
rect 22836 9868 22888 9920
rect 23572 9868 23624 9920
rect 24216 9868 24268 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 5632 9664 5684 9716
rect 8300 9664 8352 9716
rect 8760 9707 8812 9716
rect 8760 9673 8769 9707
rect 8769 9673 8803 9707
rect 8803 9673 8812 9707
rect 8760 9664 8812 9673
rect 14464 9664 14516 9716
rect 14740 9664 14792 9716
rect 15476 9664 15528 9716
rect 16488 9664 16540 9716
rect 17960 9664 18012 9716
rect 18880 9664 18932 9716
rect 3976 9503 4028 9512
rect 3976 9469 3985 9503
rect 3985 9469 4019 9503
rect 4019 9469 4028 9503
rect 4712 9571 4764 9580
rect 4712 9537 4721 9571
rect 4721 9537 4755 9571
rect 4755 9537 4764 9571
rect 4712 9528 4764 9537
rect 3976 9460 4028 9469
rect 5264 9528 5316 9580
rect 7472 9639 7524 9648
rect 7472 9605 7481 9639
rect 7481 9605 7515 9639
rect 7515 9605 7524 9639
rect 7472 9596 7524 9605
rect 8208 9596 8260 9648
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 6644 9460 6696 9512
rect 7932 9503 7984 9512
rect 7932 9469 7941 9503
rect 7941 9469 7975 9503
rect 7975 9469 7984 9503
rect 7932 9460 7984 9469
rect 8116 9571 8168 9580
rect 8116 9537 8125 9571
rect 8125 9537 8159 9571
rect 8159 9537 8168 9571
rect 8116 9528 8168 9537
rect 14648 9596 14700 9648
rect 15844 9596 15896 9648
rect 12900 9571 12952 9580
rect 12900 9537 12909 9571
rect 12909 9537 12943 9571
rect 12943 9537 12952 9571
rect 12900 9528 12952 9537
rect 12992 9571 13044 9580
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 13268 9571 13320 9580
rect 13268 9537 13277 9571
rect 13277 9537 13311 9571
rect 13311 9537 13320 9571
rect 13268 9528 13320 9537
rect 10048 9460 10100 9512
rect 15200 9528 15252 9580
rect 15292 9571 15344 9580
rect 15292 9537 15301 9571
rect 15301 9537 15335 9571
rect 15335 9537 15344 9571
rect 15292 9528 15344 9537
rect 15384 9571 15436 9580
rect 15384 9537 15393 9571
rect 15393 9537 15427 9571
rect 15427 9537 15436 9571
rect 15384 9528 15436 9537
rect 15568 9571 15620 9580
rect 15568 9537 15577 9571
rect 15577 9537 15611 9571
rect 15611 9537 15620 9571
rect 15568 9528 15620 9537
rect 16120 9571 16172 9580
rect 16120 9537 16129 9571
rect 16129 9537 16163 9571
rect 16163 9537 16172 9571
rect 16120 9528 16172 9537
rect 16856 9528 16908 9580
rect 16948 9460 17000 9512
rect 17592 9460 17644 9512
rect 18236 9503 18288 9512
rect 18236 9469 18245 9503
rect 18245 9469 18279 9503
rect 18279 9469 18288 9503
rect 18236 9460 18288 9469
rect 18328 9503 18380 9512
rect 18328 9469 18337 9503
rect 18337 9469 18371 9503
rect 18371 9469 18380 9503
rect 18328 9460 18380 9469
rect 5172 9435 5224 9444
rect 5172 9401 5181 9435
rect 5181 9401 5215 9435
rect 5215 9401 5224 9435
rect 5172 9392 5224 9401
rect 5356 9392 5408 9444
rect 9680 9392 9732 9444
rect 16856 9392 16908 9444
rect 19432 9528 19484 9580
rect 20720 9596 20772 9648
rect 20628 9528 20680 9580
rect 20904 9528 20956 9580
rect 21456 9528 21508 9580
rect 23296 9528 23348 9580
rect 24216 9571 24268 9580
rect 24216 9537 24225 9571
rect 24225 9537 24259 9571
rect 24259 9537 24268 9571
rect 24216 9528 24268 9537
rect 20996 9460 21048 9512
rect 21364 9503 21416 9512
rect 21364 9469 21373 9503
rect 21373 9469 21407 9503
rect 21407 9469 21416 9503
rect 21364 9460 21416 9469
rect 12440 9324 12492 9376
rect 13360 9324 13412 9376
rect 14924 9367 14976 9376
rect 14924 9333 14933 9367
rect 14933 9333 14967 9367
rect 14967 9333 14976 9367
rect 14924 9324 14976 9333
rect 15016 9324 15068 9376
rect 15752 9324 15804 9376
rect 19708 9392 19760 9444
rect 21088 9392 21140 9444
rect 19432 9324 19484 9376
rect 20812 9324 20864 9376
rect 21180 9367 21232 9376
rect 21180 9333 21189 9367
rect 21189 9333 21223 9367
rect 21223 9333 21232 9367
rect 21180 9324 21232 9333
rect 23480 9324 23532 9376
rect 23848 9324 23900 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 4712 9120 4764 9172
rect 8208 9120 8260 9172
rect 11796 9120 11848 9172
rect 15384 9120 15436 9172
rect 18696 9120 18748 9172
rect 21180 9120 21232 9172
rect 2688 8916 2740 8968
rect 3884 8984 3936 9036
rect 5264 9052 5316 9104
rect 12072 9052 12124 9104
rect 5172 9027 5224 9036
rect 5172 8993 5181 9027
rect 5181 8993 5215 9027
rect 5215 8993 5224 9027
rect 5172 8984 5224 8993
rect 11060 8984 11112 9036
rect 18236 8984 18288 9036
rect 3976 8959 4028 8968
rect 3976 8925 3985 8959
rect 3985 8925 4019 8959
rect 4019 8925 4028 8959
rect 3976 8916 4028 8925
rect 4712 8916 4764 8968
rect 5448 8916 5500 8968
rect 7932 8959 7984 8968
rect 7932 8925 7941 8959
rect 7941 8925 7975 8959
rect 7975 8925 7984 8959
rect 7932 8916 7984 8925
rect 8116 8959 8168 8968
rect 8116 8925 8125 8959
rect 8125 8925 8159 8959
rect 8159 8925 8168 8959
rect 8116 8916 8168 8925
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 12716 8959 12768 8968
rect 12716 8925 12725 8959
rect 12725 8925 12759 8959
rect 12759 8925 12768 8959
rect 12716 8916 12768 8925
rect 12808 8959 12860 8968
rect 12808 8925 12817 8959
rect 12817 8925 12851 8959
rect 12851 8925 12860 8959
rect 12808 8916 12860 8925
rect 18512 8959 18564 8968
rect 18512 8925 18521 8959
rect 18521 8925 18555 8959
rect 18555 8925 18564 8959
rect 18512 8916 18564 8925
rect 19432 8959 19484 8968
rect 19432 8925 19441 8959
rect 19441 8925 19475 8959
rect 19475 8925 19484 8959
rect 19432 8916 19484 8925
rect 20720 8959 20772 8968
rect 20720 8925 20729 8959
rect 20729 8925 20763 8959
rect 20763 8925 20772 8959
rect 20720 8916 20772 8925
rect 20812 8959 20864 8968
rect 20812 8925 20821 8959
rect 20821 8925 20855 8959
rect 20855 8925 20864 8959
rect 20812 8916 20864 8925
rect 20996 8959 21048 8968
rect 20996 8925 21005 8959
rect 21005 8925 21039 8959
rect 21039 8925 21048 8959
rect 20996 8916 21048 8925
rect 23480 8959 23532 8968
rect 23480 8925 23489 8959
rect 23489 8925 23523 8959
rect 23523 8925 23532 8959
rect 23480 8916 23532 8925
rect 23664 8959 23716 8968
rect 23664 8925 23673 8959
rect 23673 8925 23707 8959
rect 23707 8925 23716 8959
rect 23664 8916 23716 8925
rect 25044 8916 25096 8968
rect 5356 8848 5408 8900
rect 10140 8848 10192 8900
rect 12072 8848 12124 8900
rect 12348 8891 12400 8900
rect 12348 8857 12357 8891
rect 12357 8857 12391 8891
rect 12391 8857 12400 8891
rect 12348 8848 12400 8857
rect 16856 8848 16908 8900
rect 17776 8848 17828 8900
rect 19708 8848 19760 8900
rect 5540 8780 5592 8832
rect 6920 8780 6972 8832
rect 23296 8780 23348 8832
rect 24308 8848 24360 8900
rect 23940 8780 23992 8832
rect 24768 8780 24820 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 3976 8576 4028 8628
rect 5448 8619 5500 8628
rect 5448 8585 5457 8619
rect 5457 8585 5491 8619
rect 5491 8585 5500 8619
rect 5448 8576 5500 8585
rect 6920 8576 6972 8628
rect 4620 8508 4672 8560
rect 5264 8508 5316 8560
rect 2964 8415 3016 8424
rect 2964 8381 2973 8415
rect 2973 8381 3007 8415
rect 3007 8381 3016 8415
rect 2964 8372 3016 8381
rect 3884 8440 3936 8492
rect 5356 8483 5408 8492
rect 5356 8449 5365 8483
rect 5365 8449 5399 8483
rect 5399 8449 5408 8483
rect 5356 8440 5408 8449
rect 7932 8576 7984 8628
rect 8392 8576 8444 8628
rect 10140 8619 10192 8628
rect 10140 8585 10149 8619
rect 10149 8585 10183 8619
rect 10183 8585 10192 8619
rect 10140 8576 10192 8585
rect 10784 8576 10836 8628
rect 11888 8619 11940 8628
rect 11888 8585 11897 8619
rect 11897 8585 11931 8619
rect 11931 8585 11940 8619
rect 11888 8576 11940 8585
rect 14924 8576 14976 8628
rect 7012 8483 7064 8492
rect 7012 8449 7021 8483
rect 7021 8449 7055 8483
rect 7055 8449 7064 8483
rect 7012 8440 7064 8449
rect 7104 8483 7156 8492
rect 7104 8449 7113 8483
rect 7113 8449 7147 8483
rect 7147 8449 7156 8483
rect 7104 8440 7156 8449
rect 7472 8483 7524 8492
rect 7472 8449 7481 8483
rect 7481 8449 7515 8483
rect 7515 8449 7524 8483
rect 7472 8440 7524 8449
rect 11060 8508 11112 8560
rect 17132 8576 17184 8628
rect 18328 8576 18380 8628
rect 22928 8576 22980 8628
rect 24124 8576 24176 8628
rect 24676 8576 24728 8628
rect 24768 8576 24820 8628
rect 7012 8304 7064 8356
rect 8024 8483 8076 8492
rect 8024 8449 8033 8483
rect 8033 8449 8067 8483
rect 8067 8449 8076 8483
rect 8024 8440 8076 8449
rect 9128 8483 9180 8492
rect 9128 8449 9137 8483
rect 9137 8449 9171 8483
rect 9171 8449 9180 8483
rect 9128 8440 9180 8449
rect 9312 8483 9364 8492
rect 9312 8449 9321 8483
rect 9321 8449 9355 8483
rect 9355 8449 9364 8483
rect 9312 8440 9364 8449
rect 10048 8483 10100 8492
rect 10048 8449 10057 8483
rect 10057 8449 10091 8483
rect 10091 8449 10100 8483
rect 10048 8440 10100 8449
rect 10508 8440 10560 8492
rect 10784 8483 10836 8492
rect 10784 8449 10793 8483
rect 10793 8449 10827 8483
rect 10827 8449 10836 8483
rect 10784 8440 10836 8449
rect 11796 8483 11848 8492
rect 11796 8449 11805 8483
rect 11805 8449 11839 8483
rect 11839 8449 11848 8483
rect 11796 8440 11848 8449
rect 11980 8483 12032 8492
rect 11980 8449 11989 8483
rect 11989 8449 12023 8483
rect 12023 8449 12032 8483
rect 11980 8440 12032 8449
rect 12348 8440 12400 8492
rect 10600 8372 10652 8424
rect 23296 8551 23348 8560
rect 23296 8517 23305 8551
rect 23305 8517 23339 8551
rect 23339 8517 23348 8551
rect 23296 8508 23348 8517
rect 25044 8508 25096 8560
rect 17592 8440 17644 8492
rect 18052 8440 18104 8492
rect 17776 8415 17828 8424
rect 17776 8381 17785 8415
rect 17785 8381 17819 8415
rect 17819 8381 17828 8415
rect 17776 8372 17828 8381
rect 23388 8483 23440 8492
rect 23388 8449 23397 8483
rect 23397 8449 23431 8483
rect 23431 8449 23440 8483
rect 23388 8440 23440 8449
rect 23572 8483 23624 8492
rect 23572 8449 23581 8483
rect 23581 8449 23615 8483
rect 23615 8449 23624 8483
rect 23572 8440 23624 8449
rect 23848 8440 23900 8492
rect 23940 8483 23992 8492
rect 23940 8449 23949 8483
rect 23949 8449 23983 8483
rect 23983 8449 23992 8483
rect 23940 8440 23992 8449
rect 24032 8372 24084 8424
rect 24308 8483 24360 8492
rect 24308 8449 24317 8483
rect 24317 8449 24351 8483
rect 24351 8449 24360 8483
rect 24308 8440 24360 8449
rect 25228 8483 25280 8492
rect 25228 8449 25237 8483
rect 25237 8449 25271 8483
rect 25271 8449 25280 8483
rect 25228 8440 25280 8449
rect 27712 8440 27764 8492
rect 9680 8304 9732 8356
rect 15200 8304 15252 8356
rect 4712 8236 4764 8288
rect 7472 8236 7524 8288
rect 17132 8304 17184 8356
rect 17040 8279 17092 8288
rect 17040 8245 17049 8279
rect 17049 8245 17083 8279
rect 17083 8245 17092 8279
rect 17040 8236 17092 8245
rect 17408 8279 17460 8288
rect 17408 8245 17417 8279
rect 17417 8245 17451 8279
rect 17451 8245 17460 8279
rect 17408 8236 17460 8245
rect 18880 8236 18932 8288
rect 21088 8304 21140 8356
rect 23756 8347 23808 8356
rect 23756 8313 23765 8347
rect 23765 8313 23799 8347
rect 23799 8313 23808 8347
rect 23756 8304 23808 8313
rect 24676 8372 24728 8424
rect 24308 8304 24360 8356
rect 24124 8279 24176 8288
rect 24124 8245 24133 8279
rect 24133 8245 24167 8279
rect 24167 8245 24176 8279
rect 24124 8236 24176 8245
rect 24216 8236 24268 8288
rect 24676 8279 24728 8288
rect 24676 8245 24685 8279
rect 24685 8245 24719 8279
rect 24719 8245 24728 8279
rect 24676 8236 24728 8245
rect 25136 8304 25188 8356
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 9128 8032 9180 8084
rect 9312 8075 9364 8084
rect 9312 8041 9321 8075
rect 9321 8041 9355 8075
rect 9355 8041 9364 8075
rect 9312 8032 9364 8041
rect 11980 8075 12032 8084
rect 11980 8041 11989 8075
rect 11989 8041 12023 8075
rect 12023 8041 12032 8075
rect 11980 8032 12032 8041
rect 12716 8075 12768 8084
rect 12716 8041 12725 8075
rect 12725 8041 12759 8075
rect 12759 8041 12768 8075
rect 12716 8032 12768 8041
rect 15384 8075 15436 8084
rect 15384 8041 15393 8075
rect 15393 8041 15427 8075
rect 15427 8041 15436 8075
rect 15384 8032 15436 8041
rect 15844 8075 15896 8084
rect 15844 8041 15853 8075
rect 15853 8041 15887 8075
rect 15887 8041 15896 8075
rect 15844 8032 15896 8041
rect 16580 8032 16632 8084
rect 5632 7964 5684 8016
rect 3884 7939 3936 7948
rect 3884 7905 3893 7939
rect 3893 7905 3927 7939
rect 3927 7905 3936 7939
rect 3884 7896 3936 7905
rect 4528 7896 4580 7948
rect 4712 7939 4764 7948
rect 4712 7905 4721 7939
rect 4721 7905 4755 7939
rect 4755 7905 4764 7939
rect 4712 7896 4764 7905
rect 6920 7939 6972 7948
rect 6920 7905 6929 7939
rect 6929 7905 6963 7939
rect 6963 7905 6972 7939
rect 6920 7896 6972 7905
rect 8024 7964 8076 8016
rect 11796 7964 11848 8016
rect 18328 8032 18380 8084
rect 4344 7828 4396 7880
rect 7196 7828 7248 7880
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 11980 7896 12032 7948
rect 8576 7828 8628 7837
rect 10784 7828 10836 7880
rect 10140 7760 10192 7812
rect 12716 7828 12768 7880
rect 17868 7964 17920 8016
rect 18420 7964 18472 8016
rect 19248 7964 19300 8016
rect 13360 7896 13412 7948
rect 14464 7896 14516 7948
rect 13268 7871 13320 7880
rect 13268 7837 13277 7871
rect 13277 7837 13311 7871
rect 13311 7837 13320 7871
rect 13268 7828 13320 7837
rect 15200 7828 15252 7880
rect 15568 7871 15620 7880
rect 15568 7837 15577 7871
rect 15577 7837 15611 7871
rect 15611 7837 15620 7871
rect 15568 7828 15620 7837
rect 15660 7871 15712 7880
rect 15660 7837 15669 7871
rect 15669 7837 15703 7871
rect 15703 7837 15712 7871
rect 15660 7828 15712 7837
rect 17040 7939 17092 7948
rect 17040 7905 17049 7939
rect 17049 7905 17083 7939
rect 17083 7905 17092 7939
rect 17040 7896 17092 7905
rect 14280 7760 14332 7812
rect 17408 7828 17460 7880
rect 18052 7871 18104 7880
rect 18052 7837 18061 7871
rect 18061 7837 18095 7871
rect 18095 7837 18104 7871
rect 18052 7828 18104 7837
rect 18144 7871 18196 7880
rect 18144 7837 18153 7871
rect 18153 7837 18187 7871
rect 18187 7837 18196 7871
rect 18144 7828 18196 7837
rect 18328 7871 18380 7880
rect 18328 7837 18337 7871
rect 18337 7837 18371 7871
rect 18371 7837 18380 7871
rect 18328 7828 18380 7837
rect 18420 7871 18472 7880
rect 18420 7837 18429 7871
rect 18429 7837 18463 7871
rect 18463 7837 18472 7871
rect 18420 7828 18472 7837
rect 18512 7828 18564 7880
rect 5448 7692 5500 7744
rect 12256 7692 12308 7744
rect 13820 7692 13872 7744
rect 15016 7692 15068 7744
rect 17316 7692 17368 7744
rect 17684 7760 17736 7812
rect 18512 7692 18564 7744
rect 18604 7735 18656 7744
rect 18604 7701 18613 7735
rect 18613 7701 18647 7735
rect 18647 7701 18656 7735
rect 18604 7692 18656 7701
rect 19248 7871 19300 7880
rect 19248 7837 19257 7871
rect 19257 7837 19291 7871
rect 19291 7837 19300 7871
rect 19248 7828 19300 7837
rect 20076 7896 20128 7948
rect 19708 7871 19760 7880
rect 19708 7837 19717 7871
rect 19717 7837 19751 7871
rect 19751 7837 19760 7871
rect 19708 7828 19760 7837
rect 20444 7828 20496 7880
rect 20536 7871 20588 7880
rect 20536 7837 20545 7871
rect 20545 7837 20579 7871
rect 20579 7837 20588 7871
rect 20536 7828 20588 7837
rect 21364 7964 21416 8016
rect 21824 8032 21876 8084
rect 22560 8032 22612 8084
rect 24032 8032 24084 8084
rect 25044 8032 25096 8084
rect 22928 7964 22980 8016
rect 21640 7896 21692 7948
rect 22008 7896 22060 7948
rect 20812 7871 20864 7880
rect 20812 7837 20821 7871
rect 20821 7837 20855 7871
rect 20855 7837 20864 7871
rect 20812 7828 20864 7837
rect 20904 7871 20956 7880
rect 20904 7837 20913 7871
rect 20913 7837 20947 7871
rect 20947 7837 20956 7871
rect 20904 7828 20956 7837
rect 21180 7871 21232 7880
rect 21180 7837 21189 7871
rect 21189 7837 21223 7871
rect 21223 7837 21232 7871
rect 21180 7828 21232 7837
rect 21364 7871 21416 7880
rect 21364 7837 21373 7871
rect 21373 7837 21407 7871
rect 21407 7837 21416 7871
rect 21364 7828 21416 7837
rect 21456 7871 21508 7880
rect 21456 7837 21465 7871
rect 21465 7837 21499 7871
rect 21499 7837 21508 7871
rect 21456 7828 21508 7837
rect 22744 7828 22796 7880
rect 23388 7828 23440 7880
rect 23848 7871 23900 7880
rect 23848 7837 23857 7871
rect 23857 7837 23891 7871
rect 23891 7837 23900 7871
rect 23848 7828 23900 7837
rect 24400 7939 24452 7948
rect 24400 7905 24409 7939
rect 24409 7905 24443 7939
rect 24443 7905 24452 7939
rect 24400 7896 24452 7905
rect 24676 7939 24728 7948
rect 24676 7905 24685 7939
rect 24685 7905 24719 7939
rect 24719 7905 24728 7939
rect 24676 7896 24728 7905
rect 24124 7871 24176 7880
rect 24124 7837 24133 7871
rect 24133 7837 24167 7871
rect 24167 7837 24176 7871
rect 24124 7828 24176 7837
rect 19984 7760 20036 7812
rect 20168 7760 20220 7812
rect 21732 7803 21784 7812
rect 21732 7769 21741 7803
rect 21741 7769 21775 7803
rect 21775 7769 21784 7803
rect 21732 7760 21784 7769
rect 22652 7803 22704 7812
rect 22652 7769 22661 7803
rect 22661 7769 22695 7803
rect 22695 7769 22704 7803
rect 22652 7760 22704 7769
rect 25136 7760 25188 7812
rect 19248 7692 19300 7744
rect 20260 7692 20312 7744
rect 20812 7692 20864 7744
rect 21088 7692 21140 7744
rect 21824 7735 21876 7744
rect 21824 7701 21833 7735
rect 21833 7701 21867 7735
rect 21867 7701 21876 7735
rect 21824 7692 21876 7701
rect 23020 7735 23072 7744
rect 23020 7701 23029 7735
rect 23029 7701 23063 7735
rect 23063 7701 23072 7735
rect 23020 7692 23072 7701
rect 23480 7735 23532 7744
rect 23480 7701 23489 7735
rect 23489 7701 23523 7735
rect 23523 7701 23532 7735
rect 23480 7692 23532 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 4344 7531 4396 7540
rect 4344 7497 4353 7531
rect 4353 7497 4387 7531
rect 4387 7497 4396 7531
rect 4344 7488 4396 7497
rect 7288 7488 7340 7540
rect 8392 7420 8444 7472
rect 9588 7488 9640 7540
rect 14188 7488 14240 7540
rect 15568 7488 15620 7540
rect 17500 7488 17552 7540
rect 18512 7488 18564 7540
rect 9772 7463 9824 7472
rect 9772 7429 9781 7463
rect 9781 7429 9815 7463
rect 9815 7429 9824 7463
rect 9772 7420 9824 7429
rect 10048 7420 10100 7472
rect 5264 7352 5316 7404
rect 6276 7352 6328 7404
rect 5540 7284 5592 7336
rect 5632 7284 5684 7336
rect 6920 7395 6972 7404
rect 6920 7361 6929 7395
rect 6929 7361 6963 7395
rect 6963 7361 6972 7395
rect 6920 7352 6972 7361
rect 8208 7352 8260 7404
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 9404 7395 9456 7404
rect 9404 7361 9413 7395
rect 9413 7361 9447 7395
rect 9447 7361 9456 7395
rect 9404 7352 9456 7361
rect 8576 7284 8628 7336
rect 10324 7352 10376 7404
rect 10784 7395 10836 7404
rect 10784 7361 10793 7395
rect 10793 7361 10827 7395
rect 10827 7361 10836 7395
rect 10784 7352 10836 7361
rect 10968 7395 11020 7404
rect 10968 7361 10977 7395
rect 10977 7361 11011 7395
rect 11011 7361 11020 7395
rect 10968 7352 11020 7361
rect 11060 7395 11112 7404
rect 11060 7361 11069 7395
rect 11069 7361 11103 7395
rect 11103 7361 11112 7395
rect 11060 7352 11112 7361
rect 11796 7420 11848 7472
rect 11980 7395 12032 7404
rect 11980 7361 11989 7395
rect 11989 7361 12023 7395
rect 12023 7361 12032 7395
rect 12900 7420 12952 7472
rect 14280 7420 14332 7472
rect 11980 7352 12032 7361
rect 12624 7352 12676 7404
rect 13268 7352 13320 7404
rect 14556 7352 14608 7404
rect 14740 7395 14792 7404
rect 14740 7361 14749 7395
rect 14749 7361 14783 7395
rect 14783 7361 14792 7395
rect 14740 7352 14792 7361
rect 14832 7395 14884 7404
rect 14832 7361 14841 7395
rect 14841 7361 14875 7395
rect 14875 7361 14884 7395
rect 14832 7352 14884 7361
rect 15384 7420 15436 7472
rect 16120 7420 16172 7472
rect 18052 7420 18104 7472
rect 18788 7420 18840 7472
rect 11888 7259 11940 7268
rect 11888 7225 11897 7259
rect 11897 7225 11931 7259
rect 11931 7225 11940 7259
rect 11888 7216 11940 7225
rect 5908 7148 5960 7200
rect 9772 7148 9824 7200
rect 12716 7216 12768 7268
rect 12992 7216 13044 7268
rect 13360 7216 13412 7268
rect 14648 7327 14700 7336
rect 14648 7293 14657 7327
rect 14657 7293 14691 7327
rect 14691 7293 14700 7327
rect 14648 7284 14700 7293
rect 15752 7284 15804 7336
rect 16764 7284 16816 7336
rect 17592 7352 17644 7404
rect 17960 7352 18012 7404
rect 18604 7395 18656 7404
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 21088 7488 21140 7540
rect 21364 7488 21416 7540
rect 21916 7488 21968 7540
rect 24216 7488 24268 7540
rect 20168 7352 20220 7404
rect 20352 7395 20404 7404
rect 20352 7361 20361 7395
rect 20361 7361 20395 7395
rect 20395 7361 20404 7395
rect 20352 7352 20404 7361
rect 20444 7395 20496 7404
rect 20444 7361 20453 7395
rect 20453 7361 20487 7395
rect 20487 7361 20496 7395
rect 20444 7352 20496 7361
rect 20536 7395 20588 7404
rect 20536 7361 20545 7395
rect 20545 7361 20579 7395
rect 20579 7361 20588 7395
rect 20536 7352 20588 7361
rect 18880 7327 18932 7336
rect 18880 7293 18889 7327
rect 18889 7293 18923 7327
rect 18923 7293 18932 7327
rect 18880 7284 18932 7293
rect 19708 7284 19760 7336
rect 20260 7284 20312 7336
rect 20812 7395 20864 7404
rect 20812 7361 20821 7395
rect 20821 7361 20855 7395
rect 20855 7361 20864 7395
rect 20812 7352 20864 7361
rect 20996 7352 21048 7404
rect 21548 7352 21600 7404
rect 12532 7191 12584 7200
rect 12532 7157 12541 7191
rect 12541 7157 12575 7191
rect 12575 7157 12584 7191
rect 12532 7148 12584 7157
rect 12808 7148 12860 7200
rect 14372 7148 14424 7200
rect 18052 7148 18104 7200
rect 19984 7259 20036 7268
rect 19984 7225 19993 7259
rect 19993 7225 20027 7259
rect 20027 7225 20036 7259
rect 19984 7216 20036 7225
rect 20076 7259 20128 7268
rect 20076 7225 20085 7259
rect 20085 7225 20119 7259
rect 20119 7225 20128 7259
rect 20076 7216 20128 7225
rect 20720 7216 20772 7268
rect 20904 7216 20956 7268
rect 22744 7463 22796 7472
rect 22744 7429 22753 7463
rect 22753 7429 22787 7463
rect 22787 7429 22796 7463
rect 22744 7420 22796 7429
rect 22928 7463 22980 7472
rect 22928 7429 22937 7463
rect 22937 7429 22971 7463
rect 22971 7429 22980 7463
rect 22928 7420 22980 7429
rect 22008 7395 22060 7404
rect 22008 7361 22017 7395
rect 22017 7361 22051 7395
rect 22051 7361 22060 7395
rect 22008 7352 22060 7361
rect 22560 7352 22612 7404
rect 22560 7216 22612 7268
rect 19340 7148 19392 7200
rect 19708 7148 19760 7200
rect 24216 7395 24268 7404
rect 24216 7361 24225 7395
rect 24225 7361 24259 7395
rect 24259 7361 24268 7395
rect 24216 7352 24268 7361
rect 24308 7395 24360 7404
rect 24308 7361 24317 7395
rect 24317 7361 24351 7395
rect 24351 7361 24360 7395
rect 24308 7352 24360 7361
rect 23388 7327 23440 7336
rect 23388 7293 23397 7327
rect 23397 7293 23431 7327
rect 23431 7293 23440 7327
rect 23388 7284 23440 7293
rect 24124 7284 24176 7336
rect 27620 7216 27672 7268
rect 24032 7191 24084 7200
rect 24032 7157 24041 7191
rect 24041 7157 24075 7191
rect 24075 7157 24084 7191
rect 24032 7148 24084 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 5540 6944 5592 6996
rect 5448 6919 5500 6928
rect 5448 6885 5457 6919
rect 5457 6885 5491 6919
rect 5491 6885 5500 6919
rect 5448 6876 5500 6885
rect 5632 6808 5684 6860
rect 5816 6740 5868 6792
rect 6276 6851 6328 6860
rect 6276 6817 6285 6851
rect 6285 6817 6319 6851
rect 6319 6817 6328 6851
rect 6276 6808 6328 6817
rect 8576 6944 8628 6996
rect 9404 6944 9456 6996
rect 10508 6944 10560 6996
rect 10784 6987 10836 6996
rect 10784 6953 10793 6987
rect 10793 6953 10827 6987
rect 10827 6953 10836 6987
rect 10784 6944 10836 6953
rect 6460 6808 6512 6860
rect 6644 6740 6696 6792
rect 7104 6740 7156 6792
rect 8208 6783 8260 6792
rect 8208 6749 8217 6783
rect 8217 6749 8251 6783
rect 8251 6749 8260 6783
rect 8208 6740 8260 6749
rect 8392 6783 8444 6792
rect 8392 6749 8401 6783
rect 8401 6749 8435 6783
rect 8435 6749 8444 6783
rect 8392 6740 8444 6749
rect 9128 6783 9180 6792
rect 6920 6672 6972 6724
rect 7564 6715 7616 6724
rect 7564 6681 7573 6715
rect 7573 6681 7607 6715
rect 7607 6681 7616 6715
rect 7564 6672 7616 6681
rect 6644 6604 6696 6656
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 10048 6876 10100 6928
rect 10140 6740 10192 6792
rect 11060 6808 11112 6860
rect 11244 6876 11296 6928
rect 11888 6876 11940 6928
rect 11428 6740 11480 6792
rect 10324 6672 10376 6724
rect 11152 6715 11204 6724
rect 11152 6681 11161 6715
rect 11161 6681 11195 6715
rect 11195 6681 11204 6715
rect 11152 6672 11204 6681
rect 11704 6740 11756 6792
rect 11796 6783 11848 6792
rect 11796 6749 11805 6783
rect 11805 6749 11839 6783
rect 11839 6749 11848 6783
rect 11796 6740 11848 6749
rect 14280 6987 14332 6996
rect 14280 6953 14289 6987
rect 14289 6953 14323 6987
rect 14323 6953 14332 6987
rect 14280 6944 14332 6953
rect 13084 6876 13136 6928
rect 12256 6808 12308 6860
rect 12348 6808 12400 6860
rect 12624 6808 12676 6860
rect 12164 6740 12216 6792
rect 12808 6783 12860 6792
rect 12808 6749 12817 6783
rect 12817 6749 12851 6783
rect 12851 6749 12860 6783
rect 12808 6740 12860 6749
rect 13360 6876 13412 6928
rect 14740 6808 14792 6860
rect 14832 6808 14884 6860
rect 13360 6783 13412 6792
rect 13360 6749 13369 6783
rect 13369 6749 13403 6783
rect 13403 6749 13412 6783
rect 13360 6740 13412 6749
rect 13452 6783 13504 6792
rect 13452 6749 13461 6783
rect 13461 6749 13495 6783
rect 13495 6749 13504 6783
rect 13452 6740 13504 6749
rect 14096 6740 14148 6792
rect 14556 6783 14608 6792
rect 14556 6749 14565 6783
rect 14565 6749 14599 6783
rect 14599 6749 14608 6783
rect 14556 6740 14608 6749
rect 17684 6944 17736 6996
rect 17868 6944 17920 6996
rect 12348 6672 12400 6724
rect 13636 6715 13688 6724
rect 13636 6681 13645 6715
rect 13645 6681 13679 6715
rect 13679 6681 13688 6715
rect 13636 6672 13688 6681
rect 13820 6672 13872 6724
rect 14740 6715 14792 6724
rect 14740 6681 14749 6715
rect 14749 6681 14783 6715
rect 14783 6681 14792 6715
rect 14740 6672 14792 6681
rect 9496 6647 9548 6656
rect 9496 6613 9505 6647
rect 9505 6613 9539 6647
rect 9539 6613 9548 6647
rect 9496 6604 9548 6613
rect 10968 6604 11020 6656
rect 11612 6604 11664 6656
rect 11704 6604 11756 6656
rect 13360 6604 13412 6656
rect 13544 6604 13596 6656
rect 16212 6876 16264 6928
rect 16764 6851 16816 6860
rect 16764 6817 16773 6851
rect 16773 6817 16807 6851
rect 16807 6817 16816 6851
rect 16764 6808 16816 6817
rect 15660 6783 15712 6792
rect 15660 6749 15669 6783
rect 15669 6749 15703 6783
rect 15703 6749 15712 6783
rect 15660 6740 15712 6749
rect 15752 6783 15804 6792
rect 15752 6749 15761 6783
rect 15761 6749 15795 6783
rect 15795 6749 15804 6783
rect 15752 6740 15804 6749
rect 15844 6783 15896 6792
rect 15844 6749 15853 6783
rect 15853 6749 15887 6783
rect 15887 6749 15896 6783
rect 15844 6740 15896 6749
rect 16672 6783 16724 6792
rect 16672 6749 16681 6783
rect 16681 6749 16715 6783
rect 16715 6749 16724 6783
rect 16672 6740 16724 6749
rect 17040 6783 17092 6792
rect 17040 6749 17049 6783
rect 17049 6749 17083 6783
rect 17083 6749 17092 6783
rect 17040 6740 17092 6749
rect 17316 6783 17368 6792
rect 17316 6749 17325 6783
rect 17325 6749 17359 6783
rect 17359 6749 17368 6783
rect 17316 6740 17368 6749
rect 18420 6876 18472 6928
rect 18788 6987 18840 6996
rect 18788 6953 18797 6987
rect 18797 6953 18831 6987
rect 18831 6953 18840 6987
rect 18788 6944 18840 6953
rect 19340 6944 19392 6996
rect 21548 6987 21600 6996
rect 21548 6953 21557 6987
rect 21557 6953 21591 6987
rect 21591 6953 21600 6987
rect 21548 6944 21600 6953
rect 21732 6944 21784 6996
rect 23480 6944 23532 6996
rect 24308 6944 24360 6996
rect 19708 6876 19760 6928
rect 17776 6783 17828 6792
rect 17776 6749 17785 6783
rect 17785 6749 17819 6783
rect 17819 6749 17828 6783
rect 17776 6740 17828 6749
rect 18144 6808 18196 6860
rect 24400 6808 24452 6860
rect 18052 6783 18104 6792
rect 18052 6749 18061 6783
rect 18061 6749 18095 6783
rect 18095 6749 18104 6783
rect 18052 6740 18104 6749
rect 18328 6783 18380 6792
rect 18328 6749 18337 6783
rect 18337 6749 18371 6783
rect 18371 6749 18380 6783
rect 18328 6740 18380 6749
rect 18420 6740 18472 6792
rect 18788 6740 18840 6792
rect 19248 6740 19300 6792
rect 19432 6783 19484 6792
rect 19432 6749 19441 6783
rect 19441 6749 19475 6783
rect 19475 6749 19484 6783
rect 19432 6740 19484 6749
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 15108 6647 15160 6656
rect 15108 6613 15117 6647
rect 15117 6613 15151 6647
rect 15151 6613 15160 6647
rect 15108 6604 15160 6613
rect 16672 6604 16724 6656
rect 22008 6783 22060 6792
rect 22008 6749 22017 6783
rect 22017 6749 22051 6783
rect 22051 6749 22060 6783
rect 22008 6740 22060 6749
rect 20812 6604 20864 6656
rect 25136 6672 25188 6724
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 6460 6400 6512 6452
rect 7104 6400 7156 6452
rect 11060 6400 11112 6452
rect 12164 6400 12216 6452
rect 13176 6400 13228 6452
rect 14832 6443 14884 6452
rect 14832 6409 14841 6443
rect 14841 6409 14875 6443
rect 14875 6409 14884 6443
rect 14832 6400 14884 6409
rect 15752 6400 15804 6452
rect 17500 6400 17552 6452
rect 17868 6400 17920 6452
rect 19248 6400 19300 6452
rect 19432 6400 19484 6452
rect 20536 6400 20588 6452
rect 20904 6400 20956 6452
rect 22008 6400 22060 6452
rect 27620 6443 27672 6452
rect 27620 6409 27629 6443
rect 27629 6409 27663 6443
rect 27663 6409 27672 6443
rect 27620 6400 27672 6409
rect 7196 6332 7248 6384
rect 11980 6332 12032 6384
rect 12716 6332 12768 6384
rect 5448 6264 5500 6316
rect 6460 6307 6512 6316
rect 6460 6273 6469 6307
rect 6469 6273 6503 6307
rect 6503 6273 6512 6307
rect 6460 6264 6512 6273
rect 6644 6264 6696 6316
rect 7288 6307 7340 6316
rect 7288 6273 7297 6307
rect 7297 6273 7331 6307
rect 7331 6273 7340 6307
rect 7288 6264 7340 6273
rect 9496 6264 9548 6316
rect 5908 6239 5960 6248
rect 5908 6205 5917 6239
rect 5917 6205 5951 6239
rect 5951 6205 5960 6239
rect 5908 6196 5960 6205
rect 6276 6196 6328 6248
rect 8392 6196 8444 6248
rect 12440 6264 12492 6316
rect 12900 6307 12952 6316
rect 12900 6273 12909 6307
rect 12909 6273 12943 6307
rect 12943 6273 12952 6307
rect 14280 6332 14332 6384
rect 14556 6332 14608 6384
rect 12900 6264 12952 6273
rect 12992 6196 13044 6248
rect 13820 6128 13872 6180
rect 15108 6307 15160 6316
rect 15108 6273 15117 6307
rect 15117 6273 15151 6307
rect 15151 6273 15160 6307
rect 15108 6264 15160 6273
rect 15384 6307 15436 6316
rect 15384 6273 15393 6307
rect 15393 6273 15427 6307
rect 15427 6273 15436 6307
rect 15384 6264 15436 6273
rect 16396 6264 16448 6316
rect 21548 6264 21600 6316
rect 23020 6264 23072 6316
rect 27804 6307 27856 6316
rect 27804 6273 27813 6307
rect 27813 6273 27847 6307
rect 27847 6273 27856 6307
rect 27804 6264 27856 6273
rect 14556 6239 14608 6248
rect 14556 6205 14565 6239
rect 14565 6205 14599 6239
rect 14599 6205 14608 6239
rect 14556 6196 14608 6205
rect 17224 6196 17276 6248
rect 17684 6196 17736 6248
rect 24032 6196 24084 6248
rect 14280 6128 14332 6180
rect 15844 6128 15896 6180
rect 12348 6103 12400 6112
rect 12348 6069 12357 6103
rect 12357 6069 12391 6103
rect 12391 6069 12400 6103
rect 12348 6060 12400 6069
rect 14648 6103 14700 6112
rect 14648 6069 14657 6103
rect 14657 6069 14691 6103
rect 14691 6069 14700 6103
rect 16580 6128 16632 6180
rect 14648 6060 14700 6069
rect 16396 6060 16448 6112
rect 18420 6060 18472 6112
rect 18696 6060 18748 6112
rect 23020 6060 23072 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 6920 5856 6972 5908
rect 7380 5856 7432 5908
rect 8668 5856 8720 5908
rect 11980 5899 12032 5908
rect 11980 5865 11989 5899
rect 11989 5865 12023 5899
rect 12023 5865 12032 5899
rect 11980 5856 12032 5865
rect 12624 5856 12676 5908
rect 15384 5856 15436 5908
rect 15844 5899 15896 5908
rect 15844 5865 15853 5899
rect 15853 5865 15887 5899
rect 15887 5865 15896 5899
rect 15844 5856 15896 5865
rect 17592 5856 17644 5908
rect 27712 5856 27764 5908
rect 14004 5788 14056 5840
rect 10232 5763 10284 5772
rect 10232 5729 10241 5763
rect 10241 5729 10275 5763
rect 10275 5729 10284 5763
rect 10232 5720 10284 5729
rect 11520 5720 11572 5772
rect 17224 5720 17276 5772
rect 27528 5652 27580 5704
rect 10508 5627 10560 5636
rect 10508 5593 10517 5627
rect 10517 5593 10551 5627
rect 10551 5593 10560 5627
rect 10508 5584 10560 5593
rect 12072 5584 12124 5636
rect 13084 5584 13136 5636
rect 14372 5627 14424 5636
rect 14372 5593 14381 5627
rect 14381 5593 14415 5627
rect 14415 5593 14424 5627
rect 14372 5584 14424 5593
rect 16764 5584 16816 5636
rect 15660 5516 15712 5568
rect 17868 5584 17920 5636
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 12164 5312 12216 5364
rect 13268 5355 13320 5364
rect 13268 5321 13277 5355
rect 13277 5321 13311 5355
rect 13311 5321 13320 5355
rect 13268 5312 13320 5321
rect 13084 5244 13136 5296
rect 15660 5244 15712 5296
rect 11520 5219 11572 5228
rect 11520 5185 11529 5219
rect 11529 5185 11563 5219
rect 11563 5185 11572 5219
rect 11520 5176 11572 5185
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 7564 2592 7616 2644
rect 8668 2635 8720 2644
rect 8668 2601 8677 2635
rect 8677 2601 8711 2635
rect 8711 2601 8720 2635
rect 8668 2592 8720 2601
rect 5816 2388 5868 2440
rect 8392 2388 8444 2440
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 12898 30676 12954 31476
rect 13542 30676 13598 31476
rect 14186 30818 14242 31476
rect 14186 30790 14412 30818
rect 14186 30676 14242 30790
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 12912 28762 12940 30676
rect 13556 28762 13584 30676
rect 14384 28762 14412 30790
rect 14830 30676 14886 31476
rect 15474 30818 15530 31476
rect 15474 30790 15700 30818
rect 15474 30676 15530 30790
rect 14844 28762 14872 30676
rect 15672 28762 15700 30790
rect 16118 30676 16174 31476
rect 16762 30676 16818 31476
rect 17406 30676 17462 31476
rect 18050 30676 18106 31476
rect 18694 30676 18750 31476
rect 19338 30676 19394 31476
rect 19982 30676 20038 31476
rect 20626 30676 20682 31476
rect 21270 30676 21326 31476
rect 21914 30676 21970 31476
rect 22558 30676 22614 31476
rect 23202 30676 23258 31476
rect 23846 30676 23902 31476
rect 24490 30676 24546 31476
rect 25134 30676 25190 31476
rect 25778 30676 25834 31476
rect 26422 30676 26478 31476
rect 27066 30676 27122 31476
rect 27710 30676 27766 31476
rect 28354 30676 28410 31476
rect 28998 30676 29054 31476
rect 16132 28762 16160 30676
rect 16776 28966 16804 30676
rect 16764 28960 16816 28966
rect 16764 28902 16816 28908
rect 17420 28762 17448 30676
rect 17500 28960 17552 28966
rect 17500 28902 17552 28908
rect 12900 28756 12952 28762
rect 12900 28698 12952 28704
rect 13544 28756 13596 28762
rect 13544 28698 13596 28704
rect 14372 28756 14424 28762
rect 14372 28698 14424 28704
rect 14832 28756 14884 28762
rect 14832 28698 14884 28704
rect 15660 28756 15712 28762
rect 15660 28698 15712 28704
rect 16120 28756 16172 28762
rect 16120 28698 16172 28704
rect 17408 28756 17460 28762
rect 17408 28698 17460 28704
rect 17512 28694 17540 28902
rect 18064 28762 18092 30676
rect 18052 28756 18104 28762
rect 18052 28698 18104 28704
rect 18708 28694 18736 30676
rect 19352 28762 19380 30676
rect 19340 28756 19392 28762
rect 19340 28698 19392 28704
rect 19996 28694 20024 30676
rect 20640 28762 20668 30676
rect 20628 28756 20680 28762
rect 20628 28698 20680 28704
rect 21284 28694 21312 30676
rect 21928 28762 21956 30676
rect 22572 28762 22600 30676
rect 23216 28762 23244 30676
rect 23860 28762 23888 30676
rect 21916 28756 21968 28762
rect 21916 28698 21968 28704
rect 22560 28756 22612 28762
rect 22560 28698 22612 28704
rect 23204 28756 23256 28762
rect 23204 28698 23256 28704
rect 23848 28756 23900 28762
rect 23848 28698 23900 28704
rect 24504 28694 24532 30676
rect 25148 28762 25176 30676
rect 25792 28762 25820 30676
rect 26436 28762 26464 30676
rect 25136 28756 25188 28762
rect 25136 28698 25188 28704
rect 25780 28756 25832 28762
rect 25780 28698 25832 28704
rect 26424 28756 26476 28762
rect 26424 28698 26476 28704
rect 17224 28688 17276 28694
rect 17224 28630 17276 28636
rect 17500 28688 17552 28694
rect 17500 28630 17552 28636
rect 18696 28688 18748 28694
rect 18696 28630 18748 28636
rect 19984 28688 20036 28694
rect 19984 28630 20036 28636
rect 21272 28688 21324 28694
rect 21272 28630 21324 28636
rect 24492 28688 24544 28694
rect 24492 28630 24544 28636
rect 17132 28552 17184 28558
rect 17132 28494 17184 28500
rect 13268 28484 13320 28490
rect 13268 28426 13320 28432
rect 14648 28484 14700 28490
rect 14648 28426 14700 28432
rect 16856 28484 16908 28490
rect 16856 28426 16908 28432
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 13280 28150 13308 28426
rect 10140 28144 10192 28150
rect 10140 28086 10192 28092
rect 13268 28144 13320 28150
rect 13268 28086 13320 28092
rect 6368 28076 6420 28082
rect 6368 28018 6420 28024
rect 6920 28076 6972 28082
rect 6920 28018 6972 28024
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 6380 27674 6408 28018
rect 6460 27872 6512 27878
rect 6460 27814 6512 27820
rect 6368 27668 6420 27674
rect 6368 27610 6420 27616
rect 5448 27600 5500 27606
rect 5448 27542 5500 27548
rect 2228 27532 2280 27538
rect 2228 27474 2280 27480
rect 5264 27532 5316 27538
rect 5264 27474 5316 27480
rect 2240 26994 2268 27474
rect 3884 27464 3936 27470
rect 3884 27406 3936 27412
rect 3976 27464 4028 27470
rect 3976 27406 4028 27412
rect 4804 27464 4856 27470
rect 4804 27406 4856 27412
rect 3700 27396 3752 27402
rect 3700 27338 3752 27344
rect 3148 27056 3200 27062
rect 3148 26998 3200 27004
rect 2228 26988 2280 26994
rect 2228 26930 2280 26936
rect 1860 26920 1912 26926
rect 1860 26862 1912 26868
rect 1872 26382 1900 26862
rect 1860 26376 1912 26382
rect 1860 26318 1912 26324
rect 1952 26376 2004 26382
rect 1952 26318 2004 26324
rect 848 24812 900 24818
rect 848 24754 900 24760
rect 860 24721 888 24754
rect 846 24712 902 24721
rect 846 24647 902 24656
rect 848 24132 900 24138
rect 848 24074 900 24080
rect 860 24041 888 24074
rect 846 24032 902 24041
rect 846 23967 902 23976
rect 848 23112 900 23118
rect 846 23080 848 23089
rect 900 23080 902 23089
rect 846 23015 902 23024
rect 1398 22536 1454 22545
rect 1398 22471 1454 22480
rect 1412 22030 1440 22471
rect 1400 22024 1452 22030
rect 1400 21966 1452 21972
rect 1308 21616 1360 21622
rect 1308 21558 1360 21564
rect 1320 21185 1348 21558
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1306 21176 1362 21185
rect 1306 21111 1362 21120
rect 1412 20505 1440 21490
rect 1398 20496 1454 20505
rect 1398 20431 1454 20440
rect 846 19952 902 19961
rect 846 19887 902 19896
rect 860 19854 888 19887
rect 848 19848 900 19854
rect 848 19790 900 19796
rect 1584 19372 1636 19378
rect 1584 19314 1636 19320
rect 1872 19334 1900 26318
rect 1964 23662 1992 26318
rect 2136 24608 2188 24614
rect 2136 24550 2188 24556
rect 2148 24138 2176 24550
rect 2136 24132 2188 24138
rect 2136 24074 2188 24080
rect 2240 24070 2268 26930
rect 2320 26920 2372 26926
rect 2320 26862 2372 26868
rect 2332 26586 2360 26862
rect 2872 26784 2924 26790
rect 2872 26726 2924 26732
rect 2320 26580 2372 26586
rect 2320 26522 2372 26528
rect 2780 26308 2832 26314
rect 2884 26296 2912 26726
rect 3160 26586 3188 26998
rect 3712 26994 3740 27338
rect 3700 26988 3752 26994
rect 3700 26930 3752 26936
rect 3712 26586 3740 26930
rect 3896 26790 3924 27406
rect 3988 27130 4016 27406
rect 4068 27328 4120 27334
rect 4068 27270 4120 27276
rect 4712 27328 4764 27334
rect 4712 27270 4764 27276
rect 3976 27124 4028 27130
rect 3976 27066 4028 27072
rect 3884 26784 3936 26790
rect 3884 26726 3936 26732
rect 3148 26580 3200 26586
rect 3148 26522 3200 26528
rect 3700 26580 3752 26586
rect 3700 26522 3752 26528
rect 3056 26376 3108 26382
rect 3056 26318 3108 26324
rect 2832 26268 2912 26296
rect 2780 26250 2832 26256
rect 2792 25906 2820 26250
rect 2780 25900 2832 25906
rect 2780 25842 2832 25848
rect 2872 25832 2924 25838
rect 2872 25774 2924 25780
rect 2884 24886 2912 25774
rect 2872 24880 2924 24886
rect 2700 24818 2820 24834
rect 2872 24822 2924 24828
rect 2504 24812 2556 24818
rect 2504 24754 2556 24760
rect 2688 24812 2820 24818
rect 2740 24806 2820 24812
rect 2688 24754 2740 24760
rect 2516 24206 2544 24754
rect 2792 24410 2820 24806
rect 2964 24608 3016 24614
rect 2964 24550 3016 24556
rect 2780 24404 2832 24410
rect 2780 24346 2832 24352
rect 2976 24274 3004 24550
rect 2964 24268 3016 24274
rect 2964 24210 3016 24216
rect 2504 24200 2556 24206
rect 2504 24142 2556 24148
rect 2596 24200 2648 24206
rect 2596 24142 2648 24148
rect 2228 24064 2280 24070
rect 2228 24006 2280 24012
rect 1952 23656 2004 23662
rect 1952 23598 2004 23604
rect 2136 23044 2188 23050
rect 2136 22986 2188 22992
rect 2148 22574 2176 22986
rect 2136 22568 2188 22574
rect 2136 22510 2188 22516
rect 2148 21962 2176 22510
rect 2136 21956 2188 21962
rect 2136 21898 2188 21904
rect 2044 20800 2096 20806
rect 2044 20742 2096 20748
rect 2056 20466 2084 20742
rect 2240 20466 2268 24006
rect 2516 23798 2544 24142
rect 2504 23792 2556 23798
rect 2504 23734 2556 23740
rect 2608 23730 2636 24142
rect 2596 23724 2648 23730
rect 2596 23666 2648 23672
rect 2320 22976 2372 22982
rect 2320 22918 2372 22924
rect 2332 22642 2360 22918
rect 2320 22636 2372 22642
rect 2320 22578 2372 22584
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 2332 21554 2360 22034
rect 2608 22012 2636 23666
rect 2780 23588 2832 23594
rect 2780 23530 2832 23536
rect 2688 23180 2740 23186
rect 2688 23122 2740 23128
rect 2700 22982 2728 23122
rect 2688 22976 2740 22982
rect 2688 22918 2740 22924
rect 2792 22216 2820 23530
rect 2964 22976 3016 22982
rect 2964 22918 3016 22924
rect 2872 22772 2924 22778
rect 2872 22714 2924 22720
rect 2884 22409 2912 22714
rect 2976 22574 3004 22918
rect 2964 22568 3016 22574
rect 2964 22510 3016 22516
rect 2870 22400 2926 22409
rect 2870 22335 2926 22344
rect 2792 22188 3004 22216
rect 2778 22128 2834 22137
rect 2778 22063 2834 22072
rect 2688 22024 2740 22030
rect 2516 21984 2688 22012
rect 2320 21548 2372 21554
rect 2320 21490 2372 21496
rect 2332 21010 2360 21490
rect 2320 21004 2372 21010
rect 2320 20946 2372 20952
rect 2044 20460 2096 20466
rect 2044 20402 2096 20408
rect 2228 20460 2280 20466
rect 2228 20402 2280 20408
rect 2056 19922 2084 20402
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 2240 19854 2268 20402
rect 2228 19848 2280 19854
rect 2228 19790 2280 19796
rect 2320 19712 2372 19718
rect 2320 19654 2372 19660
rect 1492 18284 1544 18290
rect 1492 18226 1544 18232
rect 1504 17785 1532 18226
rect 1596 18086 1624 19314
rect 1872 19306 1992 19334
rect 1964 18358 1992 19306
rect 2332 18358 2360 19654
rect 1952 18352 2004 18358
rect 1872 18312 1952 18340
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1490 17776 1546 17785
rect 1490 17711 1546 17720
rect 1596 17678 1624 18022
rect 1584 17672 1636 17678
rect 1584 17614 1636 17620
rect 1872 17202 1900 18312
rect 1952 18294 2004 18300
rect 2320 18352 2372 18358
rect 2320 18294 2372 18300
rect 1952 17740 2004 17746
rect 1952 17682 2004 17688
rect 2412 17740 2464 17746
rect 2412 17682 2464 17688
rect 1860 17196 1912 17202
rect 1860 17138 1912 17144
rect 1964 17134 1992 17682
rect 2424 17338 2452 17682
rect 2412 17332 2464 17338
rect 2412 17274 2464 17280
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 848 16108 900 16114
rect 848 16050 900 16056
rect 860 15881 888 16050
rect 1860 16040 1912 16046
rect 1860 15982 1912 15988
rect 846 15872 902 15881
rect 846 15807 902 15816
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13705 1440 13874
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 1872 13326 1900 15982
rect 2412 15020 2464 15026
rect 2412 14962 2464 14968
rect 2424 14414 2452 14962
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 1964 13394 1992 13806
rect 2424 13530 2452 14350
rect 2412 13524 2464 13530
rect 2412 13466 2464 13472
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 2228 13388 2280 13394
rect 2228 13330 2280 13336
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 846 11792 902 11801
rect 846 11727 848 11736
rect 900 11727 902 11736
rect 848 11698 900 11704
rect 1964 10742 1992 13330
rect 2240 12782 2268 13330
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 2240 11830 2268 12582
rect 2516 12434 2544 21984
rect 2688 21966 2740 21972
rect 2596 20936 2648 20942
rect 2596 20878 2648 20884
rect 2608 19990 2636 20878
rect 2792 20466 2820 22063
rect 2872 22024 2924 22030
rect 2872 21966 2924 21972
rect 2884 21865 2912 21966
rect 2870 21856 2926 21865
rect 2870 21791 2926 21800
rect 2976 21622 3004 22188
rect 3068 21894 3096 26318
rect 3160 25906 3188 26522
rect 3896 26382 3924 26726
rect 3988 26586 4016 27066
rect 4080 26994 4108 27270
rect 4068 26988 4120 26994
rect 4068 26930 4120 26936
rect 4620 26988 4672 26994
rect 4620 26930 4672 26936
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 3976 26580 4028 26586
rect 3976 26522 4028 26528
rect 3884 26376 3936 26382
rect 3884 26318 3936 26324
rect 4632 26314 4660 26930
rect 4724 26518 4752 27270
rect 4816 26858 4844 27406
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 5276 27130 5304 27474
rect 5264 27124 5316 27130
rect 5264 27066 5316 27072
rect 5460 27010 5488 27542
rect 6184 27464 6236 27470
rect 6184 27406 6236 27412
rect 6000 27396 6052 27402
rect 6000 27338 6052 27344
rect 5540 27328 5592 27334
rect 5540 27270 5592 27276
rect 5816 27328 5868 27334
rect 5816 27270 5868 27276
rect 5092 26982 5488 27010
rect 4804 26852 4856 26858
rect 4804 26794 4856 26800
rect 4816 26586 4844 26794
rect 4804 26580 4856 26586
rect 4804 26522 4856 26528
rect 4712 26512 4764 26518
rect 4712 26454 4764 26460
rect 5092 26450 5120 26982
rect 5264 26920 5316 26926
rect 5264 26862 5316 26868
rect 5172 26580 5224 26586
rect 5172 26522 5224 26528
rect 5080 26444 5132 26450
rect 5080 26386 5132 26392
rect 5184 26382 5212 26522
rect 5172 26376 5224 26382
rect 5172 26318 5224 26324
rect 3424 26308 3476 26314
rect 3424 26250 3476 26256
rect 4620 26308 4672 26314
rect 4620 26250 4672 26256
rect 3148 25900 3200 25906
rect 3148 25842 3200 25848
rect 3436 24410 3464 26250
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4896 24880 4948 24886
rect 4896 24822 4948 24828
rect 4068 24812 4120 24818
rect 4068 24754 4120 24760
rect 3424 24404 3476 24410
rect 3424 24346 3476 24352
rect 4080 24342 4108 24754
rect 4712 24744 4764 24750
rect 4712 24686 4764 24692
rect 4620 24608 4672 24614
rect 4620 24550 4672 24556
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4068 24336 4120 24342
rect 4068 24278 4120 24284
rect 4436 24132 4488 24138
rect 4436 24074 4488 24080
rect 3148 24064 3200 24070
rect 3148 24006 3200 24012
rect 3160 23118 3188 24006
rect 4448 23610 4476 24074
rect 4632 23798 4660 24550
rect 4724 24206 4752 24686
rect 4804 24268 4856 24274
rect 4804 24210 4856 24216
rect 4712 24200 4764 24206
rect 4712 24142 4764 24148
rect 4620 23792 4672 23798
rect 4620 23734 4672 23740
rect 4724 23730 4752 24142
rect 4816 23866 4844 24210
rect 4908 24138 4936 24822
rect 5276 24818 5304 26862
rect 5368 24818 5396 26982
rect 5552 26382 5580 27270
rect 5724 27124 5776 27130
rect 5724 27066 5776 27072
rect 5632 27056 5684 27062
rect 5632 26998 5684 27004
rect 5644 26772 5672 26998
rect 5736 26926 5764 27066
rect 5828 27062 5856 27270
rect 5816 27056 5868 27062
rect 5816 26998 5868 27004
rect 5724 26920 5776 26926
rect 5724 26862 5776 26868
rect 5724 26784 5776 26790
rect 5644 26744 5724 26772
rect 5724 26726 5776 26732
rect 5828 26382 5856 26998
rect 6012 26994 6040 27338
rect 6092 27328 6144 27334
rect 6092 27270 6144 27276
rect 6000 26988 6052 26994
rect 6000 26930 6052 26936
rect 6104 26926 6132 27270
rect 6092 26920 6144 26926
rect 6092 26862 6144 26868
rect 6000 26784 6052 26790
rect 6000 26726 6052 26732
rect 5540 26376 5592 26382
rect 5540 26318 5592 26324
rect 5816 26376 5868 26382
rect 5816 26318 5868 26324
rect 5448 25968 5500 25974
rect 5448 25910 5500 25916
rect 5460 24818 5488 25910
rect 6012 25906 6040 26726
rect 6196 26586 6224 27406
rect 6380 26926 6408 27610
rect 6472 27470 6500 27814
rect 6932 27606 6960 28018
rect 9404 28008 9456 28014
rect 9404 27950 9456 27956
rect 7012 27872 7064 27878
rect 7012 27814 7064 27820
rect 6920 27600 6972 27606
rect 6920 27542 6972 27548
rect 6460 27464 6512 27470
rect 6460 27406 6512 27412
rect 6552 27464 6604 27470
rect 6552 27406 6604 27412
rect 6460 27328 6512 27334
rect 6460 27270 6512 27276
rect 6368 26920 6420 26926
rect 6368 26862 6420 26868
rect 6184 26580 6236 26586
rect 6184 26522 6236 26528
rect 6092 26308 6144 26314
rect 6092 26250 6144 26256
rect 6000 25900 6052 25906
rect 6000 25842 6052 25848
rect 5080 24812 5132 24818
rect 5080 24754 5132 24760
rect 5264 24812 5316 24818
rect 5264 24754 5316 24760
rect 5356 24812 5408 24818
rect 5356 24754 5408 24760
rect 5448 24812 5500 24818
rect 5448 24754 5500 24760
rect 5092 24274 5120 24754
rect 5080 24268 5132 24274
rect 5080 24210 5132 24216
rect 5276 24206 5304 24754
rect 5908 24676 5960 24682
rect 5908 24618 5960 24624
rect 5264 24200 5316 24206
rect 5264 24142 5316 24148
rect 4896 24132 4948 24138
rect 4896 24074 4948 24080
rect 5632 24132 5684 24138
rect 5632 24074 5684 24080
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4804 23860 4856 23866
rect 4804 23802 4856 23808
rect 5644 23798 5672 24074
rect 5632 23792 5684 23798
rect 5632 23734 5684 23740
rect 4712 23724 4764 23730
rect 4712 23666 4764 23672
rect 5264 23656 5316 23662
rect 4448 23582 4660 23610
rect 5264 23598 5316 23604
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23186 4660 23582
rect 4620 23180 4672 23186
rect 4620 23122 4672 23128
rect 3148 23112 3200 23118
rect 3148 23054 3200 23060
rect 3160 22642 3188 23054
rect 4252 23044 4304 23050
rect 4252 22986 4304 22992
rect 4620 23044 4672 23050
rect 4620 22986 4672 22992
rect 3792 22976 3844 22982
rect 3792 22918 3844 22924
rect 3804 22710 3832 22918
rect 4068 22772 4120 22778
rect 4068 22714 4120 22720
rect 3792 22704 3844 22710
rect 3792 22646 3844 22652
rect 3148 22636 3200 22642
rect 3148 22578 3200 22584
rect 3608 22568 3660 22574
rect 3608 22510 3660 22516
rect 3056 21888 3108 21894
rect 3056 21830 3108 21836
rect 2964 21616 3016 21622
rect 2964 21558 3016 21564
rect 2780 20460 2832 20466
rect 2780 20402 2832 20408
rect 2596 19984 2648 19990
rect 2596 19926 2648 19932
rect 2608 19378 2636 19926
rect 2688 19916 2740 19922
rect 2976 19904 3004 21558
rect 3620 21554 3648 22510
rect 3884 22432 3936 22438
rect 3884 22374 3936 22380
rect 3896 21894 3924 22374
rect 4080 22166 4108 22714
rect 4264 22710 4292 22986
rect 4252 22704 4304 22710
rect 4252 22646 4304 22652
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4068 22160 4120 22166
rect 4068 22102 4120 22108
rect 4080 22030 4108 22102
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 3884 21888 3936 21894
rect 3884 21830 3936 21836
rect 3976 21888 4028 21894
rect 3976 21830 4028 21836
rect 3988 21554 4016 21830
rect 3608 21548 3660 21554
rect 3608 21490 3660 21496
rect 3976 21548 4028 21554
rect 3976 21490 4028 21496
rect 3424 20392 3476 20398
rect 3424 20334 3476 20340
rect 3148 20256 3200 20262
rect 3148 20198 3200 20204
rect 3160 19922 3188 20198
rect 3436 19922 3464 20334
rect 3148 19916 3200 19922
rect 2976 19876 3096 19904
rect 2688 19858 2740 19864
rect 2596 19372 2648 19378
rect 2596 19314 2648 19320
rect 2700 18340 2728 19858
rect 2964 19780 3016 19786
rect 2964 19722 3016 19728
rect 2976 19378 3004 19722
rect 2964 19372 3016 19378
rect 2964 19314 3016 19320
rect 2608 18312 2728 18340
rect 2608 17678 2636 18312
rect 2872 18284 2924 18290
rect 2872 18226 2924 18232
rect 2884 17728 2912 18226
rect 2964 18216 3016 18222
rect 2964 18158 3016 18164
rect 2976 17882 3004 18158
rect 2964 17876 3016 17882
rect 2964 17818 3016 17824
rect 2884 17700 3004 17728
rect 2596 17672 2648 17678
rect 2596 17614 2648 17620
rect 2976 17610 3004 17700
rect 2964 17604 3016 17610
rect 2964 17546 3016 17552
rect 2688 17060 2740 17066
rect 2688 17002 2740 17008
rect 2700 15026 2728 17002
rect 2976 16658 3004 17546
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 2884 16250 2912 16526
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 2700 14482 2728 14962
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 2780 14544 2832 14550
rect 2780 14486 2832 14492
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 2792 13870 2820 14486
rect 2884 14482 2912 14758
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 3068 13920 3096 19876
rect 3148 19858 3200 19864
rect 3424 19916 3476 19922
rect 3424 19858 3476 19864
rect 3436 19310 3464 19858
rect 4080 19446 4108 21966
rect 4632 21894 4660 22986
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 4804 22500 4856 22506
rect 4804 22442 4856 22448
rect 4816 22030 4844 22442
rect 5276 22030 5304 23598
rect 5540 23588 5592 23594
rect 5540 23530 5592 23536
rect 5552 23186 5580 23530
rect 5540 23180 5592 23186
rect 5540 23122 5592 23128
rect 5644 23118 5672 23734
rect 5920 23730 5948 24618
rect 5908 23724 5960 23730
rect 5908 23666 5960 23672
rect 6104 23118 6132 26250
rect 5632 23112 5684 23118
rect 5632 23054 5684 23060
rect 6092 23112 6144 23118
rect 6092 23054 6144 23060
rect 6276 23044 6328 23050
rect 6276 22986 6328 22992
rect 4804 22024 4856 22030
rect 4804 21966 4856 21972
rect 5264 22024 5316 22030
rect 5264 21966 5316 21972
rect 4620 21888 4672 21894
rect 4620 21830 4672 21836
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4632 20942 4660 21830
rect 4816 21554 4844 21966
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 5276 21554 5304 21966
rect 6092 21956 6144 21962
rect 6092 21898 6144 21904
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 5264 21548 5316 21554
rect 5264 21490 5316 21496
rect 6104 21486 6132 21898
rect 4712 21480 4764 21486
rect 4712 21422 4764 21428
rect 5724 21480 5776 21486
rect 5724 21422 5776 21428
rect 6092 21480 6144 21486
rect 6092 21422 6144 21428
rect 4620 20936 4672 20942
rect 4620 20878 4672 20884
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4724 19854 4752 21422
rect 5736 20942 5764 21422
rect 6104 20942 6132 21422
rect 5264 20936 5316 20942
rect 5264 20878 5316 20884
rect 5724 20936 5776 20942
rect 5724 20878 5776 20884
rect 6092 20936 6144 20942
rect 6092 20878 6144 20884
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 4528 19780 4580 19786
rect 4528 19722 4580 19728
rect 4540 19446 4568 19722
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 5276 19446 5304 20878
rect 6288 20806 6316 22986
rect 6380 22982 6408 26862
rect 6472 26450 6500 27270
rect 6564 26994 6592 27406
rect 6932 27130 6960 27542
rect 6920 27124 6972 27130
rect 6920 27066 6972 27072
rect 6552 26988 6604 26994
rect 6552 26930 6604 26936
rect 6736 26988 6788 26994
rect 6736 26930 6788 26936
rect 6564 26858 6592 26930
rect 6552 26852 6604 26858
rect 6552 26794 6604 26800
rect 6564 26450 6592 26794
rect 6460 26444 6512 26450
rect 6460 26386 6512 26392
rect 6552 26444 6604 26450
rect 6552 26386 6604 26392
rect 6748 26382 6776 26930
rect 7024 26926 7052 27814
rect 9416 27470 9444 27950
rect 10152 27606 10180 28086
rect 10968 28076 11020 28082
rect 10968 28018 11020 28024
rect 11796 28076 11848 28082
rect 11796 28018 11848 28024
rect 12256 28076 12308 28082
rect 12256 28018 12308 28024
rect 10232 27872 10284 27878
rect 10232 27814 10284 27820
rect 10876 27872 10928 27878
rect 10876 27814 10928 27820
rect 10140 27600 10192 27606
rect 10140 27542 10192 27548
rect 10244 27470 10272 27814
rect 10888 27674 10916 27814
rect 10876 27668 10928 27674
rect 10876 27610 10928 27616
rect 10324 27600 10376 27606
rect 10322 27568 10324 27577
rect 10376 27568 10378 27577
rect 10322 27503 10378 27512
rect 10782 27568 10838 27577
rect 10782 27503 10784 27512
rect 10836 27503 10838 27512
rect 10784 27474 10836 27480
rect 7932 27464 7984 27470
rect 7932 27406 7984 27412
rect 9404 27464 9456 27470
rect 9404 27406 9456 27412
rect 10232 27464 10284 27470
rect 10232 27406 10284 27412
rect 7380 27328 7432 27334
rect 7380 27270 7432 27276
rect 7392 26994 7420 27270
rect 7944 26994 7972 27406
rect 9496 27396 9548 27402
rect 9496 27338 9548 27344
rect 8300 27328 8352 27334
rect 8300 27270 8352 27276
rect 9312 27328 9364 27334
rect 9312 27270 9364 27276
rect 8312 27062 8340 27270
rect 8300 27056 8352 27062
rect 8300 26998 8352 27004
rect 7380 26988 7432 26994
rect 7380 26930 7432 26936
rect 7932 26988 7984 26994
rect 7932 26930 7984 26936
rect 9128 26988 9180 26994
rect 9128 26930 9180 26936
rect 7012 26920 7064 26926
rect 7012 26862 7064 26868
rect 6920 26784 6972 26790
rect 6920 26726 6972 26732
rect 8208 26784 8260 26790
rect 8208 26726 8260 26732
rect 6932 26586 6960 26726
rect 6920 26580 6972 26586
rect 6920 26522 6972 26528
rect 6736 26376 6788 26382
rect 6736 26318 6788 26324
rect 6828 26240 6880 26246
rect 6828 26182 6880 26188
rect 6840 25838 6868 26182
rect 8220 25974 8248 26726
rect 9140 26382 9168 26930
rect 9324 26382 9352 27270
rect 9128 26376 9180 26382
rect 9128 26318 9180 26324
rect 9312 26376 9364 26382
rect 9312 26318 9364 26324
rect 8852 26240 8904 26246
rect 8852 26182 8904 26188
rect 8208 25968 8260 25974
rect 8208 25910 8260 25916
rect 8864 25906 8892 26182
rect 8852 25900 8904 25906
rect 8852 25842 8904 25848
rect 6828 25832 6880 25838
rect 6828 25774 6880 25780
rect 7564 25696 7616 25702
rect 7564 25638 7616 25644
rect 7656 25696 7708 25702
rect 7656 25638 7708 25644
rect 8668 25696 8720 25702
rect 8668 25638 8720 25644
rect 7576 24206 7604 25638
rect 7668 24818 7696 25638
rect 8680 24818 8708 25638
rect 7656 24812 7708 24818
rect 7656 24754 7708 24760
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 8668 24812 8720 24818
rect 8668 24754 8720 24760
rect 8404 24682 8432 24754
rect 8392 24676 8444 24682
rect 8392 24618 8444 24624
rect 8404 24410 8432 24618
rect 9312 24608 9364 24614
rect 9312 24550 9364 24556
rect 9404 24608 9456 24614
rect 9404 24550 9456 24556
rect 8392 24404 8444 24410
rect 8392 24346 8444 24352
rect 7472 24200 7524 24206
rect 7472 24142 7524 24148
rect 7564 24200 7616 24206
rect 7564 24142 7616 24148
rect 7484 23730 7512 24142
rect 7472 23724 7524 23730
rect 7472 23666 7524 23672
rect 7576 23662 7604 24142
rect 9220 24132 9272 24138
rect 9220 24074 9272 24080
rect 9232 23866 9260 24074
rect 9220 23860 9272 23866
rect 9220 23802 9272 23808
rect 9324 23730 9352 24550
rect 9416 24206 9444 24550
rect 9404 24200 9456 24206
rect 9404 24142 9456 24148
rect 9416 23798 9444 24142
rect 9404 23792 9456 23798
rect 9404 23734 9456 23740
rect 9036 23724 9088 23730
rect 9036 23666 9088 23672
rect 9312 23724 9364 23730
rect 9312 23666 9364 23672
rect 7564 23656 7616 23662
rect 7564 23598 7616 23604
rect 6920 23588 6972 23594
rect 6920 23530 6972 23536
rect 8116 23588 8168 23594
rect 8116 23530 8168 23536
rect 6932 23118 6960 23530
rect 7840 23316 7892 23322
rect 7840 23258 7892 23264
rect 6920 23112 6972 23118
rect 6920 23054 6972 23060
rect 6736 23044 6788 23050
rect 6736 22986 6788 22992
rect 6368 22976 6420 22982
rect 6368 22918 6420 22924
rect 6748 22642 6776 22986
rect 6932 22642 6960 23054
rect 7656 23044 7708 23050
rect 7656 22986 7708 22992
rect 7668 22642 7696 22986
rect 7852 22642 7880 23258
rect 8128 22982 8156 23530
rect 9048 23118 9076 23666
rect 9312 23180 9364 23186
rect 9312 23122 9364 23128
rect 9036 23112 9088 23118
rect 9036 23054 9088 23060
rect 8392 23044 8444 23050
rect 8392 22986 8444 22992
rect 8116 22976 8168 22982
rect 8116 22918 8168 22924
rect 8128 22710 8156 22918
rect 8404 22778 8432 22986
rect 8852 22976 8904 22982
rect 8852 22918 8904 22924
rect 8392 22772 8444 22778
rect 8392 22714 8444 22720
rect 8864 22710 8892 22918
rect 8116 22704 8168 22710
rect 8116 22646 8168 22652
rect 8852 22704 8904 22710
rect 8852 22646 8904 22652
rect 9048 22642 9076 23054
rect 9324 22642 9352 23122
rect 6736 22636 6788 22642
rect 6736 22578 6788 22584
rect 6920 22636 6972 22642
rect 6920 22578 6972 22584
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7656 22636 7708 22642
rect 7656 22578 7708 22584
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 9036 22636 9088 22642
rect 9036 22578 9088 22584
rect 9312 22636 9364 22642
rect 9312 22578 9364 22584
rect 7484 21622 7512 22578
rect 7472 21616 7524 21622
rect 7472 21558 7524 21564
rect 7668 21554 7696 22578
rect 9324 22030 9352 22578
rect 9312 22024 9364 22030
rect 9312 21966 9364 21972
rect 7656 21548 7708 21554
rect 7656 21490 7708 21496
rect 8576 21412 8628 21418
rect 8576 21354 8628 21360
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 6932 20924 6960 21286
rect 7104 20936 7156 20942
rect 6932 20896 7104 20924
rect 6552 20868 6604 20874
rect 6552 20810 6604 20816
rect 6276 20800 6328 20806
rect 6276 20742 6328 20748
rect 6288 20466 6316 20742
rect 6276 20460 6328 20466
rect 6276 20402 6328 20408
rect 6368 19848 6420 19854
rect 6368 19790 6420 19796
rect 5356 19712 5408 19718
rect 5356 19654 5408 19660
rect 6000 19712 6052 19718
rect 6000 19654 6052 19660
rect 4068 19440 4120 19446
rect 4068 19382 4120 19388
rect 4528 19440 4580 19446
rect 4528 19382 4580 19388
rect 5264 19440 5316 19446
rect 5264 19382 5316 19388
rect 3424 19304 3476 19310
rect 3424 19246 3476 19252
rect 4068 19304 4120 19310
rect 4068 19246 4120 19252
rect 4712 19304 4764 19310
rect 4712 19246 4764 19252
rect 3148 18216 3200 18222
rect 3148 18158 3200 18164
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 3160 17814 3188 18158
rect 3424 18080 3476 18086
rect 3424 18022 3476 18028
rect 3148 17808 3200 17814
rect 3148 17750 3200 17756
rect 3160 16114 3188 17750
rect 3436 17202 3464 18022
rect 3424 17196 3476 17202
rect 3424 17138 3476 17144
rect 3516 16652 3568 16658
rect 3516 16594 3568 16600
rect 3148 16108 3200 16114
rect 3148 16050 3200 16056
rect 3528 15026 3556 16594
rect 3896 16114 3924 18158
rect 4080 17338 4108 19246
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4724 18222 4752 19246
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4816 18426 4844 18702
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 5276 18290 5304 19382
rect 5368 19378 5396 19654
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5356 19372 5408 19378
rect 5356 19314 5408 19320
rect 5368 18766 5396 19314
rect 5356 18760 5408 18766
rect 5356 18702 5408 18708
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 4080 17202 4108 17274
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 4620 17060 4672 17066
rect 4620 17002 4672 17008
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16114 4660 17002
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4724 16114 4752 16934
rect 4804 16516 4856 16522
rect 4804 16458 4856 16464
rect 3884 16108 3936 16114
rect 3884 16050 3936 16056
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4816 16046 4844 16458
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 4804 16040 4856 16046
rect 4804 15982 4856 15988
rect 3792 15904 3844 15910
rect 3792 15846 3844 15852
rect 3804 15502 3832 15846
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3344 14618 3372 14962
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3792 14612 3844 14618
rect 3792 14554 3844 14560
rect 3332 14408 3384 14414
rect 3332 14350 3384 14356
rect 3148 14340 3200 14346
rect 3148 14282 3200 14288
rect 3160 13938 3188 14282
rect 3344 14074 3372 14350
rect 3608 14340 3660 14346
rect 3608 14282 3660 14288
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3620 14006 3648 14282
rect 3804 14074 3832 14554
rect 3896 14414 3924 14758
rect 3988 14550 4016 15982
rect 4620 15904 4672 15910
rect 5460 15858 5488 19450
rect 6012 19378 6040 19654
rect 6000 19372 6052 19378
rect 6000 19314 6052 19320
rect 6092 19168 6144 19174
rect 6092 19110 6144 19116
rect 6104 18766 6132 19110
rect 6092 18760 6144 18766
rect 6092 18702 6144 18708
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5736 16590 5764 18566
rect 6380 18290 6408 19790
rect 6564 19378 6592 20810
rect 6932 20466 6960 20896
rect 7104 20878 7156 20884
rect 8300 20868 8352 20874
rect 8300 20810 8352 20816
rect 8312 20466 8340 20810
rect 6920 20460 6972 20466
rect 6920 20402 6972 20408
rect 7932 20460 7984 20466
rect 7932 20402 7984 20408
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 7944 19854 7972 20402
rect 8312 19922 8340 20402
rect 8392 20324 8444 20330
rect 8392 20266 8444 20272
rect 8300 19916 8352 19922
rect 8300 19858 8352 19864
rect 7932 19848 7984 19854
rect 7932 19790 7984 19796
rect 8404 19514 8432 20266
rect 8392 19508 8444 19514
rect 8392 19450 8444 19456
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 8208 19372 8260 19378
rect 8208 19314 8260 19320
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 6472 18358 6500 19110
rect 6564 18766 6592 19314
rect 8220 18970 8248 19314
rect 8404 19258 8432 19450
rect 8588 19378 8616 21354
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8312 19230 8432 19258
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 8312 18766 8340 19230
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 7656 18692 7708 18698
rect 7656 18634 7708 18640
rect 6460 18352 6512 18358
rect 6460 18294 6512 18300
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 5724 16584 5776 16590
rect 5724 16526 5776 16532
rect 5736 16114 5764 16526
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 4620 15846 4672 15852
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15570 4660 15846
rect 4816 15830 5488 15858
rect 5724 15904 5776 15910
rect 5724 15846 5776 15852
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 4724 15026 4752 15302
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 3976 14544 4028 14550
rect 3976 14486 4028 14492
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 4080 14260 4108 14894
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4724 14550 4752 14962
rect 4712 14544 4764 14550
rect 4712 14486 4764 14492
rect 4160 14272 4212 14278
rect 4080 14232 4160 14260
rect 4160 14214 4212 14220
rect 3792 14068 3844 14074
rect 3792 14010 3844 14016
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 3608 14000 3660 14006
rect 3608 13942 3660 13948
rect 4080 13938 4108 14010
rect 4172 13938 4200 14214
rect 2976 13892 3096 13920
rect 3148 13932 3200 13938
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2976 13326 3004 13892
rect 3148 13874 3200 13880
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 3056 13796 3108 13802
rect 3056 13738 3108 13744
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 2976 12850 3004 13262
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2516 12406 2636 12434
rect 2228 11824 2280 11830
rect 2228 11766 2280 11772
rect 2240 11218 2268 11766
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2228 11212 2280 11218
rect 2228 11154 2280 11160
rect 2332 11150 2360 11698
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2332 10810 2360 11086
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 1952 10736 2004 10742
rect 1952 10678 2004 10684
rect 2608 10674 2636 12406
rect 3068 12306 3096 13738
rect 3240 12368 3292 12374
rect 3240 12310 3292 12316
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 3252 12238 3280 12310
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3252 11898 3280 12174
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 4080 11762 4108 13874
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4816 12434 4844 15830
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 5736 15026 5764 15846
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5724 15020 5776 15026
rect 5724 14962 5776 14968
rect 5276 14482 5304 14962
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6840 14482 6868 14894
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 6748 13938 6776 14350
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 5552 12850 5580 13806
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 4632 12406 4844 12434
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 4540 11694 4568 12038
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 2792 10810 2820 11562
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2148 10130 2176 10406
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 2608 10062 2636 10610
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2700 8974 2728 10746
rect 2976 10606 3004 11290
rect 3344 10674 3372 11630
rect 3528 11354 3556 11630
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 3976 10532 4028 10538
rect 3976 10474 4028 10480
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2976 8430 3004 9862
rect 3988 9518 4016 10474
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 3884 9036 3936 9042
rect 3884 8978 3936 8984
rect 3896 8498 3924 8978
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3988 8634 4016 8910
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 4632 8566 4660 12406
rect 5368 12306 5396 12718
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 5552 12238 5580 12786
rect 6196 12238 6224 12786
rect 6656 12238 6684 12786
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 4724 11762 4752 12174
rect 4816 11830 4844 12174
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 5092 10996 5120 11698
rect 5540 11620 5592 11626
rect 5540 11562 5592 11568
rect 5092 10968 5304 10996
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5276 9586 5304 10968
rect 5552 10606 5580 11562
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6564 10810 6592 11018
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5644 9722 5672 10610
rect 5632 9716 5684 9722
rect 5632 9658 5684 9664
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 4724 9178 4752 9522
rect 5172 9444 5224 9450
rect 5172 9386 5224 9392
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 5184 9042 5212 9386
rect 5276 9110 5304 9522
rect 6656 9518 6684 12174
rect 6748 11558 6776 13874
rect 6840 13870 6868 14418
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6840 13326 6868 13670
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6748 11286 6776 11494
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 3896 7954 3924 8434
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7970 4660 8502
rect 4724 8294 4752 8910
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5276 8566 5304 9046
rect 5368 8906 5396 9386
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5264 8560 5316 8566
rect 5264 8502 5316 8508
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4540 7954 4660 7970
rect 4724 7954 4752 8230
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 4528 7948 4660 7954
rect 4580 7942 4660 7948
rect 4712 7948 4764 7954
rect 4528 7890 4580 7896
rect 4712 7890 4764 7896
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4356 7546 4384 7822
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 5276 7410 5304 8502
rect 5368 8498 5396 8842
rect 5460 8634 5488 8910
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 5460 6934 5488 7686
rect 5552 7342 5580 8774
rect 6932 8634 6960 8774
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5644 7342 5672 7958
rect 6932 7954 6960 8570
rect 7024 8498 7052 18022
rect 7576 17678 7604 18226
rect 7668 18222 7696 18634
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 7668 17678 7696 18158
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7576 17320 7604 17614
rect 8312 17338 8340 17682
rect 8300 17332 8352 17338
rect 7576 17292 7696 17320
rect 7564 17196 7616 17202
rect 7564 17138 7616 17144
rect 7380 16584 7432 16590
rect 7380 16526 7432 16532
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7196 16108 7248 16114
rect 7196 16050 7248 16056
rect 7208 14890 7236 16050
rect 7288 15972 7340 15978
rect 7288 15914 7340 15920
rect 7300 15502 7328 15914
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 7300 15162 7328 15438
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 7196 14884 7248 14890
rect 7196 14826 7248 14832
rect 7300 14550 7328 15098
rect 7392 15026 7420 16526
rect 7484 15026 7512 16526
rect 7576 16250 7604 17138
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7288 14544 7340 14550
rect 7288 14486 7340 14492
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7116 12986 7144 13262
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7484 12434 7512 13262
rect 7392 12406 7512 12434
rect 7392 12374 7420 12406
rect 7380 12368 7432 12374
rect 7380 12310 7432 12316
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7116 11762 7144 12174
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7116 11014 7144 11698
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7208 10606 7236 11154
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7392 10674 7420 11086
rect 7668 10742 7696 17292
rect 8300 17274 8352 17280
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7852 16114 7880 17138
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 8128 15910 8156 16594
rect 8312 16114 8340 17274
rect 8404 16726 8432 19110
rect 8588 18766 8616 19314
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8680 18426 8708 18770
rect 8772 18766 8800 19654
rect 8760 18760 8812 18766
rect 8760 18702 8812 18708
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 8668 18420 8720 18426
rect 8668 18362 8720 18368
rect 9232 18290 9260 18566
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 8852 17672 8904 17678
rect 8852 17614 8904 17620
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 8680 16794 8708 17138
rect 8864 17134 8892 17614
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8944 17128 8996 17134
rect 8944 17070 8996 17076
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8392 16720 8444 16726
rect 8392 16662 8444 16668
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8128 15502 8156 15846
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 8128 15094 8156 15438
rect 8116 15088 8168 15094
rect 8116 15030 8168 15036
rect 8588 14958 8616 16526
rect 8680 15026 8708 16730
rect 8956 16590 8984 17070
rect 9324 16658 9352 21966
rect 9508 19786 9536 27338
rect 10244 26926 10272 27406
rect 10980 27130 11008 28018
rect 11704 27872 11756 27878
rect 11704 27814 11756 27820
rect 11244 27668 11296 27674
rect 11244 27610 11296 27616
rect 10968 27124 11020 27130
rect 10968 27066 11020 27072
rect 11256 26994 11284 27610
rect 11716 27470 11744 27814
rect 11808 27674 11836 28018
rect 12072 28008 12124 28014
rect 12072 27950 12124 27956
rect 11796 27668 11848 27674
rect 11796 27610 11848 27616
rect 11794 27568 11850 27577
rect 11794 27503 11850 27512
rect 11808 27470 11836 27503
rect 11336 27464 11388 27470
rect 11336 27406 11388 27412
rect 11704 27464 11756 27470
rect 11704 27406 11756 27412
rect 11796 27464 11848 27470
rect 11796 27406 11848 27412
rect 11348 27062 11376 27406
rect 11336 27056 11388 27062
rect 11336 26998 11388 27004
rect 10600 26988 10652 26994
rect 10600 26930 10652 26936
rect 11244 26988 11296 26994
rect 11244 26930 11296 26936
rect 10232 26920 10284 26926
rect 10232 26862 10284 26868
rect 9864 26580 9916 26586
rect 9864 26522 9916 26528
rect 9772 26240 9824 26246
rect 9772 26182 9824 26188
rect 9784 25294 9812 26182
rect 9876 25294 9904 26522
rect 10612 26382 10640 26930
rect 10692 26784 10744 26790
rect 10692 26726 10744 26732
rect 10600 26376 10652 26382
rect 10600 26318 10652 26324
rect 10704 25294 10732 26726
rect 11256 26450 11284 26930
rect 11348 26858 11376 26998
rect 11716 26994 11744 27406
rect 11888 27328 11940 27334
rect 11888 27270 11940 27276
rect 11980 27328 12032 27334
rect 11980 27270 12032 27276
rect 11900 26994 11928 27270
rect 11704 26988 11756 26994
rect 11704 26930 11756 26936
rect 11888 26988 11940 26994
rect 11888 26930 11940 26936
rect 11336 26852 11388 26858
rect 11336 26794 11388 26800
rect 11244 26444 11296 26450
rect 11244 26386 11296 26392
rect 11348 26382 11376 26794
rect 11992 26790 12020 27270
rect 12084 27130 12112 27950
rect 12268 27470 12296 28018
rect 14660 27713 14688 28426
rect 14646 27704 14702 27713
rect 14646 27639 14702 27648
rect 12164 27464 12216 27470
rect 12164 27406 12216 27412
rect 12256 27464 12308 27470
rect 12256 27406 12308 27412
rect 12072 27124 12124 27130
rect 12072 27066 12124 27072
rect 11980 26784 12032 26790
rect 11980 26726 12032 26732
rect 11992 26382 12020 26726
rect 11336 26376 11388 26382
rect 11336 26318 11388 26324
rect 11980 26376 12032 26382
rect 11980 26318 12032 26324
rect 10876 26240 10928 26246
rect 10876 26182 10928 26188
rect 10888 25294 10916 26182
rect 12084 25786 12112 27066
rect 12176 26994 12204 27406
rect 12164 26988 12216 26994
rect 12164 26930 12216 26936
rect 12268 26790 12296 27406
rect 12808 27396 12860 27402
rect 12808 27338 12860 27344
rect 12532 27056 12584 27062
rect 12532 26998 12584 27004
rect 12440 26852 12492 26858
rect 12440 26794 12492 26800
rect 12256 26784 12308 26790
rect 12256 26726 12308 26732
rect 12268 26042 12296 26726
rect 12452 26246 12480 26794
rect 12544 26586 12572 26998
rect 12532 26580 12584 26586
rect 12532 26522 12584 26528
rect 12624 26512 12676 26518
rect 12624 26454 12676 26460
rect 12532 26376 12584 26382
rect 12532 26318 12584 26324
rect 12440 26240 12492 26246
rect 12440 26182 12492 26188
rect 12452 26042 12480 26182
rect 12256 26036 12308 26042
rect 12256 25978 12308 25984
rect 12440 26036 12492 26042
rect 12440 25978 12492 25984
rect 12084 25758 12204 25786
rect 12072 25696 12124 25702
rect 12072 25638 12124 25644
rect 9772 25288 9824 25294
rect 9772 25230 9824 25236
rect 9864 25288 9916 25294
rect 9864 25230 9916 25236
rect 10692 25288 10744 25294
rect 10692 25230 10744 25236
rect 10876 25288 10928 25294
rect 10876 25230 10928 25236
rect 9864 25152 9916 25158
rect 9864 25094 9916 25100
rect 10692 25152 10744 25158
rect 10692 25094 10744 25100
rect 9876 24886 9904 25094
rect 9864 24880 9916 24886
rect 9864 24822 9916 24828
rect 9876 24206 9904 24822
rect 10704 24818 10732 25094
rect 10888 24954 10916 25230
rect 11060 25220 11112 25226
rect 11060 25162 11112 25168
rect 10968 25152 11020 25158
rect 10968 25094 11020 25100
rect 10980 24954 11008 25094
rect 11072 24954 11100 25162
rect 11888 25152 11940 25158
rect 11888 25094 11940 25100
rect 10876 24948 10928 24954
rect 10876 24890 10928 24896
rect 10968 24948 11020 24954
rect 10968 24890 11020 24896
rect 11060 24948 11112 24954
rect 11060 24890 11112 24896
rect 10692 24812 10744 24818
rect 10692 24754 10744 24760
rect 10876 24812 10928 24818
rect 10876 24754 10928 24760
rect 10416 24608 10468 24614
rect 10416 24550 10468 24556
rect 9864 24200 9916 24206
rect 9864 24142 9916 24148
rect 9956 24200 10008 24206
rect 10140 24200 10192 24206
rect 10008 24160 10140 24188
rect 9956 24142 10008 24148
rect 10140 24142 10192 24148
rect 10232 23724 10284 23730
rect 10232 23666 10284 23672
rect 9864 23656 9916 23662
rect 9864 23598 9916 23604
rect 9876 23322 9904 23598
rect 9864 23316 9916 23322
rect 9864 23258 9916 23264
rect 9588 22976 9640 22982
rect 9588 22918 9640 22924
rect 9600 22778 9628 22918
rect 9588 22772 9640 22778
rect 9588 22714 9640 22720
rect 9600 22030 9628 22714
rect 10244 22642 10272 23666
rect 10428 23118 10456 24550
rect 10888 24342 10916 24754
rect 10980 24682 11008 24890
rect 10968 24676 11020 24682
rect 10968 24618 11020 24624
rect 11704 24608 11756 24614
rect 11704 24550 11756 24556
rect 10876 24336 10928 24342
rect 10876 24278 10928 24284
rect 11716 24274 11744 24550
rect 11704 24268 11756 24274
rect 11704 24210 11756 24216
rect 10876 24200 10928 24206
rect 10876 24142 10928 24148
rect 10600 24132 10652 24138
rect 10600 24074 10652 24080
rect 10508 23520 10560 23526
rect 10508 23462 10560 23468
rect 10520 23118 10548 23462
rect 10612 23118 10640 24074
rect 10888 23798 10916 24142
rect 10876 23792 10928 23798
rect 10876 23734 10928 23740
rect 10888 23118 10916 23734
rect 10416 23112 10468 23118
rect 10416 23054 10468 23060
rect 10508 23112 10560 23118
rect 10508 23054 10560 23060
rect 10600 23112 10652 23118
rect 10600 23054 10652 23060
rect 10876 23112 10928 23118
rect 10876 23054 10928 23060
rect 10612 22778 10640 23054
rect 11060 22976 11112 22982
rect 11060 22918 11112 22924
rect 10600 22772 10652 22778
rect 10600 22714 10652 22720
rect 11072 22710 11100 22918
rect 11060 22704 11112 22710
rect 11060 22646 11112 22652
rect 10232 22636 10284 22642
rect 10232 22578 10284 22584
rect 10244 22030 10272 22578
rect 11900 22030 11928 25094
rect 12084 24886 12112 25638
rect 12072 24880 12124 24886
rect 12072 24822 12124 24828
rect 11980 24744 12032 24750
rect 11980 24686 12032 24692
rect 11992 24206 12020 24686
rect 12084 24206 12112 24822
rect 11980 24200 12032 24206
rect 11980 24142 12032 24148
rect 12072 24200 12124 24206
rect 12072 24142 12124 24148
rect 11992 23322 12020 24142
rect 11980 23316 12032 23322
rect 11980 23258 12032 23264
rect 12176 23186 12204 25758
rect 12440 25492 12492 25498
rect 12440 25434 12492 25440
rect 12452 25294 12480 25434
rect 12440 25288 12492 25294
rect 12440 25230 12492 25236
rect 12440 25152 12492 25158
rect 12440 25094 12492 25100
rect 12348 24744 12400 24750
rect 12348 24686 12400 24692
rect 12360 23662 12388 24686
rect 12452 24070 12480 25094
rect 12544 24750 12572 26318
rect 12636 25838 12664 26454
rect 12716 26308 12768 26314
rect 12716 26250 12768 26256
rect 12728 25906 12756 26250
rect 12820 25974 12848 27338
rect 12992 27328 13044 27334
rect 12912 27288 12992 27316
rect 12808 25968 12860 25974
rect 12808 25910 12860 25916
rect 12716 25900 12768 25906
rect 12716 25842 12768 25848
rect 12624 25832 12676 25838
rect 12624 25774 12676 25780
rect 12808 25832 12860 25838
rect 12912 25820 12940 27288
rect 12992 27270 13044 27276
rect 16868 27130 16896 28426
rect 17144 27606 17172 28494
rect 17236 27674 17264 28630
rect 26056 28552 26108 28558
rect 26056 28494 26108 28500
rect 18144 28484 18196 28490
rect 18144 28426 18196 28432
rect 18420 28484 18472 28490
rect 18420 28426 18472 28432
rect 19340 28484 19392 28490
rect 19340 28426 19392 28432
rect 20076 28484 20128 28490
rect 20076 28426 20128 28432
rect 20444 28484 20496 28490
rect 20444 28426 20496 28432
rect 20996 28484 21048 28490
rect 20996 28426 21048 28432
rect 21456 28484 21508 28490
rect 21456 28426 21508 28432
rect 22468 28484 22520 28490
rect 22468 28426 22520 28432
rect 23020 28484 23072 28490
rect 23020 28426 23072 28432
rect 23112 28484 23164 28490
rect 23112 28426 23164 28432
rect 24492 28484 24544 28490
rect 24492 28426 24544 28432
rect 25044 28484 25096 28490
rect 25044 28426 25096 28432
rect 25596 28484 25648 28490
rect 25596 28426 25648 28432
rect 17776 28416 17828 28422
rect 17776 28358 17828 28364
rect 17592 28008 17644 28014
rect 17592 27950 17644 27956
rect 17224 27668 17276 27674
rect 17224 27610 17276 27616
rect 17132 27600 17184 27606
rect 17132 27542 17184 27548
rect 17604 27470 17632 27950
rect 17788 27606 17816 28358
rect 17960 28076 18012 28082
rect 17960 28018 18012 28024
rect 17776 27600 17828 27606
rect 17776 27542 17828 27548
rect 17592 27464 17644 27470
rect 17592 27406 17644 27412
rect 17868 27464 17920 27470
rect 17972 27452 18000 28018
rect 18156 27674 18184 28426
rect 18432 28218 18460 28426
rect 18420 28212 18472 28218
rect 18420 28154 18472 28160
rect 19156 28008 19208 28014
rect 19156 27950 19208 27956
rect 19064 27940 19116 27946
rect 19064 27882 19116 27888
rect 19076 27674 19104 27882
rect 18144 27668 18196 27674
rect 18144 27610 18196 27616
rect 19064 27668 19116 27674
rect 19064 27610 19116 27616
rect 17920 27424 18000 27452
rect 17868 27406 17920 27412
rect 16856 27124 16908 27130
rect 16856 27066 16908 27072
rect 13084 26784 13136 26790
rect 13084 26726 13136 26732
rect 13096 26382 13124 26726
rect 17972 26586 18000 27424
rect 18052 27464 18104 27470
rect 18052 27406 18104 27412
rect 18970 27432 19026 27441
rect 18064 26994 18092 27406
rect 18970 27367 19026 27376
rect 18236 27328 18288 27334
rect 18236 27270 18288 27276
rect 18248 26994 18276 27270
rect 18984 27062 19012 27367
rect 18972 27056 19024 27062
rect 18972 26998 19024 27004
rect 18052 26988 18104 26994
rect 18052 26930 18104 26936
rect 18236 26988 18288 26994
rect 18236 26930 18288 26936
rect 19076 26874 19104 27610
rect 19168 26994 19196 27950
rect 19352 27130 19380 28426
rect 19628 28206 19932 28234
rect 20088 28218 20116 28426
rect 20456 28218 20484 28426
rect 19628 28150 19656 28206
rect 19432 28144 19484 28150
rect 19432 28086 19484 28092
rect 19616 28144 19668 28150
rect 19616 28086 19668 28092
rect 19444 27946 19472 28086
rect 19708 28076 19760 28082
rect 19708 28018 19760 28024
rect 19800 28076 19852 28082
rect 19800 28018 19852 28024
rect 19720 27962 19748 28018
rect 19432 27940 19484 27946
rect 19432 27882 19484 27888
rect 19536 27934 19748 27962
rect 19432 27668 19484 27674
rect 19432 27610 19484 27616
rect 19444 27334 19472 27610
rect 19536 27538 19564 27934
rect 19616 27872 19668 27878
rect 19616 27814 19668 27820
rect 19524 27532 19576 27538
rect 19524 27474 19576 27480
rect 19536 27402 19564 27474
rect 19524 27396 19576 27402
rect 19524 27338 19576 27344
rect 19432 27328 19484 27334
rect 19536 27305 19564 27338
rect 19432 27270 19484 27276
rect 19522 27296 19578 27305
rect 19340 27124 19392 27130
rect 19340 27066 19392 27072
rect 19156 26988 19208 26994
rect 19156 26930 19208 26936
rect 19248 26988 19300 26994
rect 19248 26930 19300 26936
rect 19260 26874 19288 26930
rect 19340 26920 19392 26926
rect 19076 26846 19288 26874
rect 19338 26888 19340 26897
rect 19392 26888 19394 26897
rect 19338 26823 19394 26832
rect 19444 26790 19472 27270
rect 19522 27231 19578 27240
rect 19536 26994 19564 27231
rect 19628 27130 19656 27814
rect 19812 27538 19840 28018
rect 19904 27946 19932 28206
rect 19984 28212 20036 28218
rect 19984 28154 20036 28160
rect 20076 28212 20128 28218
rect 20076 28154 20128 28160
rect 20444 28212 20496 28218
rect 20444 28154 20496 28160
rect 19996 28014 20024 28154
rect 20904 28144 20956 28150
rect 20904 28086 20956 28092
rect 19984 28008 20036 28014
rect 19984 27950 20036 27956
rect 19892 27940 19944 27946
rect 19892 27882 19944 27888
rect 20628 27940 20680 27946
rect 20628 27882 20680 27888
rect 19904 27606 19932 27882
rect 19892 27600 19944 27606
rect 19984 27600 20036 27606
rect 19892 27542 19944 27548
rect 19982 27568 19984 27577
rect 20076 27600 20128 27606
rect 20036 27568 20038 27577
rect 19800 27532 19852 27538
rect 20076 27542 20128 27548
rect 19982 27503 20038 27512
rect 19800 27474 19852 27480
rect 20088 27402 20116 27542
rect 20168 27532 20220 27538
rect 20168 27474 20220 27480
rect 20180 27441 20208 27474
rect 20352 27464 20404 27470
rect 20166 27432 20222 27441
rect 19800 27396 19852 27402
rect 19800 27338 19852 27344
rect 20076 27396 20128 27402
rect 20352 27406 20404 27412
rect 20166 27367 20222 27376
rect 20076 27338 20128 27344
rect 19616 27124 19668 27130
rect 19616 27066 19668 27072
rect 19812 27062 19840 27338
rect 20168 27328 20220 27334
rect 20260 27328 20312 27334
rect 20168 27270 20220 27276
rect 20258 27296 20260 27305
rect 20312 27296 20314 27305
rect 20180 27130 20208 27270
rect 20258 27231 20314 27240
rect 20168 27124 20220 27130
rect 20168 27066 20220 27072
rect 19800 27056 19852 27062
rect 19800 26998 19852 27004
rect 19524 26988 19576 26994
rect 19524 26930 19576 26936
rect 20168 26988 20220 26994
rect 20168 26930 20220 26936
rect 20074 26888 20130 26897
rect 20074 26823 20076 26832
rect 20128 26823 20130 26832
rect 20076 26794 20128 26800
rect 19432 26784 19484 26790
rect 19432 26726 19484 26732
rect 19800 26784 19852 26790
rect 19800 26726 19852 26732
rect 17960 26580 18012 26586
rect 17960 26522 18012 26528
rect 19812 26382 19840 26726
rect 20180 26586 20208 26930
rect 20364 26858 20392 27406
rect 20536 27396 20588 27402
rect 20640 27384 20668 27882
rect 20588 27356 20668 27384
rect 20536 27338 20588 27344
rect 20444 26988 20496 26994
rect 20444 26930 20496 26936
rect 20352 26852 20404 26858
rect 20352 26794 20404 26800
rect 20364 26586 20392 26794
rect 20168 26580 20220 26586
rect 20168 26522 20220 26528
rect 20352 26580 20404 26586
rect 20352 26522 20404 26528
rect 12992 26376 13044 26382
rect 12992 26318 13044 26324
rect 13084 26376 13136 26382
rect 13084 26318 13136 26324
rect 13176 26376 13228 26382
rect 13176 26318 13228 26324
rect 19800 26376 19852 26382
rect 19800 26318 19852 26324
rect 12860 25792 12940 25820
rect 12808 25774 12860 25780
rect 12636 25294 12664 25774
rect 12624 25288 12676 25294
rect 12624 25230 12676 25236
rect 12716 25288 12768 25294
rect 12716 25230 12768 25236
rect 12532 24744 12584 24750
rect 12532 24686 12584 24692
rect 12728 24342 12756 25230
rect 12716 24336 12768 24342
rect 12716 24278 12768 24284
rect 12440 24064 12492 24070
rect 12440 24006 12492 24012
rect 12728 23730 12756 24278
rect 12716 23724 12768 23730
rect 12716 23666 12768 23672
rect 12348 23656 12400 23662
rect 12348 23598 12400 23604
rect 12728 23322 12756 23666
rect 12820 23662 12848 25774
rect 13004 25498 13032 26318
rect 13188 26042 13216 26318
rect 20180 26246 20208 26522
rect 20456 26450 20484 26930
rect 20444 26444 20496 26450
rect 20444 26386 20496 26392
rect 20168 26240 20220 26246
rect 20168 26182 20220 26188
rect 20444 26240 20496 26246
rect 20444 26182 20496 26188
rect 13176 26036 13228 26042
rect 13176 25978 13228 25984
rect 12992 25492 13044 25498
rect 12992 25434 13044 25440
rect 13004 24698 13032 25434
rect 13188 25362 13216 25978
rect 20456 25906 20484 26182
rect 20444 25900 20496 25906
rect 20444 25842 20496 25848
rect 20536 25696 20588 25702
rect 20640 25684 20668 27356
rect 20916 25906 20944 28086
rect 21008 27674 21036 28426
rect 21180 28076 21232 28082
rect 21180 28018 21232 28024
rect 20996 27668 21048 27674
rect 20996 27610 21048 27616
rect 21192 27402 21220 28018
rect 21468 27606 21496 28426
rect 22008 28416 22060 28422
rect 22008 28358 22060 28364
rect 21916 28144 21968 28150
rect 21916 28086 21968 28092
rect 21456 27600 21508 27606
rect 21456 27542 21508 27548
rect 21640 27464 21692 27470
rect 21640 27406 21692 27412
rect 21180 27396 21232 27402
rect 21180 27338 21232 27344
rect 20994 27296 21050 27305
rect 20994 27231 21050 27240
rect 21008 26994 21036 27231
rect 21652 26994 21680 27406
rect 21928 27402 21956 28086
rect 21916 27396 21968 27402
rect 21916 27338 21968 27344
rect 22020 27130 22048 28358
rect 22376 28076 22428 28082
rect 22376 28018 22428 28024
rect 22008 27124 22060 27130
rect 22008 27066 22060 27072
rect 20996 26988 21048 26994
rect 20996 26930 21048 26936
rect 21640 26988 21692 26994
rect 21640 26930 21692 26936
rect 22192 26988 22244 26994
rect 22192 26930 22244 26936
rect 20996 26852 21048 26858
rect 20996 26794 21048 26800
rect 21008 26586 21036 26794
rect 20996 26580 21048 26586
rect 20996 26522 21048 26528
rect 21652 26450 21680 26930
rect 21640 26444 21692 26450
rect 21640 26386 21692 26392
rect 20904 25900 20956 25906
rect 20904 25842 20956 25848
rect 22008 25900 22060 25906
rect 22008 25842 22060 25848
rect 20588 25656 20668 25684
rect 20536 25638 20588 25644
rect 17408 25492 17460 25498
rect 17408 25434 17460 25440
rect 13176 25356 13228 25362
rect 13176 25298 13228 25304
rect 15568 25288 15620 25294
rect 15568 25230 15620 25236
rect 15660 25288 15712 25294
rect 15660 25230 15712 25236
rect 15936 25288 15988 25294
rect 15936 25230 15988 25236
rect 15580 24818 15608 25230
rect 15672 24954 15700 25230
rect 15660 24948 15712 24954
rect 15660 24890 15712 24896
rect 15672 24818 15700 24890
rect 15948 24886 15976 25230
rect 16120 25220 16172 25226
rect 16120 25162 16172 25168
rect 15936 24880 15988 24886
rect 15936 24822 15988 24828
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 15568 24812 15620 24818
rect 15568 24754 15620 24760
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 12912 24670 13032 24698
rect 12912 23730 12940 24670
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 13004 24206 13032 24550
rect 14844 24410 14872 24754
rect 15672 24410 15700 24754
rect 15948 24750 15976 24822
rect 16132 24818 16160 25162
rect 16948 25152 17000 25158
rect 16948 25094 17000 25100
rect 17132 25152 17184 25158
rect 17132 25094 17184 25100
rect 16856 24948 16908 24954
rect 16856 24890 16908 24896
rect 16120 24812 16172 24818
rect 16120 24754 16172 24760
rect 15936 24744 15988 24750
rect 15936 24686 15988 24692
rect 16120 24676 16172 24682
rect 16120 24618 16172 24624
rect 15844 24608 15896 24614
rect 15844 24550 15896 24556
rect 14832 24404 14884 24410
rect 14832 24346 14884 24352
rect 15660 24404 15712 24410
rect 15660 24346 15712 24352
rect 14188 24336 14240 24342
rect 14188 24278 14240 24284
rect 12992 24200 13044 24206
rect 12992 24142 13044 24148
rect 13544 24064 13596 24070
rect 13544 24006 13596 24012
rect 13556 23798 13584 24006
rect 13544 23792 13596 23798
rect 13544 23734 13596 23740
rect 12900 23724 12952 23730
rect 12900 23666 12952 23672
rect 12808 23656 12860 23662
rect 12808 23598 12860 23604
rect 12716 23316 12768 23322
rect 12716 23258 12768 23264
rect 12912 23186 12940 23666
rect 13544 23656 13596 23662
rect 13544 23598 13596 23604
rect 13176 23588 13228 23594
rect 13176 23530 13228 23536
rect 12164 23180 12216 23186
rect 12164 23122 12216 23128
rect 12900 23180 12952 23186
rect 12900 23122 12952 23128
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12716 22976 12768 22982
rect 12716 22918 12768 22924
rect 12636 22642 12664 22918
rect 12624 22636 12676 22642
rect 12624 22578 12676 22584
rect 12636 22234 12664 22578
rect 12624 22228 12676 22234
rect 12624 22170 12676 22176
rect 9588 22024 9640 22030
rect 9588 21966 9640 21972
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 11888 22024 11940 22030
rect 11888 21966 11940 21972
rect 12164 22024 12216 22030
rect 12164 21966 12216 21972
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 9496 19780 9548 19786
rect 9496 19722 9548 19728
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 9508 17678 9536 18022
rect 9600 17882 9628 21966
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 11520 21004 11572 21010
rect 11520 20946 11572 20952
rect 11152 20936 11204 20942
rect 11152 20878 11204 20884
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 11164 20534 11192 20878
rect 11152 20528 11204 20534
rect 11152 20470 11204 20476
rect 11348 20466 11376 20878
rect 11532 20534 11560 20946
rect 11612 20936 11664 20942
rect 11612 20878 11664 20884
rect 11624 20602 11652 20878
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 11520 20528 11572 20534
rect 11520 20470 11572 20476
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 11244 20460 11296 20466
rect 11244 20402 11296 20408
rect 11336 20460 11388 20466
rect 11336 20402 11388 20408
rect 11072 20262 11100 20402
rect 11256 20330 11284 20402
rect 11244 20324 11296 20330
rect 11244 20266 11296 20272
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 11612 19916 11664 19922
rect 11612 19858 11664 19864
rect 9772 19236 9824 19242
rect 9772 19178 9824 19184
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9692 18290 9720 18566
rect 9784 18358 9812 19178
rect 9772 18352 9824 18358
rect 9772 18294 9824 18300
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9680 18148 9732 18154
rect 9680 18090 9732 18096
rect 9588 17876 9640 17882
rect 9588 17818 9640 17824
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 9508 16522 9536 17614
rect 9692 17202 9720 18090
rect 9784 17202 9812 18294
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 9876 17678 9904 18226
rect 10048 18216 10100 18222
rect 10048 18158 10100 18164
rect 10060 17746 10088 18158
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 10060 17338 10088 17682
rect 10600 17536 10652 17542
rect 10600 17478 10652 17484
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 10232 17060 10284 17066
rect 10232 17002 10284 17008
rect 10244 16590 10272 17002
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 9496 16516 9548 16522
rect 9496 16458 9548 16464
rect 10244 16250 10272 16526
rect 10232 16244 10284 16250
rect 10232 16186 10284 16192
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 9312 15904 9364 15910
rect 9312 15846 9364 15852
rect 9324 15502 9352 15846
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9600 15162 9628 16050
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9692 15502 9720 15846
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9876 15434 9904 16050
rect 10612 16046 10640 17478
rect 11624 17202 11652 19858
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 11624 16726 11652 17138
rect 11612 16720 11664 16726
rect 11612 16662 11664 16668
rect 11716 16114 11744 21830
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 12084 21010 12112 21490
rect 12176 21146 12204 21966
rect 12164 21140 12216 21146
rect 12164 21082 12216 21088
rect 12072 21004 12124 21010
rect 12072 20946 12124 20952
rect 12544 20942 12572 21966
rect 12728 21894 12756 22918
rect 13188 22642 13216 23530
rect 13176 22636 13228 22642
rect 13176 22578 13228 22584
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12808 21004 12860 21010
rect 12808 20946 12860 20952
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 11888 20868 11940 20874
rect 11888 20810 11940 20816
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11808 18290 11836 20402
rect 11900 19718 11928 20810
rect 12256 20528 12308 20534
rect 12256 20470 12308 20476
rect 12164 20324 12216 20330
rect 12164 20266 12216 20272
rect 11888 19712 11940 19718
rect 11888 19654 11940 19660
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11796 18148 11848 18154
rect 11796 18090 11848 18096
rect 11808 17542 11836 18090
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11900 16674 11928 19654
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 11808 16646 11928 16674
rect 11992 16658 12020 18022
rect 12176 17882 12204 20266
rect 12268 20262 12296 20470
rect 12348 20460 12400 20466
rect 12348 20402 12400 20408
rect 12440 20460 12492 20466
rect 12440 20402 12492 20408
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 12268 19718 12296 20198
rect 12360 19990 12388 20402
rect 12452 20058 12480 20402
rect 12440 20052 12492 20058
rect 12440 19994 12492 20000
rect 12348 19984 12400 19990
rect 12348 19926 12400 19932
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12268 18222 12296 19654
rect 12360 18902 12388 19926
rect 12544 19922 12572 20878
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12440 19780 12492 19786
rect 12440 19722 12492 19728
rect 12452 19446 12480 19722
rect 12440 19440 12492 19446
rect 12440 19382 12492 19388
rect 12544 19378 12572 19858
rect 12636 19514 12664 20334
rect 12820 19854 12848 20946
rect 13188 20942 13216 22578
rect 13556 22094 13584 23598
rect 14200 23186 14228 24278
rect 14372 24200 14424 24206
rect 14372 24142 14424 24148
rect 15660 24200 15712 24206
rect 15660 24142 15712 24148
rect 14188 23180 14240 23186
rect 14188 23122 14240 23128
rect 14188 22432 14240 22438
rect 14188 22374 14240 22380
rect 13464 22066 13584 22094
rect 13176 20936 13228 20942
rect 13176 20878 13228 20884
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13280 20058 13308 20402
rect 13268 20052 13320 20058
rect 13268 19994 13320 20000
rect 12808 19848 12860 19854
rect 12728 19808 12808 19836
rect 12624 19508 12676 19514
rect 12624 19450 12676 19456
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 12636 19258 12664 19450
rect 12728 19310 12756 19808
rect 13464 19836 13492 22066
rect 14096 21888 14148 21894
rect 14096 21830 14148 21836
rect 14108 21622 14136 21830
rect 14096 21616 14148 21622
rect 14096 21558 14148 21564
rect 14004 21480 14056 21486
rect 14004 21422 14056 21428
rect 13820 21412 13872 21418
rect 13820 21354 13872 21360
rect 13544 20936 13596 20942
rect 13596 20896 13676 20924
rect 13544 20878 13596 20884
rect 13544 20800 13596 20806
rect 13544 20742 13596 20748
rect 13556 20534 13584 20742
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 13542 20360 13598 20369
rect 13542 20295 13598 20304
rect 13556 20262 13584 20295
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 13648 19854 13676 20896
rect 13832 20602 13860 21354
rect 13912 21344 13964 21350
rect 13912 21286 13964 21292
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 13924 20505 13952 21286
rect 14016 20913 14044 21422
rect 14096 20936 14148 20942
rect 14002 20904 14058 20913
rect 14096 20878 14148 20884
rect 14002 20839 14058 20848
rect 13910 20496 13966 20505
rect 13820 20460 13872 20466
rect 13910 20431 13966 20440
rect 13820 20402 13872 20408
rect 13728 20324 13780 20330
rect 13728 20266 13780 20272
rect 13740 20058 13768 20266
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 12808 19790 12860 19796
rect 13280 19808 13492 19836
rect 13636 19848 13688 19854
rect 13280 19446 13308 19808
rect 13636 19790 13688 19796
rect 13268 19440 13320 19446
rect 13268 19382 13320 19388
rect 12452 19230 12664 19258
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 12348 18896 12400 18902
rect 12348 18838 12400 18844
rect 12452 18426 12480 19230
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12544 18426 12572 19110
rect 12900 18760 12952 18766
rect 12900 18702 12952 18708
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12728 18426 12756 18566
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12532 18420 12584 18426
rect 12532 18362 12584 18368
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 12164 17876 12216 17882
rect 12164 17818 12216 17824
rect 12256 17876 12308 17882
rect 12256 17818 12308 17824
rect 12176 17785 12204 17818
rect 12162 17776 12218 17785
rect 12162 17711 12218 17720
rect 12072 17536 12124 17542
rect 12072 17478 12124 17484
rect 11980 16652 12032 16658
rect 11808 16182 11836 16646
rect 11980 16594 12032 16600
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11796 16176 11848 16182
rect 11796 16118 11848 16124
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 10048 16040 10100 16046
rect 10048 15982 10100 15988
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 9864 15428 9916 15434
rect 9864 15370 9916 15376
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9876 15026 9904 15370
rect 10060 15026 10088 15982
rect 11716 15502 11744 16050
rect 11808 15502 11836 16118
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 8668 15020 8720 15026
rect 8668 14962 8720 14968
rect 9864 15020 9916 15026
rect 9864 14962 9916 14968
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 7932 14884 7984 14890
rect 7932 14826 7984 14832
rect 7944 14006 7972 14826
rect 7932 14000 7984 14006
rect 7932 13942 7984 13948
rect 7748 12164 7800 12170
rect 7748 12106 7800 12112
rect 7760 11762 7788 12106
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7656 10736 7708 10742
rect 7656 10678 7708 10684
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7392 10062 7420 10610
rect 7668 10062 7696 10678
rect 7944 10130 7972 13942
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8312 13394 8340 13806
rect 8588 13802 8616 14894
rect 8576 13796 8628 13802
rect 8576 13738 8628 13744
rect 8588 13530 8616 13738
rect 8680 13530 8708 14962
rect 10520 14890 10548 15438
rect 10692 15088 10744 15094
rect 10692 15030 10744 15036
rect 10508 14884 10560 14890
rect 10508 14826 10560 14832
rect 10520 13938 10548 14826
rect 10704 13977 10732 15030
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11348 14346 11376 14758
rect 11336 14340 11388 14346
rect 11336 14282 11388 14288
rect 11348 14074 11376 14282
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 10690 13968 10746 13977
rect 10508 13932 10560 13938
rect 10690 13903 10746 13912
rect 10508 13874 10560 13880
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 8944 13728 8996 13734
rect 8944 13670 8996 13676
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8956 13326 8984 13670
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 8036 12850 8064 13126
rect 8024 12844 8076 12850
rect 8128 12832 8156 13262
rect 8300 13252 8352 13258
rect 8300 13194 8352 13200
rect 8312 12986 8340 13194
rect 9232 12986 9260 13262
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 8208 12844 8260 12850
rect 8128 12804 8208 12832
rect 8024 12786 8076 12792
rect 8208 12786 8260 12792
rect 8036 12730 8064 12786
rect 8036 12702 8156 12730
rect 8128 10810 8156 12702
rect 8220 11898 8248 12786
rect 8312 12306 8340 12922
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 9784 12209 9812 12718
rect 9770 12200 9826 12209
rect 9770 12135 9826 12144
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 9784 11082 9812 12135
rect 10874 12064 10930 12073
rect 10874 11999 10930 12008
rect 10508 11824 10560 11830
rect 10508 11766 10560 11772
rect 10230 11384 10286 11393
rect 10048 11348 10100 11354
rect 10230 11319 10232 11328
rect 10048 11290 10100 11296
rect 10284 11319 10286 11328
rect 10232 11290 10284 11296
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7392 9586 7420 9998
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7484 9654 7512 9930
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7012 8356 7064 8362
rect 7012 8298 7064 8304
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6920 7404 6972 7410
rect 7024 7392 7052 8298
rect 6972 7364 7052 7392
rect 6920 7346 6972 7352
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5552 7002 5580 7278
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5460 6322 5488 6870
rect 5644 6866 5672 7278
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5816 6792 5868 6798
rect 5920 6780 5948 7142
rect 6288 6866 6316 7346
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 5868 6752 5948 6780
rect 5816 6734 5868 6740
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5920 6254 5948 6752
rect 6288 6254 6316 6802
rect 6472 6458 6500 6802
rect 6644 6792 6696 6798
rect 6696 6752 6776 6780
rect 6644 6734 6696 6740
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6748 6610 6776 6752
rect 6932 6730 6960 7346
rect 7116 6798 7144 8434
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 6920 6724 6972 6730
rect 6920 6666 6972 6672
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6472 6322 6500 6394
rect 6656 6322 6684 6598
rect 6748 6582 6960 6610
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 6276 6248 6328 6254
rect 6276 6190 6328 6196
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 6932 5914 6960 6582
rect 7116 6458 7144 6734
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7208 6390 7236 7822
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7196 6384 7248 6390
rect 7196 6326 7248 6332
rect 7300 6322 7328 7482
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7392 5914 7420 9522
rect 7484 8498 7512 9590
rect 8128 9586 8156 10202
rect 8220 10198 8248 10406
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8220 9738 8248 10134
rect 8312 9994 8340 10542
rect 8404 10198 8432 10610
rect 8864 10266 8892 10610
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 8220 9722 8340 9738
rect 8220 9716 8352 9722
rect 8220 9710 8300 9716
rect 8300 9658 8352 9664
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7944 8974 7972 9454
rect 8128 8974 8156 9522
rect 8220 9178 8248 9590
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 7944 8634 7972 8910
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 7484 8294 7512 8434
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 8036 8022 8064 8434
rect 8024 8016 8076 8022
rect 8024 7958 8076 7964
rect 8220 7410 8248 9114
rect 8404 8634 8432 10134
rect 9140 9994 9168 10542
rect 9324 10266 9352 10610
rect 9968 10266 9996 10950
rect 10060 10606 10088 11290
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 10152 10062 10180 11154
rect 10520 11150 10548 11766
rect 10888 11762 10916 11999
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10598 11248 10654 11257
rect 10598 11183 10654 11192
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10612 10470 10640 11183
rect 10796 11150 10824 11290
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10888 10810 10916 11086
rect 11072 11082 11100 13806
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11164 11218 11192 12038
rect 11348 11898 11376 12174
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 11072 10674 11100 11018
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10612 10266 10640 10406
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 9128 9988 9180 9994
rect 9128 9930 9180 9936
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 8772 9722 8800 9862
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 9140 8498 9168 9930
rect 9588 9920 9640 9926
rect 9586 9888 9588 9897
rect 9680 9920 9732 9926
rect 9640 9888 9642 9897
rect 9680 9862 9732 9868
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9586 9823 9642 9832
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9140 8090 9168 8434
rect 9324 8090 9352 8434
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8220 6798 8248 7346
rect 8404 6798 8432 7414
rect 8588 7342 8616 7822
rect 9600 7546 9628 9823
rect 9692 9450 9720 9862
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9692 8362 9720 9386
rect 9680 8356 9732 8362
rect 9680 8298 9732 8304
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9784 7478 9812 9862
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 10060 8498 10088 9454
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 10152 8634 10180 8842
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10060 7478 10088 8434
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 9772 7472 9824 7478
rect 9772 7414 9824 7420
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8588 7002 8616 7278
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 9140 6798 9168 7346
rect 9416 7002 9444 7346
rect 9784 7206 9812 7414
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 10060 6934 10088 7414
rect 10048 6928 10100 6934
rect 10048 6870 10100 6876
rect 10152 6798 10180 7754
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 7564 6724 7616 6730
rect 7564 6666 7616 6672
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 7576 2650 7604 6666
rect 8404 6254 8432 6734
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9508 6322 9536 6598
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8680 2650 8708 5850
rect 10244 5778 10272 8910
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10336 6730 10364 7346
rect 10520 7002 10548 8434
rect 10612 8430 10640 10202
rect 11164 10062 11192 11154
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11348 10985 11376 11086
rect 11334 10976 11390 10985
rect 11334 10911 11390 10920
rect 11348 10538 11376 10911
rect 11440 10674 11468 12786
rect 11808 12714 11836 14962
rect 11900 13462 11928 16526
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 11992 14074 12020 15438
rect 12084 15162 12112 17478
rect 12268 16590 12296 17818
rect 12452 17626 12480 18362
rect 12532 18284 12584 18290
rect 12716 18284 12768 18290
rect 12532 18226 12584 18232
rect 12636 18244 12716 18272
rect 12544 17882 12572 18226
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12360 17598 12480 17626
rect 12360 17542 12388 17598
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12164 16516 12216 16522
rect 12164 16458 12216 16464
rect 12176 15706 12204 16458
rect 12164 15700 12216 15706
rect 12164 15642 12216 15648
rect 12360 15162 12388 16730
rect 12072 15156 12124 15162
rect 12072 15098 12124 15104
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12452 15026 12480 17598
rect 12532 17604 12584 17610
rect 12532 17546 12584 17552
rect 12544 16590 12572 17546
rect 12636 16998 12664 18244
rect 12716 18226 12768 18232
rect 12912 18222 12940 18702
rect 13004 18290 13032 19246
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13188 18358 13216 18566
rect 13176 18352 13228 18358
rect 13176 18294 13228 18300
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 12900 18216 12952 18222
rect 12820 18176 12900 18204
rect 12820 17746 12848 18176
rect 12900 18158 12952 18164
rect 12898 17776 12954 17785
rect 12808 17740 12860 17746
rect 12898 17711 12954 17720
rect 12808 17682 12860 17688
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 12636 16590 12664 16934
rect 12728 16658 12756 17070
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12072 15020 12124 15026
rect 12440 15020 12492 15026
rect 12124 14980 12204 15008
rect 12072 14962 12124 14968
rect 12072 14884 12124 14890
rect 12072 14826 12124 14832
rect 12084 14618 12112 14826
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12176 14090 12204 14980
rect 12440 14962 12492 14968
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 12084 14062 12204 14090
rect 12268 14074 12296 14758
rect 12256 14068 12308 14074
rect 12084 13954 12112 14062
rect 12256 14010 12308 14016
rect 11992 13926 12112 13954
rect 11992 13870 12020 13926
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 12440 13864 12492 13870
rect 12544 13852 12572 16526
rect 12728 16182 12756 16594
rect 12716 16176 12768 16182
rect 12716 16118 12768 16124
rect 12912 15026 12940 17711
rect 13280 17270 13308 19382
rect 13648 19174 13676 19790
rect 13728 19236 13780 19242
rect 13728 19178 13780 19184
rect 13636 19168 13688 19174
rect 13636 19110 13688 19116
rect 13740 18766 13768 19178
rect 13832 18970 13860 20402
rect 14016 19990 14044 20839
rect 14004 19984 14056 19990
rect 14004 19926 14056 19932
rect 13912 19848 13964 19854
rect 13912 19790 13964 19796
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13924 18834 13952 19790
rect 14004 19780 14056 19786
rect 14108 19768 14136 20878
rect 14200 19922 14228 22374
rect 14280 22228 14332 22234
rect 14280 22170 14332 22176
rect 14292 21962 14320 22170
rect 14384 22098 14412 24142
rect 15672 23866 15700 24142
rect 15660 23860 15712 23866
rect 15660 23802 15712 23808
rect 15016 23520 15068 23526
rect 15016 23462 15068 23468
rect 14556 23180 14608 23186
rect 14556 23122 14608 23128
rect 14372 22092 14424 22098
rect 14372 22034 14424 22040
rect 14568 21978 14596 23122
rect 15028 23118 15056 23462
rect 15016 23112 15068 23118
rect 15016 23054 15068 23060
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 14280 21956 14332 21962
rect 14280 21898 14332 21904
rect 14384 21950 14596 21978
rect 14660 21962 14688 22918
rect 14740 22092 14792 22098
rect 14740 22034 14792 22040
rect 14648 21956 14700 21962
rect 14292 21690 14320 21898
rect 14280 21684 14332 21690
rect 14280 21626 14332 21632
rect 14384 21486 14412 21950
rect 14648 21898 14700 21904
rect 14556 21888 14608 21894
rect 14556 21830 14608 21836
rect 14372 21480 14424 21486
rect 14372 21422 14424 21428
rect 14464 21344 14516 21350
rect 14464 21286 14516 21292
rect 14372 20936 14424 20942
rect 14372 20878 14424 20884
rect 14280 20800 14332 20806
rect 14280 20742 14332 20748
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 14056 19740 14136 19768
rect 14004 19722 14056 19728
rect 14016 19310 14044 19722
rect 14096 19440 14148 19446
rect 14096 19382 14148 19388
rect 14004 19304 14056 19310
rect 14004 19246 14056 19252
rect 14108 19122 14136 19382
rect 14016 19094 14136 19122
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 13924 18358 13952 18770
rect 13912 18352 13964 18358
rect 13912 18294 13964 18300
rect 14016 18204 14044 19094
rect 14096 18692 14148 18698
rect 14096 18634 14148 18640
rect 13924 18176 14044 18204
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 13268 17264 13320 17270
rect 13268 17206 13320 17212
rect 13268 17060 13320 17066
rect 13268 17002 13320 17008
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 13188 16250 13216 16526
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 13280 14414 13308 17002
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13372 15570 13400 16390
rect 13360 15564 13412 15570
rect 13360 15506 13412 15512
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 13372 14278 13400 14962
rect 13464 14414 13492 17818
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13832 16114 13860 17138
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13832 15706 13860 15846
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12992 14272 13044 14278
rect 12992 14214 13044 14220
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 12820 13938 12848 14214
rect 13004 14006 13032 14214
rect 12992 14000 13044 14006
rect 12992 13942 13044 13948
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12492 13824 12572 13852
rect 12440 13806 12492 13812
rect 12084 13530 12112 13806
rect 12348 13796 12400 13802
rect 12348 13738 12400 13744
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 11888 13456 11940 13462
rect 11888 13398 11940 13404
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 12176 12866 12204 13670
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 12268 12986 12296 13262
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12084 12764 12112 12854
rect 12176 12838 12296 12866
rect 12360 12850 12388 13738
rect 13372 13734 13400 14214
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12084 12736 12204 12764
rect 11796 12708 11848 12714
rect 11796 12650 11848 12656
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 11520 12096 11572 12102
rect 11520 12038 11572 12044
rect 11532 11898 11560 12038
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11978 11792 12034 11801
rect 11704 11756 11756 11762
rect 11978 11727 11980 11736
rect 11704 11698 11756 11704
rect 12032 11727 12034 11736
rect 11980 11698 12032 11704
rect 11716 11665 11744 11698
rect 11702 11656 11758 11665
rect 11702 11591 11758 11600
rect 12084 11354 12112 12582
rect 12176 11762 12204 12736
rect 12268 12730 12296 12838
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12268 12702 12388 12730
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 12268 11762 12296 12242
rect 12164 11756 12216 11762
rect 12164 11698 12216 11704
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 12176 11626 12204 11698
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 11520 11280 11572 11286
rect 11520 11222 11572 11228
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11532 10996 11560 11222
rect 11624 11121 11652 11222
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11610 11112 11666 11121
rect 11610 11047 11666 11056
rect 11716 11070 11928 11098
rect 11716 10996 11744 11070
rect 11900 11014 11928 11070
rect 11532 10968 11744 10996
rect 11796 11008 11848 11014
rect 11796 10950 11848 10956
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11440 9994 11468 10610
rect 11808 10606 11836 10950
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11624 10033 11652 10542
rect 11610 10024 11666 10033
rect 11428 9988 11480 9994
rect 11610 9959 11666 9968
rect 11428 9930 11480 9936
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11072 9042 11100 9862
rect 11808 9178 11836 10542
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10796 8498 10824 8570
rect 11072 8566 11100 8978
rect 11900 8634 11928 10610
rect 11992 9994 12020 11154
rect 12084 11082 12112 11290
rect 12254 11248 12310 11257
rect 12254 11183 12310 11192
rect 12268 11150 12296 11183
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 11980 9988 12032 9994
rect 11980 9930 12032 9936
rect 12084 9110 12112 11018
rect 12176 10810 12204 11018
rect 12360 10810 12388 12702
rect 12452 12345 12480 13466
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12624 13252 12676 13258
rect 12624 13194 12676 13200
rect 12636 12986 12664 13194
rect 12820 13190 12848 13330
rect 13924 13326 13952 18176
rect 14108 18086 14136 18634
rect 14200 18290 14228 19858
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14096 18080 14148 18086
rect 14096 18022 14148 18028
rect 14004 16992 14056 16998
rect 14004 16934 14056 16940
rect 14016 15978 14044 16934
rect 14108 16250 14136 18022
rect 14200 17678 14228 18226
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 14096 16244 14148 16250
rect 14096 16186 14148 16192
rect 14292 15994 14320 20742
rect 14384 19446 14412 20878
rect 14476 20806 14504 21286
rect 14568 20942 14596 21830
rect 14648 21480 14700 21486
rect 14648 21422 14700 21428
rect 14556 20936 14608 20942
rect 14556 20878 14608 20884
rect 14464 20800 14516 20806
rect 14464 20742 14516 20748
rect 14554 20496 14610 20505
rect 14554 20431 14610 20440
rect 14568 20398 14596 20431
rect 14556 20392 14608 20398
rect 14556 20334 14608 20340
rect 14372 19440 14424 19446
rect 14372 19382 14424 19388
rect 14372 19304 14424 19310
rect 14372 19246 14424 19252
rect 14384 18766 14412 19246
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14476 18766 14504 19110
rect 14660 18850 14688 21422
rect 14752 21350 14780 22034
rect 15028 22030 15056 23054
rect 15016 22024 15068 22030
rect 15016 21966 15068 21972
rect 15292 22024 15344 22030
rect 15292 21966 15344 21972
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14844 21486 14872 21830
rect 15028 21690 15056 21966
rect 15016 21684 15068 21690
rect 15016 21626 15068 21632
rect 15304 21554 15332 21966
rect 15292 21548 15344 21554
rect 15292 21490 15344 21496
rect 14832 21480 14884 21486
rect 14832 21422 14884 21428
rect 14936 21406 15240 21434
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 14832 21344 14884 21350
rect 14936 21298 14964 21406
rect 14884 21292 14964 21298
rect 14832 21286 14964 21292
rect 15016 21344 15068 21350
rect 15016 21286 15068 21292
rect 14844 21270 14964 21286
rect 15028 21026 15056 21286
rect 15212 21146 15240 21406
rect 15384 21412 15436 21418
rect 15384 21354 15436 21360
rect 15108 21140 15160 21146
rect 15108 21082 15160 21088
rect 15200 21140 15252 21146
rect 15200 21082 15252 21088
rect 15120 21049 15148 21082
rect 14752 21010 15056 21026
rect 14740 21004 15056 21010
rect 14792 20998 15056 21004
rect 15106 21040 15162 21049
rect 15106 20975 15162 20984
rect 14740 20946 14792 20952
rect 14924 20936 14976 20942
rect 14924 20878 14976 20884
rect 14740 20868 14792 20874
rect 14740 20810 14792 20816
rect 14752 20398 14780 20810
rect 14936 20602 14964 20878
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 15396 20788 15424 21354
rect 15476 20800 15528 20806
rect 15396 20760 15476 20788
rect 14924 20596 14976 20602
rect 14924 20538 14976 20544
rect 15108 20596 15160 20602
rect 15108 20538 15160 20544
rect 15016 20460 15068 20466
rect 15016 20402 15068 20408
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 14752 19922 14780 20334
rect 15028 19990 15056 20402
rect 15016 19984 15068 19990
rect 15016 19926 15068 19932
rect 14740 19916 14792 19922
rect 14740 19858 14792 19864
rect 15028 19514 15056 19926
rect 15120 19786 15148 20538
rect 15212 20466 15240 20742
rect 15396 20466 15424 20760
rect 15476 20742 15528 20748
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15292 20460 15344 20466
rect 15292 20402 15344 20408
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15476 20460 15528 20466
rect 15476 20402 15528 20408
rect 15108 19780 15160 19786
rect 15108 19722 15160 19728
rect 15016 19508 15068 19514
rect 15016 19450 15068 19456
rect 15120 19446 15148 19722
rect 15212 19718 15240 20402
rect 15304 20058 15332 20402
rect 15488 20369 15516 20402
rect 15474 20360 15530 20369
rect 15474 20295 15530 20304
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 15200 19712 15252 19718
rect 15200 19654 15252 19660
rect 15108 19440 15160 19446
rect 15108 19382 15160 19388
rect 14660 18822 14780 18850
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14476 18578 14504 18702
rect 14384 18550 14504 18578
rect 14384 17202 14412 18550
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14476 17814 14504 18022
rect 14464 17808 14516 17814
rect 14464 17750 14516 17756
rect 14476 17202 14504 17750
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 14660 17202 14688 17682
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 14556 17060 14608 17066
rect 14556 17002 14608 17008
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14384 16522 14412 16934
rect 14372 16516 14424 16522
rect 14424 16476 14504 16504
rect 14372 16458 14424 16464
rect 14476 16114 14504 16476
rect 14568 16454 14596 17002
rect 14556 16448 14608 16454
rect 14556 16390 14608 16396
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 14004 15972 14056 15978
rect 14292 15966 14412 15994
rect 14004 15914 14056 15920
rect 14096 15904 14148 15910
rect 14096 15846 14148 15852
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14004 14476 14056 14482
rect 14004 14418 14056 14424
rect 14016 13394 14044 14418
rect 14004 13388 14056 13394
rect 14004 13330 14056 13336
rect 13912 13320 13964 13326
rect 13912 13262 13964 13268
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 12728 12918 12756 13126
rect 12716 12912 12768 12918
rect 12716 12854 12768 12860
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 12438 12336 12494 12345
rect 12438 12271 12440 12280
rect 12492 12271 12494 12280
rect 12532 12300 12584 12306
rect 12440 12242 12492 12248
rect 12532 12242 12584 12248
rect 12544 12084 12572 12242
rect 12636 12102 12664 12786
rect 12820 12434 12848 13126
rect 12820 12406 12940 12434
rect 12808 12300 12860 12306
rect 12728 12260 12808 12288
rect 12452 12056 12572 12084
rect 12624 12096 12676 12102
rect 12452 11762 12480 12056
rect 12624 12038 12676 12044
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12440 11756 12492 11762
rect 12440 11698 12492 11704
rect 12452 11354 12480 11698
rect 12544 11354 12572 11766
rect 12728 11626 12756 12260
rect 12808 12242 12860 12248
rect 12912 12186 12940 12406
rect 13358 12336 13414 12345
rect 13358 12271 13414 12280
rect 12820 12170 12940 12186
rect 12808 12164 12940 12170
rect 12860 12158 12940 12164
rect 13268 12164 13320 12170
rect 12808 12106 12860 12112
rect 13268 12106 13320 12112
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 12716 11620 12768 11626
rect 12716 11562 12768 11568
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12268 10130 12296 10610
rect 12348 10532 12400 10538
rect 12348 10474 12400 10480
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 12360 9994 12388 10474
rect 12452 10062 12480 10746
rect 12544 10742 12572 10950
rect 12532 10736 12584 10742
rect 12532 10678 12584 10684
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12348 9988 12400 9994
rect 12348 9930 12400 9936
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12072 9104 12124 9110
rect 12072 9046 12124 9052
rect 12072 8900 12124 8906
rect 12072 8842 12124 8848
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11060 8560 11112 8566
rect 11060 8502 11112 8508
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10796 7886 10824 8434
rect 11808 8022 11836 8434
rect 11992 8090 12020 8434
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 11796 8016 11848 8022
rect 11796 7958 11848 7964
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 11808 7478 11836 7958
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 11796 7472 11848 7478
rect 11796 7414 11848 7420
rect 11992 7410 12020 7890
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 10796 7002 10824 7346
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 10324 6724 10376 6730
rect 10324 6666 10376 6672
rect 10232 5772 10284 5778
rect 10232 5714 10284 5720
rect 10520 5642 10548 6938
rect 10980 6662 11008 7346
rect 11072 6866 11100 7346
rect 11888 7268 11940 7274
rect 11888 7210 11940 7216
rect 11794 7032 11850 7041
rect 11794 6967 11850 6976
rect 11244 6928 11296 6934
rect 11164 6888 11244 6916
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 11072 6458 11100 6802
rect 11164 6730 11192 6888
rect 11244 6870 11296 6876
rect 11426 6896 11482 6905
rect 11426 6831 11482 6840
rect 11440 6798 11468 6831
rect 11808 6798 11836 6967
rect 11900 6934 11928 7210
rect 11888 6928 11940 6934
rect 11888 6870 11940 6876
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11716 6662 11744 6734
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11624 6497 11652 6598
rect 11610 6488 11666 6497
rect 11060 6452 11112 6458
rect 11610 6423 11666 6432
rect 11060 6394 11112 6400
rect 11992 6390 12020 7346
rect 11980 6384 12032 6390
rect 11980 6326 12032 6332
rect 11992 5914 12020 6326
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 10508 5636 10560 5642
rect 10508 5578 10560 5584
rect 11532 5234 11560 5714
rect 12084 5642 12112 8842
rect 12360 8498 12388 8842
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12268 6866 12296 7686
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 12348 6860 12400 6866
rect 12452 6848 12480 9318
rect 12544 7206 12572 10542
rect 12636 9994 12664 10678
rect 12728 10606 12756 11562
rect 12912 10810 12940 12038
rect 13188 11354 13216 12038
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 13096 10985 13124 11086
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 13082 10976 13138 10985
rect 13082 10911 13138 10920
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12992 10532 13044 10538
rect 12992 10474 13044 10480
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12820 10130 12848 10406
rect 12900 10192 12952 10198
rect 12900 10134 12952 10140
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12624 9988 12676 9994
rect 12624 9930 12676 9936
rect 12636 7410 12664 9930
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12820 8974 12848 9862
rect 12912 9586 12940 10134
rect 13004 9586 13032 10474
rect 13096 10198 13124 10911
rect 13084 10192 13136 10198
rect 13084 10134 13136 10140
rect 13096 10062 13124 10134
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12728 8090 12756 8910
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12728 7274 12756 7822
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12400 6820 12480 6848
rect 12348 6802 12400 6808
rect 12164 6792 12216 6798
rect 12544 6746 12572 7142
rect 12622 6896 12678 6905
rect 12622 6831 12624 6840
rect 12676 6831 12678 6840
rect 12624 6802 12676 6808
rect 12164 6734 12216 6740
rect 12176 6458 12204 6734
rect 12348 6724 12400 6730
rect 12348 6666 12400 6672
rect 12452 6718 12572 6746
rect 12360 6633 12388 6666
rect 12346 6624 12402 6633
rect 12346 6559 12402 6568
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12072 5636 12124 5642
rect 12072 5578 12124 5584
rect 12176 5370 12204 6394
rect 12452 6322 12480 6718
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12348 6112 12400 6118
rect 12346 6080 12348 6089
rect 12400 6080 12402 6089
rect 12346 6015 12402 6024
rect 12636 5914 12664 6802
rect 12728 6390 12756 7210
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12820 6798 12848 7142
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12912 6322 12940 7414
rect 12992 7268 13044 7274
rect 12992 7210 13044 7216
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12912 6225 12940 6258
rect 13004 6254 13032 7210
rect 13082 7032 13138 7041
rect 13082 6967 13138 6976
rect 13096 6934 13124 6967
rect 13084 6928 13136 6934
rect 13084 6870 13136 6876
rect 13188 6458 13216 11018
rect 13280 11014 13308 12106
rect 13268 11008 13320 11014
rect 13268 10950 13320 10956
rect 13280 9586 13308 10950
rect 13372 9625 13400 12271
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13542 11792 13598 11801
rect 13542 11727 13598 11736
rect 13358 9616 13414 9625
rect 13268 9580 13320 9586
rect 13358 9551 13414 9560
rect 13268 9522 13320 9528
rect 13280 8072 13308 9522
rect 13372 9382 13400 9551
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13280 8044 13400 8072
rect 13266 7984 13322 7993
rect 13372 7954 13400 8044
rect 13266 7919 13322 7928
rect 13360 7948 13412 7954
rect 13280 7886 13308 7919
rect 13360 7890 13412 7896
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 12992 6248 13044 6254
rect 12898 6216 12954 6225
rect 12992 6190 13044 6196
rect 12898 6151 12954 6160
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 13084 5636 13136 5642
rect 13084 5578 13136 5584
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 13096 5302 13124 5578
rect 13280 5370 13308 7346
rect 13372 7274 13400 7890
rect 13360 7268 13412 7274
rect 13360 7210 13412 7216
rect 13556 7041 13584 11727
rect 13832 11558 13860 11834
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13832 7750 13860 11494
rect 14108 11121 14136 15846
rect 14292 15162 14320 15846
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14384 15094 14412 15966
rect 14372 15088 14424 15094
rect 14278 15056 14334 15065
rect 14372 15030 14424 15036
rect 14278 14991 14280 15000
rect 14332 14991 14334 15000
rect 14280 14962 14332 14968
rect 14752 14958 14780 18822
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 15108 18284 15160 18290
rect 15108 18226 15160 18232
rect 15120 17678 15148 18226
rect 15200 17808 15252 17814
rect 15200 17750 15252 17756
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 14844 16998 14872 17614
rect 15016 17536 15068 17542
rect 15016 17478 15068 17484
rect 14832 16992 14884 16998
rect 14832 16934 14884 16940
rect 15028 16114 15056 17478
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 15120 16250 15148 16390
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 15212 16046 15240 17750
rect 15396 17678 15424 18702
rect 15672 18358 15700 23802
rect 15856 23730 15884 24550
rect 15936 24132 15988 24138
rect 15936 24074 15988 24080
rect 15844 23724 15896 23730
rect 15844 23666 15896 23672
rect 15752 23520 15804 23526
rect 15752 23462 15804 23468
rect 15764 23118 15792 23462
rect 15752 23112 15804 23118
rect 15752 23054 15804 23060
rect 15660 18352 15712 18358
rect 15660 18294 15712 18300
rect 15764 17678 15792 23054
rect 15844 21072 15896 21078
rect 15844 21014 15896 21020
rect 15856 18290 15884 21014
rect 15948 18426 15976 24074
rect 16132 23730 16160 24618
rect 16396 24132 16448 24138
rect 16396 24074 16448 24080
rect 16408 23798 16436 24074
rect 16396 23792 16448 23798
rect 16396 23734 16448 23740
rect 16120 23724 16172 23730
rect 16120 23666 16172 23672
rect 16868 23594 16896 24890
rect 16960 24750 16988 25094
rect 16948 24744 17000 24750
rect 16948 24686 17000 24692
rect 17040 24336 17092 24342
rect 17040 24278 17092 24284
rect 17052 23730 17080 24278
rect 17144 23730 17172 25094
rect 17420 24954 17448 25434
rect 20548 25430 20576 25638
rect 20536 25424 20588 25430
rect 20536 25366 20588 25372
rect 22020 25294 22048 25842
rect 22008 25288 22060 25294
rect 22008 25230 22060 25236
rect 17592 25220 17644 25226
rect 17592 25162 17644 25168
rect 17408 24948 17460 24954
rect 17408 24890 17460 24896
rect 17604 24818 17632 25162
rect 22020 24954 22048 25230
rect 22204 25226 22232 26930
rect 22284 26920 22336 26926
rect 22284 26862 22336 26868
rect 22296 26625 22324 26862
rect 22282 26616 22338 26625
rect 22388 26586 22416 28018
rect 22480 27674 22508 28426
rect 23032 28218 23060 28426
rect 23020 28212 23072 28218
rect 23020 28154 23072 28160
rect 22468 27668 22520 27674
rect 22468 27610 22520 27616
rect 23124 27606 23152 28426
rect 24400 28008 24452 28014
rect 24400 27950 24452 27956
rect 23112 27600 23164 27606
rect 23112 27542 23164 27548
rect 24412 27554 24440 27950
rect 24504 27674 24532 28426
rect 24584 28076 24636 28082
rect 24768 28076 24820 28082
rect 24584 28018 24636 28024
rect 24688 28036 24768 28064
rect 24596 27674 24624 28018
rect 24492 27668 24544 27674
rect 24492 27610 24544 27616
rect 24584 27668 24636 27674
rect 24584 27610 24636 27616
rect 24412 27526 24532 27554
rect 24504 27470 24532 27526
rect 22560 27464 22612 27470
rect 22560 27406 22612 27412
rect 23296 27464 23348 27470
rect 23296 27406 23348 27412
rect 24032 27464 24084 27470
rect 24032 27406 24084 27412
rect 24492 27464 24544 27470
rect 24492 27406 24544 27412
rect 22572 26761 22600 27406
rect 23020 27396 23072 27402
rect 23020 27338 23072 27344
rect 22652 27328 22704 27334
rect 22650 27296 22652 27305
rect 22704 27296 22706 27305
rect 22650 27231 22706 27240
rect 22664 26858 22692 27231
rect 23032 27062 23060 27338
rect 23110 27296 23166 27305
rect 23110 27231 23166 27240
rect 23124 27062 23152 27231
rect 23308 27130 23336 27406
rect 23388 27396 23440 27402
rect 23388 27338 23440 27344
rect 23296 27124 23348 27130
rect 23296 27066 23348 27072
rect 22836 27056 22888 27062
rect 23020 27056 23072 27062
rect 22888 27004 22968 27010
rect 22836 26998 22968 27004
rect 23020 26998 23072 27004
rect 23112 27056 23164 27062
rect 23112 26998 23164 27004
rect 22848 26982 22968 26998
rect 22652 26852 22704 26858
rect 22652 26794 22704 26800
rect 22558 26752 22614 26761
rect 22558 26687 22614 26696
rect 22282 26551 22338 26560
rect 22376 26580 22428 26586
rect 22376 26522 22428 26528
rect 22468 26376 22520 26382
rect 22572 26364 22600 26687
rect 22664 26466 22692 26794
rect 22940 26586 22968 26982
rect 23112 26784 23164 26790
rect 23112 26726 23164 26732
rect 23018 26616 23074 26625
rect 22928 26580 22980 26586
rect 23018 26551 23074 26560
rect 22928 26522 22980 26528
rect 22664 26438 22784 26466
rect 22756 26382 22784 26438
rect 22940 26382 22968 26522
rect 23032 26518 23060 26551
rect 23020 26512 23072 26518
rect 23020 26454 23072 26460
rect 22652 26376 22704 26382
rect 22572 26336 22652 26364
rect 22468 26318 22520 26324
rect 22652 26318 22704 26324
rect 22744 26376 22796 26382
rect 22744 26318 22796 26324
rect 22928 26376 22980 26382
rect 22928 26318 22980 26324
rect 22284 26308 22336 26314
rect 22284 26250 22336 26256
rect 22192 25220 22244 25226
rect 22192 25162 22244 25168
rect 22008 24948 22060 24954
rect 22008 24890 22060 24896
rect 22204 24886 22232 25162
rect 19156 24880 19208 24886
rect 19156 24822 19208 24828
rect 22192 24880 22244 24886
rect 22192 24822 22244 24828
rect 17592 24812 17644 24818
rect 17592 24754 17644 24760
rect 17224 24608 17276 24614
rect 17224 24550 17276 24556
rect 17236 23730 17264 24550
rect 17604 24342 17632 24754
rect 18052 24676 18104 24682
rect 18052 24618 18104 24624
rect 17868 24608 17920 24614
rect 17868 24550 17920 24556
rect 17592 24336 17644 24342
rect 17592 24278 17644 24284
rect 17500 24064 17552 24070
rect 17500 24006 17552 24012
rect 17512 23798 17540 24006
rect 17500 23792 17552 23798
rect 17500 23734 17552 23740
rect 17040 23724 17092 23730
rect 17040 23666 17092 23672
rect 17132 23724 17184 23730
rect 17132 23666 17184 23672
rect 17224 23724 17276 23730
rect 17224 23666 17276 23672
rect 16856 23588 16908 23594
rect 16856 23530 16908 23536
rect 16856 23248 16908 23254
rect 16856 23190 16908 23196
rect 16868 22574 16896 23190
rect 17052 23118 17080 23666
rect 17880 23662 17908 24550
rect 18064 24274 18092 24618
rect 18052 24268 18104 24274
rect 18052 24210 18104 24216
rect 18512 24268 18564 24274
rect 18512 24210 18564 24216
rect 18236 23860 18288 23866
rect 18236 23802 18288 23808
rect 18052 23724 18104 23730
rect 18052 23666 18104 23672
rect 17868 23656 17920 23662
rect 17868 23598 17920 23604
rect 17408 23588 17460 23594
rect 17408 23530 17460 23536
rect 17132 23520 17184 23526
rect 17132 23462 17184 23468
rect 17040 23112 17092 23118
rect 17040 23054 17092 23060
rect 16856 22568 16908 22574
rect 16856 22510 16908 22516
rect 16212 22092 16264 22098
rect 16212 22034 16264 22040
rect 16224 21554 16252 22034
rect 16948 21888 17000 21894
rect 16948 21830 17000 21836
rect 16212 21548 16264 21554
rect 16212 21490 16264 21496
rect 16396 21548 16448 21554
rect 16396 21490 16448 21496
rect 16212 20936 16264 20942
rect 16264 20896 16344 20924
rect 16212 20878 16264 20884
rect 16316 19446 16344 20896
rect 16408 20856 16436 21490
rect 16764 21480 16816 21486
rect 16764 21422 16816 21428
rect 16580 21412 16632 21418
rect 16580 21354 16632 21360
rect 16592 21078 16620 21354
rect 16580 21072 16632 21078
rect 16580 21014 16632 21020
rect 16486 20904 16542 20913
rect 16408 20848 16486 20856
rect 16408 20828 16488 20848
rect 16408 20262 16436 20828
rect 16540 20839 16542 20848
rect 16488 20810 16540 20816
rect 16592 20534 16620 21014
rect 16776 21010 16804 21422
rect 16764 21004 16816 21010
rect 16764 20946 16816 20952
rect 16580 20528 16632 20534
rect 16580 20470 16632 20476
rect 16776 20466 16804 20946
rect 16960 20602 16988 21830
rect 17052 21622 17080 23054
rect 17040 21616 17092 21622
rect 17040 21558 17092 21564
rect 17040 21344 17092 21350
rect 17040 21286 17092 21292
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 17052 20534 17080 21286
rect 17144 21010 17172 23462
rect 17224 22228 17276 22234
rect 17224 22170 17276 22176
rect 17236 22098 17264 22170
rect 17224 22092 17276 22098
rect 17224 22034 17276 22040
rect 17236 21690 17264 22034
rect 17316 21956 17368 21962
rect 17316 21898 17368 21904
rect 17224 21684 17276 21690
rect 17224 21626 17276 21632
rect 17328 21622 17356 21898
rect 17316 21616 17368 21622
rect 17316 21558 17368 21564
rect 17224 21412 17276 21418
rect 17224 21354 17276 21360
rect 17236 21146 17264 21354
rect 17224 21140 17276 21146
rect 17224 21082 17276 21088
rect 17132 21004 17184 21010
rect 17132 20946 17184 20952
rect 17040 20528 17092 20534
rect 17040 20470 17092 20476
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 16488 20392 16540 20398
rect 16488 20334 16540 20340
rect 16396 20256 16448 20262
rect 16396 20198 16448 20204
rect 16500 19718 16528 20334
rect 16488 19712 16540 19718
rect 16488 19654 16540 19660
rect 16304 19440 16356 19446
rect 16304 19382 16356 19388
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 16132 17814 16160 18226
rect 16120 17808 16172 17814
rect 16120 17750 16172 17756
rect 16316 17678 16344 19382
rect 17316 18624 17368 18630
rect 17316 18566 17368 18572
rect 17040 18420 17092 18426
rect 17040 18362 17092 18368
rect 16396 18216 16448 18222
rect 16396 18158 16448 18164
rect 16408 17814 16436 18158
rect 16856 18080 16908 18086
rect 16856 18022 16908 18028
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16396 17808 16448 17814
rect 16396 17750 16448 17756
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15752 17672 15804 17678
rect 15752 17614 15804 17620
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 15396 16794 15424 17614
rect 15660 17604 15712 17610
rect 15660 17546 15712 17552
rect 15476 17264 15528 17270
rect 15528 17224 15608 17252
rect 15476 17206 15528 17212
rect 15384 16788 15436 16794
rect 15384 16730 15436 16736
rect 15580 16504 15608 17224
rect 15672 17202 15700 17546
rect 15764 17338 15792 17614
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 15752 17332 15804 17338
rect 15752 17274 15804 17280
rect 15856 17218 15884 17478
rect 15764 17202 15884 17218
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15752 17196 15884 17202
rect 15804 17190 15884 17196
rect 16028 17196 16080 17202
rect 15752 17138 15804 17144
rect 16028 17138 16080 17144
rect 16040 16794 16068 17138
rect 16316 16998 16344 17614
rect 16408 17542 16436 17750
rect 16592 17678 16620 17818
rect 16868 17678 16896 18022
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 16120 16788 16172 16794
rect 16120 16730 16172 16736
rect 16132 16674 16160 16730
rect 16040 16646 16160 16674
rect 16040 16590 16068 16646
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 15660 16516 15712 16522
rect 15580 16476 15660 16504
rect 15660 16458 15712 16464
rect 15200 16040 15252 16046
rect 15200 15982 15252 15988
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 14740 14952 14792 14958
rect 14740 14894 14792 14900
rect 14094 11112 14150 11121
rect 14094 11047 14150 11056
rect 14004 10804 14056 10810
rect 14004 10746 14056 10752
rect 13912 10532 13964 10538
rect 13912 10474 13964 10480
rect 13924 10266 13952 10474
rect 14016 10266 14044 10746
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 14108 10062 14136 10678
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 14200 7546 14228 14894
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 14384 13258 14412 13670
rect 14372 13252 14424 13258
rect 14372 13194 14424 13200
rect 14476 11354 14504 14894
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 14556 14340 14608 14346
rect 14556 14282 14608 14288
rect 14568 13190 14596 14282
rect 14660 13870 14688 14418
rect 14844 14006 14872 14962
rect 15016 14952 15068 14958
rect 15016 14894 15068 14900
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 14936 14618 14964 14758
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14832 14000 14884 14006
rect 14832 13942 14884 13948
rect 14936 13938 14964 14214
rect 15028 13938 15056 14894
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14660 12986 14688 13806
rect 14832 13252 14884 13258
rect 14832 13194 14884 13200
rect 14648 12980 14700 12986
rect 14648 12922 14700 12928
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14568 11150 14596 12786
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14752 11150 14780 11698
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14740 11144 14792 11150
rect 14844 11121 14872 13194
rect 14936 11218 14964 13874
rect 15120 13802 15148 15846
rect 16040 15366 16068 16526
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 16028 15360 16080 15366
rect 16028 15302 16080 15308
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 15304 14618 15332 14894
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15212 13841 15240 14350
rect 15396 13870 15424 14418
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15384 13864 15436 13870
rect 15198 13832 15254 13841
rect 15108 13796 15160 13802
rect 15384 13806 15436 13812
rect 15198 13767 15254 13776
rect 15108 13738 15160 13744
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15304 12850 15332 13670
rect 15292 12844 15344 12850
rect 15476 12844 15528 12850
rect 15292 12786 15344 12792
rect 15396 12804 15476 12832
rect 15200 12776 15252 12782
rect 15198 12744 15200 12753
rect 15252 12744 15254 12753
rect 15198 12679 15254 12688
rect 15396 11642 15424 12804
rect 15476 12786 15528 12792
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15580 12374 15608 12786
rect 15568 12368 15620 12374
rect 15120 11614 15424 11642
rect 15488 12328 15568 12356
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 14740 11086 14792 11092
rect 14830 11112 14886 11121
rect 14830 11047 14886 11056
rect 14936 10810 14964 11154
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 14832 10736 14884 10742
rect 14832 10678 14884 10684
rect 14372 10668 14424 10674
rect 14424 10628 14504 10656
rect 14372 10610 14424 10616
rect 14476 10062 14504 10628
rect 14844 10266 14872 10678
rect 15028 10674 15056 10950
rect 15120 10810 15148 11614
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15304 10810 15332 11086
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15396 10742 15424 11154
rect 15488 11082 15516 12328
rect 15568 12310 15620 12316
rect 15566 11792 15622 11801
rect 15566 11727 15568 11736
rect 15620 11727 15622 11736
rect 15568 11698 15620 11704
rect 15566 11520 15622 11529
rect 15566 11455 15622 11464
rect 15580 11150 15608 11455
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15476 11076 15528 11082
rect 15476 11018 15528 11024
rect 15384 10736 15436 10742
rect 15384 10678 15436 10684
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 14936 10062 14964 10610
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15304 10130 15332 10202
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 14476 9722 14504 9998
rect 14464 9716 14516 9722
rect 14740 9716 14792 9722
rect 14464 9658 14516 9664
rect 14660 9664 14740 9674
rect 14660 9658 14792 9664
rect 14660 9654 14780 9658
rect 14648 9648 14780 9654
rect 14700 9646 14780 9648
rect 14648 9590 14700 9596
rect 14464 7948 14516 7954
rect 14464 7890 14516 7896
rect 14280 7812 14332 7818
rect 14280 7754 14332 7760
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14292 7478 14320 7754
rect 14280 7472 14332 7478
rect 14280 7414 14332 7420
rect 13542 7032 13598 7041
rect 14292 7002 14320 7414
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 13542 6967 13598 6976
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 13360 6928 13412 6934
rect 13360 6870 13412 6876
rect 13372 6798 13400 6870
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13452 6792 13504 6798
rect 14096 6792 14148 6798
rect 13452 6734 13504 6740
rect 14016 6740 14096 6746
rect 14016 6734 14148 6740
rect 13372 6662 13400 6734
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13464 6644 13492 6734
rect 13636 6724 13688 6730
rect 13636 6666 13688 6672
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 14016 6718 14136 6734
rect 13544 6656 13596 6662
rect 13464 6616 13544 6644
rect 13464 6497 13492 6616
rect 13648 6633 13676 6666
rect 13544 6598 13596 6604
rect 13634 6624 13690 6633
rect 13634 6559 13690 6568
rect 13450 6488 13506 6497
rect 13450 6423 13506 6432
rect 13832 6186 13860 6666
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 14016 5846 14044 6718
rect 14280 6384 14332 6390
rect 14280 6326 14332 6332
rect 14292 6186 14320 6326
rect 14280 6180 14332 6186
rect 14280 6122 14332 6128
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 14384 5642 14412 7142
rect 14476 6202 14504 7890
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14568 6798 14596 7346
rect 14660 7342 14688 9590
rect 14936 9382 14964 9998
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 15028 9382 15056 9862
rect 15212 9586 15240 9862
rect 15304 9586 15332 10066
rect 15396 10062 15424 10542
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15488 9722 15516 11018
rect 15568 10736 15620 10742
rect 15568 10678 15620 10684
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 15580 9586 15608 10678
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15568 9580 15620 9586
rect 15568 9522 15620 9528
rect 14924 9376 14976 9382
rect 14924 9318 14976 9324
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 14936 8634 14964 9318
rect 15396 9178 15424 9522
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 15200 8356 15252 8362
rect 15200 8298 15252 8304
rect 15212 7886 15240 8298
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14568 6390 14596 6734
rect 14660 6712 14688 7278
rect 14752 6866 14780 7346
rect 14844 6866 14872 7346
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14832 6860 14884 6866
rect 14884 6820 14964 6848
rect 14832 6802 14884 6808
rect 14740 6724 14792 6730
rect 14660 6684 14740 6712
rect 14740 6666 14792 6672
rect 14752 6633 14780 6666
rect 14936 6644 14964 6820
rect 14738 6624 14794 6633
rect 14738 6559 14794 6568
rect 14844 6616 14964 6644
rect 14844 6458 14872 6616
rect 15028 6474 15056 7686
rect 15396 7478 15424 8026
rect 15672 7886 15700 14010
rect 16118 13968 16174 13977
rect 16118 13903 16174 13912
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 15948 13462 15976 13806
rect 16132 13802 16160 13903
rect 16120 13796 16172 13802
rect 16120 13738 16172 13744
rect 15936 13456 15988 13462
rect 15936 13398 15988 13404
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 15764 12850 15792 13126
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15764 10266 15792 12786
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 15844 11756 15896 11762
rect 15844 11698 15896 11704
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15856 11665 15884 11698
rect 15842 11656 15898 11665
rect 15842 11591 15898 11600
rect 15948 10810 15976 11698
rect 16040 11150 16068 12174
rect 16132 12073 16160 13126
rect 16224 12442 16252 13262
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16316 12918 16344 13126
rect 16304 12912 16356 12918
rect 16304 12854 16356 12860
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 16118 12064 16174 12073
rect 16118 11999 16174 12008
rect 16224 11898 16252 12378
rect 16592 12374 16620 15438
rect 16684 15337 16712 15846
rect 16868 15706 16896 17138
rect 17052 16590 17080 18362
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 16948 15972 17000 15978
rect 16948 15914 17000 15920
rect 16856 15700 16908 15706
rect 16856 15642 16908 15648
rect 16960 15638 16988 15914
rect 16948 15632 17000 15638
rect 16948 15574 17000 15580
rect 17052 15570 17080 16526
rect 17144 16250 17172 17138
rect 17132 16244 17184 16250
rect 17132 16186 17184 16192
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17236 16114 17264 16186
rect 17224 16108 17276 16114
rect 17224 16050 17276 16056
rect 17132 15972 17184 15978
rect 17132 15914 17184 15920
rect 17040 15564 17092 15570
rect 17040 15506 17092 15512
rect 16764 15496 16816 15502
rect 16816 15456 16988 15484
rect 16764 15438 16816 15444
rect 16764 15360 16816 15366
rect 16670 15328 16726 15337
rect 16764 15302 16816 15308
rect 16670 15263 16726 15272
rect 16776 15162 16804 15302
rect 16960 15162 16988 15456
rect 16764 15156 16816 15162
rect 16948 15156 17000 15162
rect 16764 15098 16816 15104
rect 16868 15116 16948 15144
rect 16868 14550 16896 15116
rect 16948 15098 17000 15104
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16856 14544 16908 14550
rect 16856 14486 16908 14492
rect 16868 14414 16896 14486
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16488 12368 16540 12374
rect 16488 12310 16540 12316
rect 16580 12368 16632 12374
rect 16580 12310 16632 12316
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16316 11898 16344 12174
rect 16394 12064 16450 12073
rect 16394 11999 16450 12008
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 16210 11656 16266 11665
rect 16120 11620 16172 11626
rect 16210 11591 16266 11600
rect 16120 11562 16172 11568
rect 16132 11529 16160 11562
rect 16118 11520 16174 11529
rect 16118 11455 16174 11464
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 15936 10804 15988 10810
rect 15936 10746 15988 10752
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15750 10024 15806 10033
rect 15750 9959 15806 9968
rect 15764 9382 15792 9959
rect 15856 9654 15884 10610
rect 16040 9897 16068 11086
rect 16120 11008 16172 11014
rect 16120 10950 16172 10956
rect 16132 10674 16160 10950
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16224 10266 16252 11591
rect 16316 11082 16344 11834
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16026 9888 16082 9897
rect 16026 9823 16082 9832
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15568 7880 15620 7886
rect 15568 7822 15620 7828
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 15580 7546 15608 7822
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15384 7472 15436 7478
rect 15384 7414 15436 7420
rect 15764 7342 15792 9318
rect 15842 8120 15898 8129
rect 15842 8055 15844 8064
rect 15896 8055 15898 8064
rect 15844 8026 15896 8032
rect 16132 7478 16160 9522
rect 16120 7472 16172 7478
rect 16120 7414 16172 7420
rect 15752 7336 15804 7342
rect 15752 7278 15804 7284
rect 15658 7032 15714 7041
rect 15658 6967 15714 6976
rect 15672 6798 15700 6967
rect 16224 6934 16252 10202
rect 16212 6928 16264 6934
rect 16212 6870 16264 6876
rect 15660 6792 15712 6798
rect 15106 6760 15162 6769
rect 15660 6734 15712 6740
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15106 6695 15162 6704
rect 15120 6662 15148 6695
rect 15108 6656 15160 6662
rect 15108 6598 15160 6604
rect 14832 6452 14884 6458
rect 15028 6446 15148 6474
rect 15764 6458 15792 6734
rect 14832 6394 14884 6400
rect 14556 6384 14608 6390
rect 14556 6326 14608 6332
rect 15120 6322 15148 6446
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 14556 6248 14608 6254
rect 14476 6196 14556 6202
rect 14476 6190 14608 6196
rect 14476 6174 14596 6190
rect 14648 6112 14700 6118
rect 14646 6080 14648 6089
rect 14700 6080 14702 6089
rect 14646 6015 14702 6024
rect 15396 5914 15424 6258
rect 15856 6186 15884 6734
rect 16408 6322 16436 11999
rect 16500 11626 16528 12310
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16592 11762 16620 12038
rect 16684 11762 16712 13330
rect 16960 13326 16988 14758
rect 17052 14618 17080 14962
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 17144 14498 17172 15914
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 17052 14482 17172 14498
rect 17040 14476 17172 14482
rect 17092 14470 17172 14476
rect 17040 14418 17092 14424
rect 17236 14414 17264 15846
rect 17328 14822 17356 18566
rect 17420 17746 17448 23530
rect 17960 23520 18012 23526
rect 17960 23462 18012 23468
rect 17592 21548 17644 21554
rect 17592 21490 17644 21496
rect 17604 21010 17632 21490
rect 17592 21004 17644 21010
rect 17592 20946 17644 20952
rect 17776 20936 17828 20942
rect 17828 20896 17908 20924
rect 17776 20878 17828 20884
rect 17880 20346 17908 20896
rect 17972 20466 18000 23462
rect 18064 23322 18092 23666
rect 18248 23594 18276 23802
rect 18236 23588 18288 23594
rect 18236 23530 18288 23536
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 18248 23254 18276 23530
rect 18328 23520 18380 23526
rect 18328 23462 18380 23468
rect 18236 23248 18288 23254
rect 18236 23190 18288 23196
rect 18236 22432 18288 22438
rect 18236 22374 18288 22380
rect 18144 21548 18196 21554
rect 18144 21490 18196 21496
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 18064 20942 18092 21422
rect 18052 20936 18104 20942
rect 18052 20878 18104 20884
rect 18156 20874 18184 21490
rect 18144 20868 18196 20874
rect 18144 20810 18196 20816
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 17880 20318 18092 20346
rect 17500 20256 17552 20262
rect 17500 20198 17552 20204
rect 17512 17746 17540 20198
rect 17960 19916 18012 19922
rect 17960 19858 18012 19864
rect 17684 18216 17736 18222
rect 17684 18158 17736 18164
rect 17592 18148 17644 18154
rect 17592 18090 17644 18096
rect 17408 17740 17460 17746
rect 17408 17682 17460 17688
rect 17500 17740 17552 17746
rect 17500 17682 17552 17688
rect 17604 17678 17632 18090
rect 17696 17678 17724 18158
rect 17972 17746 18000 19858
rect 18064 19378 18092 20318
rect 18052 19372 18104 19378
rect 18052 19314 18104 19320
rect 18064 17882 18092 19314
rect 18248 18884 18276 22374
rect 18340 21554 18368 23462
rect 18420 22976 18472 22982
rect 18420 22918 18472 22924
rect 18432 22778 18460 22918
rect 18420 22772 18472 22778
rect 18420 22714 18472 22720
rect 18418 22536 18474 22545
rect 18418 22471 18474 22480
rect 18432 22438 18460 22471
rect 18420 22432 18472 22438
rect 18420 22374 18472 22380
rect 18328 21548 18380 21554
rect 18328 21490 18380 21496
rect 18420 21548 18472 21554
rect 18420 21490 18472 21496
rect 18328 21140 18380 21146
rect 18328 21082 18380 21088
rect 18340 20806 18368 21082
rect 18432 21010 18460 21490
rect 18420 21004 18472 21010
rect 18420 20946 18472 20952
rect 18328 20800 18380 20806
rect 18328 20742 18380 20748
rect 18420 20800 18472 20806
rect 18420 20742 18472 20748
rect 18156 18856 18276 18884
rect 18156 18766 18184 18856
rect 18144 18760 18196 18766
rect 18144 18702 18196 18708
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 18052 17672 18104 17678
rect 18052 17614 18104 17620
rect 17408 17060 17460 17066
rect 17408 17002 17460 17008
rect 17420 16114 17448 17002
rect 17408 16108 17460 16114
rect 17408 16050 17460 16056
rect 17420 15910 17448 16050
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17132 14272 17184 14278
rect 17132 14214 17184 14220
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 17052 12714 17080 13194
rect 17040 12708 17092 12714
rect 17040 12650 17092 12656
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16868 12306 16896 12582
rect 17052 12434 17080 12650
rect 16960 12406 17080 12434
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16672 11756 16724 11762
rect 16724 11716 16896 11744
rect 16672 11698 16724 11704
rect 16488 11620 16540 11626
rect 16488 11562 16540 11568
rect 16592 11354 16620 11698
rect 16580 11348 16632 11354
rect 16764 11348 16816 11354
rect 16580 11290 16632 11296
rect 16684 11308 16764 11336
rect 16684 10538 16712 11308
rect 16764 11290 16816 11296
rect 16868 11218 16896 11716
rect 16856 11212 16908 11218
rect 16776 11172 16856 11200
rect 16776 10742 16804 11172
rect 16856 11154 16908 11160
rect 16854 11112 16910 11121
rect 16854 11047 16856 11056
rect 16908 11047 16910 11056
rect 16856 11018 16908 11024
rect 16764 10736 16816 10742
rect 16764 10678 16816 10684
rect 16960 10554 16988 12406
rect 17144 12238 17172 14214
rect 17420 13462 17448 14894
rect 17604 14890 17632 17614
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17696 15314 17724 17478
rect 18064 17338 18092 17614
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 17960 17060 18012 17066
rect 17960 17002 18012 17008
rect 17972 16402 18000 17002
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 17788 16374 18000 16402
rect 17788 16046 17816 16374
rect 18064 16250 18092 16934
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 18052 16244 18104 16250
rect 18052 16186 18104 16192
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17696 15286 17816 15314
rect 17788 14958 17816 15286
rect 17776 14952 17828 14958
rect 17776 14894 17828 14900
rect 17592 14884 17644 14890
rect 17592 14826 17644 14832
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17696 13841 17724 14350
rect 17682 13832 17738 13841
rect 17682 13767 17738 13776
rect 17788 13734 17816 14894
rect 17776 13728 17828 13734
rect 17776 13670 17828 13676
rect 17880 13462 17908 16186
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 18064 15094 18092 16050
rect 18052 15088 18104 15094
rect 18052 15030 18104 15036
rect 18156 15026 18184 18158
rect 18248 17746 18276 18856
rect 18340 18698 18368 20742
rect 18432 20602 18460 20742
rect 18420 20596 18472 20602
rect 18420 20538 18472 20544
rect 18524 19972 18552 24210
rect 19064 24064 19116 24070
rect 19064 24006 19116 24012
rect 19076 23730 19104 24006
rect 19168 23798 19196 24822
rect 19892 24812 19944 24818
rect 19892 24754 19944 24760
rect 22008 24812 22060 24818
rect 22008 24754 22060 24760
rect 19156 23792 19208 23798
rect 19156 23734 19208 23740
rect 18604 23724 18656 23730
rect 18604 23666 18656 23672
rect 18788 23724 18840 23730
rect 18788 23666 18840 23672
rect 19064 23724 19116 23730
rect 19064 23666 19116 23672
rect 18616 22438 18644 23666
rect 18696 22704 18748 22710
rect 18694 22672 18696 22681
rect 18748 22672 18750 22681
rect 18694 22607 18750 22616
rect 18604 22432 18656 22438
rect 18604 22374 18656 22380
rect 18616 21554 18644 22374
rect 18604 21548 18656 21554
rect 18604 21490 18656 21496
rect 18800 21146 18828 23666
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18892 22778 18920 22918
rect 18880 22772 18932 22778
rect 18880 22714 18932 22720
rect 18970 22672 19026 22681
rect 18880 22636 18932 22642
rect 18970 22607 18972 22616
rect 18880 22578 18932 22584
rect 19024 22607 19026 22616
rect 18972 22578 19024 22584
rect 18892 22506 18920 22578
rect 18880 22500 18932 22506
rect 18880 22442 18932 22448
rect 19076 22098 19104 23666
rect 19064 22092 19116 22098
rect 19064 22034 19116 22040
rect 18880 21616 18932 21622
rect 18880 21558 18932 21564
rect 18788 21140 18840 21146
rect 18788 21082 18840 21088
rect 18788 20936 18840 20942
rect 18788 20878 18840 20884
rect 18696 20868 18748 20874
rect 18696 20810 18748 20816
rect 18604 20460 18656 20466
rect 18604 20402 18656 20408
rect 18432 19944 18552 19972
rect 18432 18766 18460 19944
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18328 18692 18380 18698
rect 18328 18634 18380 18640
rect 18236 17740 18288 17746
rect 18236 17682 18288 17688
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18340 17202 18368 17614
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17408 13456 17460 13462
rect 17408 13398 17460 13404
rect 17868 13456 17920 13462
rect 17868 13398 17920 13404
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17868 13320 17920 13326
rect 17868 13262 17920 13268
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17040 12096 17092 12102
rect 17236 12073 17264 12174
rect 17040 12038 17092 12044
rect 17222 12064 17278 12073
rect 17052 11830 17080 12038
rect 17222 11999 17278 12008
rect 17040 11824 17092 11830
rect 17040 11766 17092 11772
rect 17052 10674 17080 11766
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17224 10736 17276 10742
rect 17224 10678 17276 10684
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 16672 10532 16724 10538
rect 16960 10526 17080 10554
rect 16672 10474 16724 10480
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16500 9722 16528 9998
rect 16488 9716 16540 9722
rect 16684 9704 16712 10474
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16868 10130 16896 10406
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16764 9988 16816 9994
rect 16764 9930 16816 9936
rect 16856 9988 16908 9994
rect 16856 9930 16908 9936
rect 16776 9897 16804 9930
rect 16762 9888 16818 9897
rect 16762 9823 16818 9832
rect 16488 9658 16540 9664
rect 16592 9676 16712 9704
rect 16592 9625 16620 9676
rect 16578 9616 16634 9625
rect 16868 9586 16896 9930
rect 16578 9551 16634 9560
rect 16856 9580 16908 9586
rect 16592 8090 16620 9551
rect 16856 9522 16908 9528
rect 16960 9518 16988 9998
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16856 9444 16908 9450
rect 16856 9386 16908 9392
rect 16868 9330 16896 9386
rect 17052 9330 17080 10526
rect 17132 9920 17184 9926
rect 17132 9862 17184 9868
rect 16868 9302 17080 9330
rect 16868 8906 16896 9302
rect 16856 8900 16908 8906
rect 16856 8842 16908 8848
rect 17144 8634 17172 9862
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17144 8362 17172 8570
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 17040 8288 17092 8294
rect 17040 8230 17092 8236
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 15844 6180 15896 6186
rect 15844 6122 15896 6128
rect 15856 5914 15884 6122
rect 16408 6118 16436 6258
rect 16592 6186 16620 8026
rect 17052 7954 17080 8230
rect 17040 7948 17092 7954
rect 17040 7890 17092 7896
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16776 6866 16804 7278
rect 16764 6860 16816 6866
rect 16764 6802 16816 6808
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16684 6662 16712 6734
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16580 6180 16632 6186
rect 16580 6122 16632 6128
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 16776 5642 16804 6802
rect 17040 6792 17092 6798
rect 17038 6760 17040 6769
rect 17092 6760 17094 6769
rect 17038 6695 17094 6704
rect 17236 6254 17264 10678
rect 17328 10538 17356 11494
rect 17316 10532 17368 10538
rect 17316 10474 17368 10480
rect 17328 10062 17356 10474
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17420 7886 17448 8230
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17316 7744 17368 7750
rect 17316 7686 17368 7692
rect 17328 6798 17356 7686
rect 17512 7546 17540 13262
rect 17880 12782 17908 13262
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17776 11824 17828 11830
rect 17776 11766 17828 11772
rect 17788 11121 17816 11766
rect 17774 11112 17830 11121
rect 17774 11047 17830 11056
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17604 8498 17632 9454
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17512 6458 17540 7482
rect 17604 7410 17632 8434
rect 17696 7818 17724 9998
rect 17788 9674 17816 11047
rect 17972 10062 18000 14418
rect 18144 14340 18196 14346
rect 18144 14282 18196 14288
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 18064 12850 18092 13330
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 18064 12374 18092 12786
rect 18052 12368 18104 12374
rect 18052 12310 18104 12316
rect 18052 12232 18104 12238
rect 18050 12200 18052 12209
rect 18104 12200 18106 12209
rect 18050 12135 18106 12144
rect 18064 11286 18092 12135
rect 18052 11280 18104 11286
rect 18052 11222 18104 11228
rect 18052 11144 18104 11150
rect 18050 11112 18052 11121
rect 18104 11112 18106 11121
rect 18050 11047 18106 11056
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 17972 9722 18000 9998
rect 18064 9994 18092 10406
rect 18156 10266 18184 14282
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18328 13932 18380 13938
rect 18432 13920 18460 18702
rect 18512 18692 18564 18698
rect 18512 18634 18564 18640
rect 18524 13938 18552 18634
rect 18616 14618 18644 20402
rect 18708 19378 18736 20810
rect 18800 20806 18828 20878
rect 18788 20800 18840 20806
rect 18788 20742 18840 20748
rect 18800 19514 18828 20742
rect 18892 20602 18920 21558
rect 19076 21554 19104 22034
rect 19064 21548 19116 21554
rect 19064 21490 19116 21496
rect 19064 21140 19116 21146
rect 19064 21082 19116 21088
rect 19076 20942 19104 21082
rect 19168 20942 19196 23734
rect 19904 23662 19932 24754
rect 21456 24676 21508 24682
rect 21456 24618 21508 24624
rect 21364 24608 21416 24614
rect 21364 24550 21416 24556
rect 21272 24200 21324 24206
rect 21270 24168 21272 24177
rect 21324 24168 21326 24177
rect 20352 24132 20404 24138
rect 20352 24074 20404 24080
rect 20536 24132 20588 24138
rect 21270 24103 21326 24112
rect 20536 24074 20588 24080
rect 20364 23798 20392 24074
rect 20548 23866 20576 24074
rect 20536 23860 20588 23866
rect 20536 23802 20588 23808
rect 21376 23798 21404 24550
rect 21468 24206 21496 24618
rect 22020 24410 22048 24754
rect 22192 24608 22244 24614
rect 22192 24550 22244 24556
rect 22008 24404 22060 24410
rect 22008 24346 22060 24352
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 21548 24200 21600 24206
rect 21548 24142 21600 24148
rect 21560 23866 21588 24142
rect 22204 24070 22232 24550
rect 22008 24064 22060 24070
rect 22008 24006 22060 24012
rect 22192 24064 22244 24070
rect 22192 24006 22244 24012
rect 22296 24018 22324 26250
rect 22480 25974 22508 26318
rect 22468 25968 22520 25974
rect 22468 25910 22520 25916
rect 22664 25906 22692 26318
rect 23124 26314 23152 26726
rect 23308 26450 23336 27066
rect 23400 26790 23428 27338
rect 24044 26858 24072 27406
rect 24308 27396 24360 27402
rect 24228 27356 24308 27384
rect 24228 26994 24256 27356
rect 24308 27338 24360 27344
rect 24504 27062 24532 27406
rect 24492 27056 24544 27062
rect 24492 26998 24544 27004
rect 24216 26988 24268 26994
rect 24216 26930 24268 26936
rect 24400 26988 24452 26994
rect 24400 26930 24452 26936
rect 24032 26852 24084 26858
rect 24032 26794 24084 26800
rect 23388 26784 23440 26790
rect 23388 26726 23440 26732
rect 23296 26444 23348 26450
rect 23296 26386 23348 26392
rect 23112 26308 23164 26314
rect 23112 26250 23164 26256
rect 23400 25974 23428 26726
rect 23572 26512 23624 26518
rect 23572 26454 23624 26460
rect 23584 26353 23612 26454
rect 23570 26344 23626 26353
rect 23570 26279 23626 26288
rect 23020 25968 23072 25974
rect 23020 25910 23072 25916
rect 23388 25968 23440 25974
rect 23388 25910 23440 25916
rect 22652 25900 22704 25906
rect 22652 25842 22704 25848
rect 22376 24608 22428 24614
rect 22376 24550 22428 24556
rect 22388 24274 22416 24550
rect 22376 24268 22428 24274
rect 22376 24210 22428 24216
rect 21548 23860 21600 23866
rect 21548 23802 21600 23808
rect 20352 23792 20404 23798
rect 20352 23734 20404 23740
rect 21364 23792 21416 23798
rect 21364 23734 21416 23740
rect 19892 23656 19944 23662
rect 21560 23644 21588 23802
rect 22020 23798 22048 24006
rect 22204 23882 22232 24006
rect 22296 23990 22416 24018
rect 22204 23854 22324 23882
rect 22008 23792 22060 23798
rect 22008 23734 22060 23740
rect 21640 23656 21692 23662
rect 21560 23616 21640 23644
rect 19892 23598 19944 23604
rect 21640 23598 21692 23604
rect 21916 23520 21968 23526
rect 21916 23462 21968 23468
rect 21928 23118 21956 23462
rect 22296 23322 22324 23854
rect 22284 23316 22336 23322
rect 22284 23258 22336 23264
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 19432 23112 19484 23118
rect 19432 23054 19484 23060
rect 21180 23112 21232 23118
rect 21180 23054 21232 23060
rect 21916 23112 21968 23118
rect 21916 23054 21968 23060
rect 19340 22976 19392 22982
rect 19340 22918 19392 22924
rect 19352 22760 19380 22918
rect 19260 22732 19380 22760
rect 19260 22545 19288 22732
rect 19246 22536 19302 22545
rect 19246 22471 19302 22480
rect 19352 22438 19380 22732
rect 19444 22506 19472 23054
rect 19524 22636 19576 22642
rect 19524 22578 19576 22584
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 19432 22500 19484 22506
rect 19432 22442 19484 22448
rect 19340 22432 19392 22438
rect 19340 22374 19392 22380
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19444 21486 19472 21830
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19064 20936 19116 20942
rect 19064 20878 19116 20884
rect 19156 20936 19208 20942
rect 19208 20896 19288 20924
rect 19156 20878 19208 20884
rect 19260 20788 19288 20896
rect 19260 20760 19380 20788
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 18708 18766 18736 19110
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18708 17678 18736 18702
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18892 17524 18920 20538
rect 19352 20466 19380 20760
rect 18972 20460 19024 20466
rect 18972 20402 19024 20408
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 18984 20262 19012 20402
rect 19260 20346 19288 20402
rect 19260 20318 19380 20346
rect 18972 20256 19024 20262
rect 18972 20198 19024 20204
rect 18984 19990 19012 20198
rect 19352 20058 19380 20318
rect 19444 20058 19472 21422
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 18972 19984 19024 19990
rect 18972 19926 19024 19932
rect 19444 19496 19472 19994
rect 19352 19468 19472 19496
rect 19352 19394 19380 19468
rect 19536 19446 19564 22578
rect 20732 22098 20760 22578
rect 21192 22574 21220 23054
rect 22008 23044 22060 23050
rect 22008 22986 22060 22992
rect 22020 22710 22048 22986
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 22008 22704 22060 22710
rect 22008 22646 22060 22652
rect 21180 22568 21232 22574
rect 21180 22510 21232 22516
rect 22112 22522 22140 22918
rect 22296 22778 22324 23122
rect 22284 22772 22336 22778
rect 22284 22714 22336 22720
rect 22388 22710 22416 23990
rect 22560 23656 22612 23662
rect 22560 23598 22612 23604
rect 22376 22704 22428 22710
rect 22376 22646 22428 22652
rect 22388 22522 22416 22646
rect 21192 22234 21220 22510
rect 22112 22494 22416 22522
rect 21180 22228 21232 22234
rect 21180 22170 21232 22176
rect 20720 22092 20772 22098
rect 20720 22034 20772 22040
rect 22192 22024 22244 22030
rect 22192 21966 22244 21972
rect 21088 21956 21140 21962
rect 21088 21898 21140 21904
rect 19616 21616 19668 21622
rect 19616 21558 19668 21564
rect 18984 19378 19380 19394
rect 19524 19440 19576 19446
rect 19524 19382 19576 19388
rect 18972 19372 19380 19378
rect 19024 19366 19380 19372
rect 19432 19372 19484 19378
rect 18972 19314 19024 19320
rect 19432 19314 19484 19320
rect 19444 19258 19472 19314
rect 19536 19310 19564 19382
rect 19352 19230 19472 19258
rect 19524 19304 19576 19310
rect 19524 19246 19576 19252
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 18984 18698 19012 19110
rect 18972 18692 19024 18698
rect 18972 18634 19024 18640
rect 18984 17542 19012 18634
rect 19248 18624 19300 18630
rect 19248 18566 19300 18572
rect 19260 18222 19288 18566
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 19156 17740 19208 17746
rect 19156 17682 19208 17688
rect 18708 17496 18920 17524
rect 18972 17536 19024 17542
rect 18708 17338 18736 17496
rect 18972 17478 19024 17484
rect 18696 17332 18748 17338
rect 18696 17274 18748 17280
rect 18708 15706 18736 17274
rect 19064 17196 19116 17202
rect 19064 17138 19116 17144
rect 18880 16244 18932 16250
rect 18880 16186 18932 16192
rect 18892 16114 18920 16186
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 18696 15700 18748 15706
rect 18696 15642 18748 15648
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18380 13892 18460 13920
rect 18512 13932 18564 13938
rect 18328 13874 18380 13880
rect 18512 13874 18564 13880
rect 18248 13410 18276 13874
rect 18248 13382 18368 13410
rect 18236 12912 18288 12918
rect 18236 12854 18288 12860
rect 18248 12209 18276 12854
rect 18234 12200 18290 12209
rect 18234 12135 18290 12144
rect 18236 12096 18288 12102
rect 18340 12084 18368 13382
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18432 12238 18460 12786
rect 18524 12306 18552 12786
rect 18708 12434 18736 15642
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 18800 12753 18828 14826
rect 19076 14278 19104 17138
rect 19168 16998 19196 17682
rect 19352 17678 19380 19230
rect 19628 19122 19656 21558
rect 19984 21412 20036 21418
rect 19984 21354 20036 21360
rect 19892 21072 19944 21078
rect 19890 21040 19892 21049
rect 19944 21040 19946 21049
rect 19890 20975 19946 20984
rect 19996 20942 20024 21354
rect 20444 21072 20496 21078
rect 20442 21040 20444 21049
rect 20496 21040 20498 21049
rect 20442 20975 20498 20984
rect 19708 20936 19760 20942
rect 19708 20878 19760 20884
rect 19892 20936 19944 20942
rect 19892 20878 19944 20884
rect 19984 20936 20036 20942
rect 19984 20878 20036 20884
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 19720 20330 19748 20878
rect 19800 20800 19852 20806
rect 19800 20742 19852 20748
rect 19812 20534 19840 20742
rect 19800 20528 19852 20534
rect 19800 20470 19852 20476
rect 19904 20380 19932 20878
rect 20088 20534 20116 20878
rect 20076 20528 20128 20534
rect 20076 20470 20128 20476
rect 20536 20528 20588 20534
rect 20536 20470 20588 20476
rect 19812 20352 19932 20380
rect 20548 20369 20576 20470
rect 20996 20392 21048 20398
rect 20534 20360 20590 20369
rect 19708 20324 19760 20330
rect 19708 20266 19760 20272
rect 19720 20058 19748 20266
rect 19708 20052 19760 20058
rect 19708 19994 19760 20000
rect 19812 19825 19840 20352
rect 20996 20334 21048 20340
rect 20534 20295 20590 20304
rect 19798 19816 19854 19825
rect 19798 19751 19854 19760
rect 19812 19718 19840 19751
rect 19800 19712 19852 19718
rect 19800 19654 19852 19660
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19800 19372 19852 19378
rect 19800 19314 19852 19320
rect 19444 19094 19656 19122
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 19340 17536 19392 17542
rect 19340 17478 19392 17484
rect 19352 17202 19380 17478
rect 19340 17196 19392 17202
rect 19340 17138 19392 17144
rect 19156 16992 19208 16998
rect 19156 16934 19208 16940
rect 19340 15972 19392 15978
rect 19340 15914 19392 15920
rect 19248 14544 19300 14550
rect 19248 14486 19300 14492
rect 19064 14272 19116 14278
rect 19064 14214 19116 14220
rect 18880 13796 18932 13802
rect 18880 13738 18932 13744
rect 18786 12744 18842 12753
rect 18892 12714 18920 13738
rect 18786 12679 18842 12688
rect 18880 12708 18932 12714
rect 18800 12442 18828 12679
rect 18880 12650 18932 12656
rect 18616 12406 18736 12434
rect 18788 12436 18840 12442
rect 18512 12300 18564 12306
rect 18512 12242 18564 12248
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 18510 12200 18566 12209
rect 18510 12135 18566 12144
rect 18288 12056 18368 12084
rect 18236 12038 18288 12044
rect 18248 11694 18276 12038
rect 18236 11688 18288 11694
rect 18236 11630 18288 11636
rect 18328 11620 18380 11626
rect 18328 11562 18380 11568
rect 18340 11354 18368 11562
rect 18524 11393 18552 12135
rect 18510 11384 18566 11393
rect 18328 11348 18380 11354
rect 18510 11319 18566 11328
rect 18328 11290 18380 11296
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 18432 10062 18460 10950
rect 18512 10668 18564 10674
rect 18512 10610 18564 10616
rect 18524 10130 18552 10610
rect 18616 10198 18644 12406
rect 19076 12434 19104 14214
rect 19156 12776 19208 12782
rect 19156 12718 19208 12724
rect 19168 12646 19196 12718
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 18788 12378 18840 12384
rect 18984 12406 19104 12434
rect 18788 12232 18840 12238
rect 18788 12174 18840 12180
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18708 11762 18736 12038
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18708 11150 18736 11698
rect 18800 11558 18828 12174
rect 18880 11756 18932 11762
rect 18880 11698 18932 11704
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18892 10810 18920 11698
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 18788 10600 18840 10606
rect 18788 10542 18840 10548
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 18604 10192 18656 10198
rect 18604 10134 18656 10140
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 18052 9988 18104 9994
rect 18052 9930 18104 9936
rect 17960 9716 18012 9722
rect 17788 9646 17908 9674
rect 17960 9658 18012 9664
rect 17776 8900 17828 8906
rect 17776 8842 17828 8848
rect 17788 8430 17816 8842
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17880 8106 17908 9646
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 18248 9042 18276 9454
rect 18236 9036 18288 9042
rect 18236 8978 18288 8984
rect 18340 8634 18368 9454
rect 18708 9178 18736 10542
rect 18800 10266 18828 10542
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 18892 9722 18920 10542
rect 18984 10470 19012 12406
rect 19156 12368 19208 12374
rect 19156 12310 19208 12316
rect 19168 12238 19196 12310
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 19076 11762 19104 12038
rect 19064 11756 19116 11762
rect 19064 11698 19116 11704
rect 19076 11218 19104 11698
rect 19260 11354 19288 14486
rect 19352 14346 19380 15914
rect 19444 14550 19472 19094
rect 19708 18692 19760 18698
rect 19708 18634 19760 18640
rect 19720 18086 19748 18634
rect 19708 18080 19760 18086
rect 19708 18022 19760 18028
rect 19524 16516 19576 16522
rect 19524 16458 19576 16464
rect 19536 15434 19564 16458
rect 19616 16244 19668 16250
rect 19616 16186 19668 16192
rect 19628 15638 19656 16186
rect 19616 15632 19668 15638
rect 19616 15574 19668 15580
rect 19524 15428 19576 15434
rect 19524 15370 19576 15376
rect 19720 14822 19748 18022
rect 19812 17814 19840 19314
rect 19800 17808 19852 17814
rect 19800 17750 19852 17756
rect 19904 17202 19932 19654
rect 20444 19372 20496 19378
rect 20548 19360 20576 20295
rect 20628 20256 20680 20262
rect 20626 20224 20628 20233
rect 20904 20256 20956 20262
rect 20680 20224 20682 20233
rect 20904 20198 20956 20204
rect 20626 20159 20682 20168
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20496 19332 20576 19360
rect 20444 19314 20496 19320
rect 20640 18358 20668 19994
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20732 19378 20760 19790
rect 20812 19780 20864 19786
rect 20812 19722 20864 19728
rect 20824 19514 20852 19722
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20824 19378 20852 19450
rect 20916 19417 20944 20198
rect 21008 19802 21036 20334
rect 21100 20262 21128 21898
rect 21456 21140 21508 21146
rect 21456 21082 21508 21088
rect 21468 20942 21496 21082
rect 22204 21078 22232 21966
rect 22192 21072 22244 21078
rect 22192 21014 22244 21020
rect 21548 21004 21600 21010
rect 21600 20964 21772 20992
rect 21548 20946 21600 20952
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21744 20924 21772 20964
rect 21824 20936 21876 20942
rect 21744 20896 21824 20924
rect 21548 20868 21600 20874
rect 21548 20810 21600 20816
rect 21560 20466 21588 20810
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 21548 20460 21600 20466
rect 21548 20402 21600 20408
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 21100 19922 21128 20198
rect 21192 20058 21220 20402
rect 21376 20369 21404 20402
rect 21456 20392 21508 20398
rect 21362 20360 21418 20369
rect 21456 20334 21508 20340
rect 21362 20295 21418 20304
rect 21180 20052 21232 20058
rect 21180 19994 21232 20000
rect 21468 19922 21496 20334
rect 21088 19916 21140 19922
rect 21088 19858 21140 19864
rect 21456 19916 21508 19922
rect 21456 19858 21508 19864
rect 21364 19848 21416 19854
rect 21008 19796 21364 19802
rect 21008 19790 21416 19796
rect 21008 19774 21404 19790
rect 21560 19786 21588 20402
rect 21638 20224 21694 20233
rect 21638 20159 21694 20168
rect 21652 19786 21680 20159
rect 20902 19408 20958 19417
rect 20720 19372 20772 19378
rect 20720 19314 20772 19320
rect 20812 19372 20864 19378
rect 20902 19343 20958 19352
rect 20812 19314 20864 19320
rect 20732 18426 20760 19314
rect 21376 18426 21404 19774
rect 21548 19780 21600 19786
rect 21548 19722 21600 19728
rect 21640 19780 21692 19786
rect 21640 19722 21692 19728
rect 21744 19666 21772 20896
rect 21824 20878 21876 20884
rect 21916 20800 21968 20806
rect 21916 20742 21968 20748
rect 22100 20800 22152 20806
rect 22100 20742 22152 20748
rect 21824 20392 21876 20398
rect 21824 20334 21876 20340
rect 21468 19638 21772 19666
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 20628 18352 20680 18358
rect 20628 18294 20680 18300
rect 20352 18284 20404 18290
rect 20352 18226 20404 18232
rect 19892 17196 19944 17202
rect 19892 17138 19944 17144
rect 19800 17128 19852 17134
rect 19800 17070 19852 17076
rect 20168 17128 20220 17134
rect 20168 17070 20220 17076
rect 19812 16454 19840 17070
rect 20180 16658 20208 17070
rect 20168 16652 20220 16658
rect 20168 16594 20220 16600
rect 20168 16516 20220 16522
rect 20168 16458 20220 16464
rect 19800 16448 19852 16454
rect 19800 16390 19852 16396
rect 19984 16448 20036 16454
rect 19984 16390 20036 16396
rect 19892 16176 19944 16182
rect 19892 16118 19944 16124
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19708 14816 19760 14822
rect 19708 14758 19760 14764
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19352 13394 19380 14282
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19352 12714 19380 13194
rect 19340 12708 19392 12714
rect 19340 12650 19392 12656
rect 19352 12442 19380 12650
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19338 12336 19394 12345
rect 19338 12271 19340 12280
rect 19392 12271 19394 12280
rect 19340 12242 19392 12248
rect 19444 11898 19472 14350
rect 19616 13932 19668 13938
rect 19616 13874 19668 13880
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19536 11898 19564 12718
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 19536 11762 19564 11834
rect 19524 11756 19576 11762
rect 19524 11698 19576 11704
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19064 11212 19116 11218
rect 19064 11154 19116 11160
rect 19260 10674 19288 11290
rect 19628 10674 19656 13874
rect 19720 11762 19748 14758
rect 19812 14414 19840 15302
rect 19800 14408 19852 14414
rect 19800 14350 19852 14356
rect 19800 12776 19852 12782
rect 19800 12718 19852 12724
rect 19812 12170 19840 12718
rect 19904 12442 19932 16118
rect 19996 15502 20024 16390
rect 20180 16250 20208 16458
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 20272 15570 20300 15846
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 20272 15026 20300 15506
rect 20364 15434 20392 18226
rect 20996 17808 21048 17814
rect 20996 17750 21048 17756
rect 21008 17678 21036 17750
rect 20720 17672 20772 17678
rect 20640 17632 20720 17660
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20456 16046 20484 16526
rect 20444 16040 20496 16046
rect 20444 15982 20496 15988
rect 20352 15428 20404 15434
rect 20352 15370 20404 15376
rect 20640 15094 20668 17632
rect 20720 17614 20772 17620
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 20916 17338 20944 17614
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 20904 17332 20956 17338
rect 20904 17274 20956 17280
rect 20824 16794 20852 17274
rect 20996 17264 21048 17270
rect 20996 17206 21048 17212
rect 21008 16998 21036 17206
rect 21284 17202 21312 17614
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20812 16788 20864 16794
rect 20812 16730 20864 16736
rect 20732 16561 20760 16730
rect 20916 16658 20944 16934
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 21088 16652 21140 16658
rect 21468 16640 21496 19638
rect 21638 19544 21694 19553
rect 21638 19479 21640 19488
rect 21692 19479 21694 19488
rect 21640 19450 21692 19456
rect 21732 19440 21784 19446
rect 21732 19382 21784 19388
rect 21640 19168 21692 19174
rect 21640 19110 21692 19116
rect 21088 16594 21140 16600
rect 21376 16612 21496 16640
rect 20718 16552 20774 16561
rect 20718 16487 20774 16496
rect 20732 15570 20760 16487
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 20916 16114 20944 16390
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20824 15162 20852 15438
rect 20812 15156 20864 15162
rect 21008 15144 21036 16390
rect 21100 16046 21128 16594
rect 21088 16040 21140 16046
rect 21088 15982 21140 15988
rect 21088 15360 21140 15366
rect 21088 15302 21140 15308
rect 20812 15098 20864 15104
rect 20916 15116 21036 15144
rect 20628 15088 20680 15094
rect 20680 15036 20760 15042
rect 20628 15030 20760 15036
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 20260 15020 20312 15026
rect 20640 15014 20760 15030
rect 20916 15026 20944 15116
rect 21100 15026 21128 15302
rect 20260 14962 20312 14968
rect 19996 13841 20024 14962
rect 20732 14958 20760 15014
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 21088 15020 21140 15026
rect 21088 14962 21140 14968
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 20076 14816 20128 14822
rect 20076 14758 20128 14764
rect 20088 14482 20116 14758
rect 20640 14550 20668 14894
rect 20628 14544 20680 14550
rect 20628 14486 20680 14492
rect 20076 14476 20128 14482
rect 20076 14418 20128 14424
rect 20904 14476 20956 14482
rect 20904 14418 20956 14424
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 19982 13832 20038 13841
rect 19982 13767 20038 13776
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19996 13297 20024 13330
rect 19982 13288 20038 13297
rect 19982 13223 20038 13232
rect 20076 13184 20128 13190
rect 20076 13126 20128 13132
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20088 12918 20116 13126
rect 20076 12912 20128 12918
rect 20076 12854 20128 12860
rect 19892 12436 19944 12442
rect 19892 12378 19944 12384
rect 20088 12322 20116 12854
rect 19904 12306 20116 12322
rect 19892 12300 20116 12306
rect 19944 12294 20116 12300
rect 19892 12242 19944 12248
rect 19800 12164 19852 12170
rect 19800 12106 19852 12112
rect 20088 12050 20116 12294
rect 20272 12238 20300 13126
rect 20628 12980 20680 12986
rect 20628 12922 20680 12928
rect 20534 12336 20590 12345
rect 20534 12271 20536 12280
rect 20588 12271 20590 12280
rect 20536 12242 20588 12248
rect 20640 12238 20668 12922
rect 20824 12782 20852 14010
rect 20916 13802 20944 14418
rect 21008 14414 21036 14962
rect 21180 14884 21232 14890
rect 21180 14826 21232 14832
rect 21192 14482 21220 14826
rect 21376 14618 21404 16612
rect 21652 16590 21680 19110
rect 21744 17202 21772 19382
rect 21836 18834 21864 20334
rect 21824 18828 21876 18834
rect 21824 18770 21876 18776
rect 21928 17762 21956 20742
rect 22112 20534 22140 20742
rect 22100 20528 22152 20534
rect 22100 20470 22152 20476
rect 22204 20380 22232 21014
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22468 20936 22520 20942
rect 22468 20878 22520 20884
rect 22388 20602 22416 20878
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 22112 20352 22232 20380
rect 22112 19854 22140 20352
rect 22388 20074 22416 20538
rect 22296 20046 22416 20074
rect 22296 19990 22324 20046
rect 22284 19984 22336 19990
rect 22284 19926 22336 19932
rect 22192 19916 22244 19922
rect 22192 19858 22244 19864
rect 22008 19848 22060 19854
rect 22008 19790 22060 19796
rect 22100 19848 22152 19854
rect 22100 19790 22152 19796
rect 22020 19718 22048 19790
rect 22008 19712 22060 19718
rect 22100 19712 22152 19718
rect 22060 19672 22100 19700
rect 22008 19654 22060 19660
rect 22100 19654 22152 19660
rect 22204 19334 22232 19858
rect 22376 19848 22428 19854
rect 22374 19816 22376 19825
rect 22428 19816 22430 19825
rect 22284 19780 22336 19786
rect 22374 19751 22430 19760
rect 22284 19722 22336 19728
rect 22112 19306 22232 19334
rect 22008 18284 22060 18290
rect 22112 18272 22140 19306
rect 22296 19242 22324 19722
rect 22376 19440 22428 19446
rect 22480 19428 22508 20878
rect 22572 20534 22600 23598
rect 22664 23050 22692 25842
rect 23032 25498 23060 25910
rect 24228 25906 24256 26930
rect 24308 26784 24360 26790
rect 24306 26752 24308 26761
rect 24360 26752 24362 26761
rect 24306 26687 24362 26696
rect 24320 26382 24348 26687
rect 24308 26376 24360 26382
rect 24308 26318 24360 26324
rect 24412 26314 24440 26930
rect 24492 26920 24544 26926
rect 24492 26862 24544 26868
rect 24504 26314 24532 26862
rect 24596 26790 24624 27610
rect 24688 26994 24716 28036
rect 24768 28018 24820 28024
rect 24860 27872 24912 27878
rect 24860 27814 24912 27820
rect 24872 27690 24900 27814
rect 24780 27662 24900 27690
rect 24952 27668 25004 27674
rect 24780 27470 24808 27662
rect 24952 27610 25004 27616
rect 24860 27532 24912 27538
rect 24860 27474 24912 27480
rect 24768 27464 24820 27470
rect 24768 27406 24820 27412
rect 24872 27130 24900 27474
rect 24964 27452 24992 27610
rect 25056 27606 25084 28426
rect 25228 28008 25280 28014
rect 25228 27950 25280 27956
rect 25136 27940 25188 27946
rect 25136 27882 25188 27888
rect 25148 27674 25176 27882
rect 25136 27668 25188 27674
rect 25136 27610 25188 27616
rect 25044 27600 25096 27606
rect 25044 27542 25096 27548
rect 25044 27464 25096 27470
rect 24964 27424 25044 27452
rect 25044 27406 25096 27412
rect 24952 27328 25004 27334
rect 24952 27270 25004 27276
rect 25136 27328 25188 27334
rect 25136 27270 25188 27276
rect 24860 27124 24912 27130
rect 24860 27066 24912 27072
rect 24964 26994 24992 27270
rect 24676 26988 24728 26994
rect 24676 26930 24728 26936
rect 24952 26988 25004 26994
rect 24952 26930 25004 26936
rect 24688 26790 24716 26930
rect 24584 26784 24636 26790
rect 24584 26726 24636 26732
rect 24676 26784 24728 26790
rect 24676 26726 24728 26732
rect 24676 26580 24728 26586
rect 24676 26522 24728 26528
rect 24400 26308 24452 26314
rect 24400 26250 24452 26256
rect 24492 26308 24544 26314
rect 24492 26250 24544 26256
rect 24216 25900 24268 25906
rect 24216 25842 24268 25848
rect 23020 25492 23072 25498
rect 23020 25434 23072 25440
rect 23756 24880 23808 24886
rect 23756 24822 23808 24828
rect 22928 24812 22980 24818
rect 22928 24754 22980 24760
rect 23112 24812 23164 24818
rect 23112 24754 23164 24760
rect 22940 24177 22968 24754
rect 23124 24410 23152 24754
rect 23480 24608 23532 24614
rect 23480 24550 23532 24556
rect 23492 24410 23520 24550
rect 23112 24404 23164 24410
rect 23112 24346 23164 24352
rect 23480 24404 23532 24410
rect 23480 24346 23532 24352
rect 23768 24206 23796 24822
rect 24688 24342 24716 26522
rect 25044 26444 25096 26450
rect 25044 26386 25096 26392
rect 25056 25906 25084 26386
rect 25148 26382 25176 27270
rect 25136 26376 25188 26382
rect 25136 26318 25188 26324
rect 25240 26314 25268 27950
rect 25320 27872 25372 27878
rect 25320 27814 25372 27820
rect 25332 26994 25360 27814
rect 25504 27668 25556 27674
rect 25504 27610 25556 27616
rect 25412 27464 25464 27470
rect 25412 27406 25464 27412
rect 25320 26988 25372 26994
rect 25320 26930 25372 26936
rect 25424 26450 25452 27406
rect 25516 26926 25544 27610
rect 25608 27130 25636 28426
rect 25780 28076 25832 28082
rect 25780 28018 25832 28024
rect 25596 27124 25648 27130
rect 25596 27066 25648 27072
rect 25792 26994 25820 28018
rect 25872 27396 25924 27402
rect 25872 27338 25924 27344
rect 25884 27130 25912 27338
rect 25964 27328 26016 27334
rect 25964 27270 26016 27276
rect 25872 27124 25924 27130
rect 25872 27066 25924 27072
rect 25976 26994 26004 27270
rect 26068 27130 26096 28494
rect 26424 28484 26476 28490
rect 26424 28426 26476 28432
rect 26332 28076 26384 28082
rect 26332 28018 26384 28024
rect 26148 27940 26200 27946
rect 26148 27882 26200 27888
rect 26160 27538 26188 27882
rect 26148 27532 26200 27538
rect 26148 27474 26200 27480
rect 26240 27464 26292 27470
rect 26240 27406 26292 27412
rect 26252 27130 26280 27406
rect 26344 27130 26372 28018
rect 26436 27674 26464 28426
rect 27080 28218 27108 30676
rect 27068 28212 27120 28218
rect 27068 28154 27120 28160
rect 26424 27668 26476 27674
rect 26424 27610 26476 27616
rect 27724 27606 27752 30676
rect 27712 27600 27764 27606
rect 27712 27542 27764 27548
rect 28368 27402 28396 30676
rect 29012 28082 29040 30676
rect 29000 28076 29052 28082
rect 29000 28018 29052 28024
rect 28356 27396 28408 27402
rect 28356 27338 28408 27344
rect 26056 27124 26108 27130
rect 26056 27066 26108 27072
rect 26240 27124 26292 27130
rect 26240 27066 26292 27072
rect 26332 27124 26384 27130
rect 26332 27066 26384 27072
rect 25780 26988 25832 26994
rect 25780 26930 25832 26936
rect 25964 26988 26016 26994
rect 25964 26930 26016 26936
rect 25504 26920 25556 26926
rect 25504 26862 25556 26868
rect 25412 26444 25464 26450
rect 25412 26386 25464 26392
rect 25516 26330 25544 26862
rect 26252 26450 26280 27066
rect 26516 26988 26568 26994
rect 26516 26930 26568 26936
rect 26240 26444 26292 26450
rect 26240 26386 26292 26392
rect 25228 26308 25280 26314
rect 25228 26250 25280 26256
rect 25332 26302 25544 26330
rect 25596 26376 25648 26382
rect 25596 26318 25648 26324
rect 26332 26376 26384 26382
rect 26332 26318 26384 26324
rect 25136 25968 25188 25974
rect 25136 25910 25188 25916
rect 24860 25900 24912 25906
rect 24860 25842 24912 25848
rect 25044 25900 25096 25906
rect 25044 25842 25096 25848
rect 24676 24336 24728 24342
rect 24676 24278 24728 24284
rect 23756 24200 23808 24206
rect 22926 24168 22982 24177
rect 23756 24142 23808 24148
rect 22926 24103 22982 24112
rect 22940 23186 22968 24103
rect 24872 24070 24900 25842
rect 25044 24744 25096 24750
rect 25044 24686 25096 24692
rect 25056 24274 25084 24686
rect 25044 24268 25096 24274
rect 25044 24210 25096 24216
rect 25148 24206 25176 25910
rect 25240 24818 25268 26250
rect 25332 25294 25360 26302
rect 25412 26240 25464 26246
rect 25412 26182 25464 26188
rect 25424 26042 25452 26182
rect 25412 26036 25464 26042
rect 25412 25978 25464 25984
rect 25608 25974 25636 26318
rect 25688 26240 25740 26246
rect 25688 26182 25740 26188
rect 25596 25968 25648 25974
rect 25596 25910 25648 25916
rect 25608 25770 25636 25910
rect 25504 25764 25556 25770
rect 25504 25706 25556 25712
rect 25596 25764 25648 25770
rect 25596 25706 25648 25712
rect 25516 25650 25544 25706
rect 25516 25622 25636 25650
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25228 24812 25280 24818
rect 25228 24754 25280 24760
rect 24952 24200 25004 24206
rect 25136 24200 25188 24206
rect 25004 24148 25084 24154
rect 24952 24142 25084 24148
rect 25136 24142 25188 24148
rect 24964 24126 25084 24142
rect 24492 24064 24544 24070
rect 24492 24006 24544 24012
rect 24768 24064 24820 24070
rect 24768 24006 24820 24012
rect 24860 24064 24912 24070
rect 24860 24006 24912 24012
rect 23480 23860 23532 23866
rect 23480 23802 23532 23808
rect 23296 23656 23348 23662
rect 23296 23598 23348 23604
rect 23492 23644 23520 23802
rect 23572 23656 23624 23662
rect 23492 23616 23572 23644
rect 23308 23322 23336 23598
rect 23296 23316 23348 23322
rect 23296 23258 23348 23264
rect 22928 23180 22980 23186
rect 22928 23122 22980 23128
rect 23112 23112 23164 23118
rect 23112 23054 23164 23060
rect 22652 23044 22704 23050
rect 22652 22986 22704 22992
rect 23020 22976 23072 22982
rect 23020 22918 23072 22924
rect 23032 22778 23060 22918
rect 23020 22772 23072 22778
rect 23020 22714 23072 22720
rect 23124 22574 23152 23054
rect 23112 22568 23164 22574
rect 23112 22510 23164 22516
rect 22652 21140 22704 21146
rect 22652 21082 22704 21088
rect 22560 20528 22612 20534
rect 22560 20470 22612 20476
rect 22572 20398 22600 20470
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22664 20058 22692 21082
rect 22652 20052 22704 20058
rect 22652 19994 22704 20000
rect 23296 20052 23348 20058
rect 23296 19994 23348 20000
rect 22560 19916 22612 19922
rect 22560 19858 22612 19864
rect 22572 19553 22600 19858
rect 22928 19712 22980 19718
rect 22928 19654 22980 19660
rect 22558 19544 22614 19553
rect 22558 19479 22614 19488
rect 22428 19400 22508 19428
rect 22376 19382 22428 19388
rect 22284 19236 22336 19242
rect 22284 19178 22336 19184
rect 22744 18692 22796 18698
rect 22744 18634 22796 18640
rect 22560 18420 22612 18426
rect 22560 18362 22612 18368
rect 22060 18244 22140 18272
rect 22008 18226 22060 18232
rect 21836 17734 21956 17762
rect 21732 17196 21784 17202
rect 21732 17138 21784 17144
rect 21744 16658 21772 17138
rect 21732 16652 21784 16658
rect 21732 16594 21784 16600
rect 21640 16584 21692 16590
rect 21454 16552 21510 16561
rect 21640 16526 21692 16532
rect 21454 16487 21456 16496
rect 21508 16487 21510 16496
rect 21456 16458 21508 16464
rect 21640 16040 21692 16046
rect 21640 15982 21692 15988
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 21468 15026 21496 15506
rect 21652 15502 21680 15982
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 21652 15026 21680 15438
rect 21456 15020 21508 15026
rect 21640 15020 21692 15026
rect 21508 14980 21588 15008
rect 21456 14962 21508 14968
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21180 14476 21232 14482
rect 21180 14418 21232 14424
rect 20996 14408 21048 14414
rect 20996 14350 21048 14356
rect 20904 13796 20956 13802
rect 20904 13738 20956 13744
rect 21456 13796 21508 13802
rect 21456 13738 21508 13744
rect 21468 13394 21496 13738
rect 21456 13388 21508 13394
rect 21456 13330 21508 13336
rect 21560 13326 21588 14980
rect 21640 14962 21692 14968
rect 21836 14890 21864 17734
rect 21916 17672 21968 17678
rect 21916 17614 21968 17620
rect 21824 14884 21876 14890
rect 21824 14826 21876 14832
rect 21928 14804 21956 17614
rect 22008 14816 22060 14822
rect 21928 14776 22008 14804
rect 22008 14758 22060 14764
rect 22020 14346 22048 14758
rect 22112 14482 22140 18244
rect 22468 18148 22520 18154
rect 22468 18090 22520 18096
rect 22284 18080 22336 18086
rect 22284 18022 22336 18028
rect 22296 17542 22324 18022
rect 22480 17746 22508 18090
rect 22468 17740 22520 17746
rect 22468 17682 22520 17688
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 22468 17536 22520 17542
rect 22468 17478 22520 17484
rect 22284 16448 22336 16454
rect 22284 16390 22336 16396
rect 22296 16182 22324 16390
rect 22284 16176 22336 16182
rect 22284 16118 22336 16124
rect 22192 15088 22244 15094
rect 22192 15030 22244 15036
rect 22100 14476 22152 14482
rect 22100 14418 22152 14424
rect 21824 14340 21876 14346
rect 21824 14282 21876 14288
rect 22008 14340 22060 14346
rect 22008 14282 22060 14288
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21284 12986 21312 13262
rect 21836 13161 21864 14282
rect 22100 13932 22152 13938
rect 22204 13920 22232 15030
rect 22376 15020 22428 15026
rect 22376 14962 22428 14968
rect 22388 14074 22416 14962
rect 22376 14068 22428 14074
rect 22376 14010 22428 14016
rect 22152 13892 22232 13920
rect 22100 13874 22152 13880
rect 22284 13864 22336 13870
rect 22284 13806 22336 13812
rect 22008 13796 22060 13802
rect 22060 13756 22232 13784
rect 22008 13738 22060 13744
rect 22098 13696 22154 13705
rect 22098 13631 22154 13640
rect 22008 13456 22060 13462
rect 22008 13398 22060 13404
rect 21822 13152 21878 13161
rect 21822 13087 21878 13096
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 20904 12844 20956 12850
rect 20904 12786 20956 12792
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20720 12300 20772 12306
rect 20720 12242 20772 12248
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 20088 12022 20300 12050
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 19708 11756 19760 11762
rect 19708 11698 19760 11704
rect 19720 10742 19748 11698
rect 19708 10736 19760 10742
rect 19708 10678 19760 10684
rect 19248 10668 19300 10674
rect 19248 10610 19300 10616
rect 19616 10668 19668 10674
rect 19616 10610 19668 10616
rect 20180 10606 20208 11834
rect 20272 11354 20300 12022
rect 20732 11558 20760 12242
rect 20824 12238 20852 12718
rect 20812 12232 20864 12238
rect 20812 12174 20864 12180
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20732 10810 20760 10950
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20536 10668 20588 10674
rect 20588 10628 20760 10656
rect 20536 10610 20588 10616
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 20168 10600 20220 10606
rect 20168 10542 20220 10548
rect 19248 10532 19300 10538
rect 19248 10474 19300 10480
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18880 9716 18932 9722
rect 18880 9658 18932 9664
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 17788 8078 17908 8106
rect 17684 7812 17736 7818
rect 17684 7754 17736 7760
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17236 5778 17264 6190
rect 17604 5914 17632 7346
rect 17696 7002 17724 7754
rect 17684 6996 17736 7002
rect 17684 6938 17736 6944
rect 17696 6780 17724 6938
rect 17788 6882 17816 8078
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17880 7002 17908 7958
rect 18064 7886 18092 8434
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18340 7886 18368 8026
rect 18420 8016 18472 8022
rect 18420 7958 18472 7964
rect 18432 7886 18460 7958
rect 18524 7886 18552 8910
rect 18880 8288 18932 8294
rect 18880 8230 18932 8236
rect 18052 7880 18104 7886
rect 18144 7880 18196 7886
rect 18052 7822 18104 7828
rect 18142 7848 18144 7857
rect 18328 7880 18380 7886
rect 18196 7848 18198 7857
rect 18064 7478 18092 7822
rect 18328 7822 18380 7828
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18142 7783 18198 7792
rect 18052 7472 18104 7478
rect 17958 7440 18014 7449
rect 18052 7414 18104 7420
rect 17958 7375 17960 7384
rect 18012 7375 18014 7384
rect 17960 7346 18012 7352
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 17868 6996 17920 7002
rect 17868 6938 17920 6944
rect 17788 6854 17908 6882
rect 17776 6792 17828 6798
rect 17696 6752 17776 6780
rect 17776 6734 17828 6740
rect 17880 6458 17908 6854
rect 18064 6798 18092 7142
rect 18156 6866 18184 7783
rect 18326 7440 18382 7449
rect 18326 7375 18382 7384
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 18340 6798 18368 7375
rect 18432 6934 18460 7822
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18604 7744 18656 7750
rect 18604 7686 18656 7692
rect 18524 7546 18552 7686
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18616 7410 18644 7686
rect 18788 7472 18840 7478
rect 18788 7414 18840 7420
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18800 7002 18828 7414
rect 18892 7342 18920 8230
rect 19260 8022 19288 10474
rect 19996 10470 20024 10542
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19984 10464 20036 10470
rect 19984 10406 20036 10412
rect 19904 10198 19932 10406
rect 19892 10192 19944 10198
rect 19892 10134 19944 10140
rect 20180 10130 20208 10542
rect 20168 10124 20220 10130
rect 20168 10066 20220 10072
rect 20732 9654 20760 10628
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 20628 9580 20680 9586
rect 20824 9568 20852 12174
rect 20916 9994 20944 12786
rect 21088 12436 21140 12442
rect 21140 12396 21220 12424
rect 21088 12378 21140 12384
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 20996 11688 21048 11694
rect 20996 11630 21048 11636
rect 21008 11150 21036 11630
rect 20996 11144 21048 11150
rect 20996 11086 21048 11092
rect 21008 10742 21036 11086
rect 20996 10736 21048 10742
rect 20996 10678 21048 10684
rect 20996 10260 21048 10266
rect 20996 10202 21048 10208
rect 20904 9988 20956 9994
rect 20904 9930 20956 9936
rect 20904 9580 20956 9586
rect 20824 9540 20904 9568
rect 20628 9522 20680 9528
rect 20904 9522 20956 9528
rect 19444 9382 19472 9522
rect 20640 9466 20668 9522
rect 21008 9518 21036 10202
rect 20996 9512 21048 9518
rect 19708 9444 19760 9450
rect 20640 9438 20760 9466
rect 20996 9454 21048 9460
rect 19708 9386 19760 9392
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19444 8974 19472 9318
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 19720 8906 19748 9386
rect 20732 8974 20760 9438
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 20824 8974 20852 9318
rect 21008 8974 21036 9454
rect 21100 9450 21128 12174
rect 21192 11150 21220 12396
rect 21284 12306 21312 12922
rect 22020 12850 22048 13398
rect 22112 13326 22140 13631
rect 22204 13546 22232 13756
rect 22296 13705 22324 13806
rect 22376 13796 22428 13802
rect 22376 13738 22428 13744
rect 22282 13696 22338 13705
rect 22282 13631 22338 13640
rect 22204 13518 22324 13546
rect 22296 13326 22324 13518
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 22284 13320 22336 13326
rect 22284 13262 22336 13268
rect 21824 12844 21876 12850
rect 21824 12786 21876 12792
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 21836 12374 21864 12786
rect 22020 12442 22048 12786
rect 22112 12646 22140 13262
rect 22284 13184 22336 13190
rect 22190 13152 22246 13161
rect 22284 13126 22336 13132
rect 22190 13087 22246 13096
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 22008 12436 22060 12442
rect 22008 12378 22060 12384
rect 21824 12368 21876 12374
rect 21824 12310 21876 12316
rect 21272 12300 21324 12306
rect 21272 12242 21324 12248
rect 21376 12170 21588 12186
rect 21376 12164 21600 12170
rect 21376 12158 21548 12164
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21180 11144 21232 11150
rect 21180 11086 21232 11092
rect 21284 10606 21312 11494
rect 21376 11121 21404 12158
rect 21548 12106 21600 12112
rect 22008 11212 22060 11218
rect 22008 11154 22060 11160
rect 21732 11144 21784 11150
rect 21362 11112 21418 11121
rect 21732 11086 21784 11092
rect 21362 11047 21418 11056
rect 21456 11076 21508 11082
rect 21272 10600 21324 10606
rect 21272 10542 21324 10548
rect 21088 9444 21140 9450
rect 21088 9386 21140 9392
rect 21180 9376 21232 9382
rect 21180 9318 21232 9324
rect 21192 9178 21220 9318
rect 21180 9172 21232 9178
rect 21180 9114 21232 9120
rect 20720 8968 20772 8974
rect 20720 8910 20772 8916
rect 20812 8968 20864 8974
rect 20812 8910 20864 8916
rect 20996 8968 21048 8974
rect 20996 8910 21048 8916
rect 19708 8900 19760 8906
rect 19708 8842 19760 8848
rect 19248 8016 19300 8022
rect 19248 7958 19300 7964
rect 19720 7886 19748 8842
rect 20076 7948 20128 7954
rect 20076 7890 20128 7896
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19260 7750 19288 7822
rect 19984 7812 20036 7818
rect 19984 7754 20036 7760
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 18420 6928 18472 6934
rect 18892 6882 18920 7278
rect 18420 6870 18472 6876
rect 18800 6854 18920 6882
rect 18800 6798 18828 6854
rect 19260 6798 19288 7686
rect 19708 7336 19760 7342
rect 19628 7284 19708 7290
rect 19628 7278 19760 7284
rect 19628 7262 19748 7278
rect 19996 7274 20024 7754
rect 20088 7274 20116 7890
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20168 7812 20220 7818
rect 20168 7754 20220 7760
rect 20180 7410 20208 7754
rect 20260 7744 20312 7750
rect 20260 7686 20312 7692
rect 20168 7404 20220 7410
rect 20168 7346 20220 7352
rect 20272 7342 20300 7686
rect 20350 7440 20406 7449
rect 20456 7410 20484 7822
rect 20548 7721 20576 7822
rect 20534 7712 20590 7721
rect 20534 7647 20590 7656
rect 20350 7375 20352 7384
rect 20404 7375 20406 7384
rect 20444 7404 20496 7410
rect 20352 7346 20404 7352
rect 20444 7346 20496 7352
rect 20536 7404 20588 7410
rect 20536 7346 20588 7352
rect 20260 7336 20312 7342
rect 20260 7278 20312 7284
rect 19984 7268 20036 7274
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19352 7002 19380 7142
rect 19340 6996 19392 7002
rect 19340 6938 19392 6944
rect 19628 6798 19656 7262
rect 19984 7210 20036 7216
rect 20076 7268 20128 7274
rect 20076 7210 20128 7216
rect 19708 7200 19760 7206
rect 19708 7142 19760 7148
rect 19720 6934 19748 7142
rect 19708 6928 19760 6934
rect 19708 6870 19760 6876
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 18328 6792 18380 6798
rect 18328 6734 18380 6740
rect 18420 6792 18472 6798
rect 18788 6792 18840 6798
rect 18420 6734 18472 6740
rect 18694 6760 18750 6769
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 17684 6248 17736 6254
rect 17682 6216 17684 6225
rect 17736 6216 17738 6225
rect 17682 6151 17738 6160
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 17224 5772 17276 5778
rect 17224 5714 17276 5720
rect 17880 5642 17908 6394
rect 18432 6118 18460 6734
rect 18788 6734 18840 6740
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 18694 6695 18750 6704
rect 18708 6118 18736 6695
rect 19260 6458 19288 6734
rect 19444 6458 19472 6734
rect 20548 6458 20576 7346
rect 20732 7274 20760 8910
rect 20824 7970 20852 8910
rect 21088 8356 21140 8362
rect 21088 8298 21140 8304
rect 20824 7942 21036 7970
rect 20812 7880 20864 7886
rect 20810 7848 20812 7857
rect 20904 7880 20956 7886
rect 20864 7848 20866 7857
rect 20904 7822 20956 7828
rect 20810 7783 20866 7792
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 20824 7410 20852 7686
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20720 7268 20772 7274
rect 20720 7210 20772 7216
rect 20824 6662 20852 7346
rect 20916 7274 20944 7822
rect 21008 7410 21036 7942
rect 21100 7750 21128 8298
rect 21180 7880 21232 7886
rect 21284 7857 21312 10542
rect 21376 9518 21404 11047
rect 21456 11018 21508 11024
rect 21468 10674 21496 11018
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 21468 10266 21496 10610
rect 21456 10260 21508 10266
rect 21456 10202 21508 10208
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 21456 9580 21508 9586
rect 21456 9522 21508 9528
rect 21364 9512 21416 9518
rect 21364 9454 21416 9460
rect 21376 8022 21404 9454
rect 21364 8016 21416 8022
rect 21364 7958 21416 7964
rect 21468 7886 21496 9522
rect 21652 7954 21680 10066
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 21364 7880 21416 7886
rect 21180 7822 21232 7828
rect 21270 7848 21326 7857
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 21086 7576 21142 7585
rect 21086 7511 21088 7520
rect 21140 7511 21142 7520
rect 21088 7482 21140 7488
rect 21192 7449 21220 7822
rect 21364 7822 21416 7828
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 21270 7783 21326 7792
rect 21376 7546 21404 7822
rect 21744 7818 21772 11086
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21732 7812 21784 7818
rect 21732 7754 21784 7760
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21178 7440 21234 7449
rect 20996 7404 21048 7410
rect 21178 7375 21234 7384
rect 21548 7404 21600 7410
rect 20996 7346 21048 7352
rect 21548 7346 21600 7352
rect 20904 7268 20956 7274
rect 20904 7210 20956 7216
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 20916 6458 20944 7210
rect 21560 7002 21588 7346
rect 21744 7002 21772 7754
rect 21836 7750 21864 8026
rect 22020 7954 22048 11154
rect 22204 11082 22232 13087
rect 22296 12714 22324 13126
rect 22388 12918 22416 13738
rect 22376 12912 22428 12918
rect 22376 12854 22428 12860
rect 22284 12708 22336 12714
rect 22284 12650 22336 12656
rect 22480 12102 22508 17478
rect 22572 16572 22600 18362
rect 22756 17066 22784 18634
rect 22744 17060 22796 17066
rect 22744 17002 22796 17008
rect 22940 16590 22968 19654
rect 23020 18080 23072 18086
rect 23020 18022 23072 18028
rect 22652 16584 22704 16590
rect 22572 16544 22652 16572
rect 22652 16526 22704 16532
rect 22836 16584 22888 16590
rect 22836 16526 22888 16532
rect 22928 16584 22980 16590
rect 22928 16526 22980 16532
rect 22848 15706 22876 16526
rect 22836 15700 22888 15706
rect 22836 15642 22888 15648
rect 22560 14612 22612 14618
rect 22560 14554 22612 14560
rect 22572 13870 22600 14554
rect 22940 14498 22968 16526
rect 22664 14470 22968 14498
rect 22664 14414 22692 14470
rect 22652 14408 22704 14414
rect 22652 14350 22704 14356
rect 22928 14272 22980 14278
rect 22650 14240 22706 14249
rect 22928 14214 22980 14220
rect 22650 14175 22706 14184
rect 22560 13864 22612 13870
rect 22560 13806 22612 13812
rect 22468 12096 22520 12102
rect 22468 12038 22520 12044
rect 22192 11076 22244 11082
rect 22192 11018 22244 11024
rect 22468 11008 22520 11014
rect 22468 10950 22520 10956
rect 22480 10198 22508 10950
rect 22560 10260 22612 10266
rect 22560 10202 22612 10208
rect 22468 10192 22520 10198
rect 22468 10134 22520 10140
rect 22572 8090 22600 10202
rect 22560 8084 22612 8090
rect 22560 8026 22612 8032
rect 22008 7948 22060 7954
rect 22008 7890 22060 7896
rect 21824 7744 21876 7750
rect 21824 7686 21876 7692
rect 21914 7712 21970 7721
rect 21914 7647 21970 7656
rect 21928 7546 21956 7647
rect 21916 7540 21968 7546
rect 21916 7482 21968 7488
rect 22020 7410 22048 7890
rect 22572 7410 22600 8026
rect 22664 7818 22692 14175
rect 22940 13938 22968 14214
rect 22928 13932 22980 13938
rect 22928 13874 22980 13880
rect 22744 13524 22796 13530
rect 22744 13466 22796 13472
rect 22756 12986 22784 13466
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22928 13320 22980 13326
rect 22928 13262 22980 13268
rect 22744 12980 22796 12986
rect 22744 12922 22796 12928
rect 22848 11898 22876 13262
rect 22836 11892 22888 11898
rect 22836 11834 22888 11840
rect 22836 11756 22888 11762
rect 22836 11698 22888 11704
rect 22744 11620 22796 11626
rect 22744 11562 22796 11568
rect 22756 10062 22784 11562
rect 22848 10742 22876 11698
rect 22836 10736 22888 10742
rect 22836 10678 22888 10684
rect 22744 10056 22796 10062
rect 22744 9998 22796 10004
rect 22848 9926 22876 10678
rect 22836 9920 22888 9926
rect 22836 9862 22888 9868
rect 22940 8634 22968 13262
rect 23032 11558 23060 18022
rect 23112 16992 23164 16998
rect 23112 16934 23164 16940
rect 23124 16794 23152 16934
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 23204 16448 23256 16454
rect 23204 16390 23256 16396
rect 23216 16250 23244 16390
rect 23204 16244 23256 16250
rect 23204 16186 23256 16192
rect 23308 16130 23336 19994
rect 23492 19922 23520 23616
rect 23572 23598 23624 23604
rect 24032 23656 24084 23662
rect 24032 23598 24084 23604
rect 24044 23322 24072 23598
rect 24032 23316 24084 23322
rect 24032 23258 24084 23264
rect 24504 23186 24532 24006
rect 24780 23186 24808 24006
rect 25056 23662 25084 24126
rect 25332 24018 25360 25230
rect 25608 25158 25636 25622
rect 25596 25152 25648 25158
rect 25596 25094 25648 25100
rect 25608 24750 25636 25094
rect 25596 24744 25648 24750
rect 25596 24686 25648 24692
rect 25608 24274 25636 24686
rect 25596 24268 25648 24274
rect 25596 24210 25648 24216
rect 25148 23990 25360 24018
rect 25044 23656 25096 23662
rect 25044 23598 25096 23604
rect 24492 23180 24544 23186
rect 24492 23122 24544 23128
rect 24768 23180 24820 23186
rect 24768 23122 24820 23128
rect 24216 23112 24268 23118
rect 24216 23054 24268 23060
rect 24228 22234 24256 23054
rect 24860 22976 24912 22982
rect 24860 22918 24912 22924
rect 24676 22500 24728 22506
rect 24676 22442 24728 22448
rect 24216 22228 24268 22234
rect 24216 22170 24268 22176
rect 24228 21350 24256 22170
rect 24688 22030 24716 22442
rect 24872 22030 24900 22918
rect 25148 22778 25176 23990
rect 25504 23792 25556 23798
rect 25504 23734 25556 23740
rect 25412 23656 25464 23662
rect 25412 23598 25464 23604
rect 25424 23118 25452 23598
rect 25412 23112 25464 23118
rect 25412 23054 25464 23060
rect 25412 22976 25464 22982
rect 25412 22918 25464 22924
rect 25136 22772 25188 22778
rect 25136 22714 25188 22720
rect 24952 22500 25004 22506
rect 24952 22442 25004 22448
rect 24584 22024 24636 22030
rect 24584 21966 24636 21972
rect 24676 22024 24728 22030
rect 24676 21966 24728 21972
rect 24860 22024 24912 22030
rect 24860 21966 24912 21972
rect 24596 21894 24624 21966
rect 24584 21888 24636 21894
rect 24584 21830 24636 21836
rect 24596 21554 24624 21830
rect 24688 21622 24716 21966
rect 24768 21888 24820 21894
rect 24768 21830 24820 21836
rect 24676 21616 24728 21622
rect 24676 21558 24728 21564
rect 24780 21554 24808 21830
rect 24584 21548 24636 21554
rect 24584 21490 24636 21496
rect 24768 21548 24820 21554
rect 24768 21490 24820 21496
rect 24676 21480 24728 21486
rect 24676 21422 24728 21428
rect 24216 21344 24268 21350
rect 24216 21286 24268 21292
rect 23572 20936 23624 20942
rect 23572 20878 23624 20884
rect 23584 20602 23612 20878
rect 24032 20868 24084 20874
rect 24032 20810 24084 20816
rect 23572 20596 23624 20602
rect 23572 20538 23624 20544
rect 24044 20398 24072 20810
rect 24032 20392 24084 20398
rect 24032 20334 24084 20340
rect 23480 19916 23532 19922
rect 23480 19858 23532 19864
rect 23388 18828 23440 18834
rect 23492 18816 23520 19858
rect 23440 18788 23520 18816
rect 23388 18770 23440 18776
rect 23216 16102 23336 16130
rect 23400 16114 23428 18770
rect 24044 18698 24072 20334
rect 24228 18970 24256 21286
rect 24688 20942 24716 21422
rect 24964 21418 24992 22442
rect 25148 22094 25176 22714
rect 25228 22500 25280 22506
rect 25228 22442 25280 22448
rect 25240 22234 25268 22442
rect 25228 22228 25280 22234
rect 25228 22170 25280 22176
rect 25320 22228 25372 22234
rect 25320 22170 25372 22176
rect 25148 22066 25268 22094
rect 25136 21888 25188 21894
rect 25136 21830 25188 21836
rect 25148 21690 25176 21830
rect 25240 21690 25268 22066
rect 25136 21684 25188 21690
rect 25136 21626 25188 21632
rect 25228 21684 25280 21690
rect 25228 21626 25280 21632
rect 24952 21412 25004 21418
rect 24952 21354 25004 21360
rect 25044 21004 25096 21010
rect 25148 20992 25176 21626
rect 25096 20964 25176 20992
rect 25044 20946 25096 20952
rect 24676 20936 24728 20942
rect 24676 20878 24728 20884
rect 24688 19922 24716 20878
rect 25240 20534 25268 21626
rect 25332 21622 25360 22170
rect 25424 22166 25452 22918
rect 25412 22160 25464 22166
rect 25412 22102 25464 22108
rect 25320 21616 25372 21622
rect 25320 21558 25372 21564
rect 25412 21616 25464 21622
rect 25412 21558 25464 21564
rect 25424 20874 25452 21558
rect 25412 20868 25464 20874
rect 25412 20810 25464 20816
rect 25228 20528 25280 20534
rect 25228 20470 25280 20476
rect 24676 19916 24728 19922
rect 24676 19858 24728 19864
rect 25516 19718 25544 23734
rect 25596 23724 25648 23730
rect 25596 23666 25648 23672
rect 25608 23254 25636 23666
rect 25596 23248 25648 23254
rect 25596 23190 25648 23196
rect 25608 22778 25636 23190
rect 25596 22772 25648 22778
rect 25596 22714 25648 22720
rect 25700 22710 25728 26182
rect 26344 25906 26372 26318
rect 26424 26308 26476 26314
rect 26424 26250 26476 26256
rect 26436 25906 26464 26250
rect 26528 26042 26556 26930
rect 26792 26852 26844 26858
rect 26792 26794 26844 26800
rect 26804 26586 26832 26794
rect 27068 26784 27120 26790
rect 27068 26726 27120 26732
rect 27712 26784 27764 26790
rect 27712 26726 27764 26732
rect 26792 26580 26844 26586
rect 26792 26522 26844 26528
rect 26792 26376 26844 26382
rect 26792 26318 26844 26324
rect 26516 26036 26568 26042
rect 26516 25978 26568 25984
rect 26332 25900 26384 25906
rect 26332 25842 26384 25848
rect 26424 25900 26476 25906
rect 26424 25842 26476 25848
rect 26344 25498 26372 25842
rect 25872 25492 25924 25498
rect 25872 25434 25924 25440
rect 26332 25492 26384 25498
rect 26332 25434 26384 25440
rect 25884 24818 25912 25434
rect 26240 25424 26292 25430
rect 26240 25366 26292 25372
rect 26252 24886 26280 25366
rect 26332 25220 26384 25226
rect 26332 25162 26384 25168
rect 26344 24954 26372 25162
rect 26332 24948 26384 24954
rect 26332 24890 26384 24896
rect 26240 24880 26292 24886
rect 26240 24822 26292 24828
rect 25780 24812 25832 24818
rect 25780 24754 25832 24760
rect 25872 24812 25924 24818
rect 25872 24754 25924 24760
rect 25792 23322 25820 24754
rect 25884 24614 25912 24754
rect 25872 24608 25924 24614
rect 25872 24550 25924 24556
rect 25884 24410 25912 24550
rect 25872 24404 25924 24410
rect 25872 24346 25924 24352
rect 25964 24268 26016 24274
rect 25964 24210 26016 24216
rect 25872 24132 25924 24138
rect 25872 24074 25924 24080
rect 25884 23798 25912 24074
rect 25976 23798 26004 24210
rect 26056 24064 26108 24070
rect 26056 24006 26108 24012
rect 25872 23792 25924 23798
rect 25872 23734 25924 23740
rect 25964 23792 26016 23798
rect 25964 23734 26016 23740
rect 26068 23730 26096 24006
rect 26252 23882 26280 24822
rect 26344 24342 26372 24890
rect 26332 24336 26384 24342
rect 26332 24278 26384 24284
rect 26160 23866 26280 23882
rect 26436 23866 26464 25842
rect 26804 25838 26832 26318
rect 26792 25832 26844 25838
rect 26792 25774 26844 25780
rect 27080 25158 27108 26726
rect 27724 26625 27752 26726
rect 27710 26616 27766 26625
rect 27710 26551 27766 26560
rect 27528 26512 27580 26518
rect 27528 26454 27580 26460
rect 27342 26344 27398 26353
rect 27342 26279 27398 26288
rect 27068 25152 27120 25158
rect 27068 25094 27120 25100
rect 26884 24608 26936 24614
rect 26884 24550 26936 24556
rect 26896 24206 26924 24550
rect 27080 24206 27108 25094
rect 27160 24608 27212 24614
rect 27160 24550 27212 24556
rect 27172 24274 27200 24550
rect 27160 24268 27212 24274
rect 27160 24210 27212 24216
rect 27356 24206 27384 26279
rect 27540 25945 27568 26454
rect 27526 25936 27582 25945
rect 27526 25871 27582 25880
rect 27528 25288 27580 25294
rect 27528 25230 27580 25236
rect 27710 25256 27766 25265
rect 27436 25220 27488 25226
rect 27436 25162 27488 25168
rect 26884 24200 26936 24206
rect 26884 24142 26936 24148
rect 27068 24200 27120 24206
rect 27068 24142 27120 24148
rect 27344 24200 27396 24206
rect 27344 24142 27396 24148
rect 27068 24064 27120 24070
rect 27068 24006 27120 24012
rect 26148 23860 26280 23866
rect 26200 23854 26280 23860
rect 26148 23802 26200 23808
rect 26056 23724 26108 23730
rect 26056 23666 26108 23672
rect 25780 23316 25832 23322
rect 25780 23258 25832 23264
rect 25688 22704 25740 22710
rect 25688 22646 25740 22652
rect 25596 22568 25648 22574
rect 25596 22510 25648 22516
rect 25608 22030 25636 22510
rect 25700 22506 25728 22646
rect 25688 22500 25740 22506
rect 25688 22442 25740 22448
rect 25792 22438 25820 23258
rect 26068 23118 26096 23666
rect 26252 23186 26280 23854
rect 26424 23860 26476 23866
rect 26424 23802 26476 23808
rect 26976 23724 27028 23730
rect 26976 23666 27028 23672
rect 26988 23322 27016 23666
rect 26976 23316 27028 23322
rect 26976 23258 27028 23264
rect 26240 23180 26292 23186
rect 26240 23122 26292 23128
rect 26608 23180 26660 23186
rect 26608 23122 26660 23128
rect 26056 23112 26108 23118
rect 26056 23054 26108 23060
rect 26620 23050 26648 23122
rect 26608 23044 26660 23050
rect 26608 22986 26660 22992
rect 26148 22976 26200 22982
rect 26148 22918 26200 22924
rect 26160 22778 26188 22918
rect 26148 22772 26200 22778
rect 26148 22714 26200 22720
rect 26056 22704 26108 22710
rect 26056 22646 26108 22652
rect 25964 22636 26016 22642
rect 25964 22578 26016 22584
rect 25780 22432 25832 22438
rect 25780 22374 25832 22380
rect 25688 22092 25740 22098
rect 25740 22052 25820 22080
rect 25688 22034 25740 22040
rect 25596 22024 25648 22030
rect 25596 21966 25648 21972
rect 25792 22012 25820 22052
rect 25872 22024 25924 22030
rect 25792 21984 25872 22012
rect 25688 21888 25740 21894
rect 25688 21830 25740 21836
rect 25700 19786 25728 21830
rect 25688 19780 25740 19786
rect 25688 19722 25740 19728
rect 24860 19712 24912 19718
rect 24860 19654 24912 19660
rect 25504 19712 25556 19718
rect 25504 19654 25556 19660
rect 24216 18964 24268 18970
rect 24216 18906 24268 18912
rect 24032 18692 24084 18698
rect 24032 18634 24084 18640
rect 24044 17610 24072 18634
rect 24492 17740 24544 17746
rect 24492 17682 24544 17688
rect 24032 17604 24084 17610
rect 24032 17546 24084 17552
rect 23480 17196 23532 17202
rect 23480 17138 23532 17144
rect 23388 16108 23440 16114
rect 23216 15638 23244 16102
rect 23388 16050 23440 16056
rect 23492 15638 23520 17138
rect 24044 16726 24072 17546
rect 24216 17536 24268 17542
rect 24216 17478 24268 17484
rect 24228 17202 24256 17478
rect 24216 17196 24268 17202
rect 24216 17138 24268 17144
rect 24032 16720 24084 16726
rect 24032 16662 24084 16668
rect 23572 16584 23624 16590
rect 23572 16526 23624 16532
rect 23848 16584 23900 16590
rect 23848 16526 23900 16532
rect 23584 15706 23612 16526
rect 23756 16040 23808 16046
rect 23756 15982 23808 15988
rect 23572 15700 23624 15706
rect 23572 15642 23624 15648
rect 23204 15632 23256 15638
rect 23110 15600 23166 15609
rect 23204 15574 23256 15580
rect 23480 15632 23532 15638
rect 23480 15574 23532 15580
rect 23110 15535 23166 15544
rect 23124 15502 23152 15535
rect 23112 15496 23164 15502
rect 23112 15438 23164 15444
rect 23124 14618 23152 15438
rect 23112 14612 23164 14618
rect 23112 14554 23164 14560
rect 23124 13870 23152 14554
rect 23112 13864 23164 13870
rect 23112 13806 23164 13812
rect 23216 12170 23244 15574
rect 23572 15496 23624 15502
rect 23572 15438 23624 15444
rect 23388 15156 23440 15162
rect 23388 15098 23440 15104
rect 23296 14884 23348 14890
rect 23296 14826 23348 14832
rect 23308 14634 23336 14826
rect 23400 14822 23428 15098
rect 23584 14890 23612 15438
rect 23768 15434 23796 15982
rect 23756 15428 23808 15434
rect 23756 15370 23808 15376
rect 23768 15094 23796 15370
rect 23860 15162 23888 16526
rect 24044 16250 24072 16662
rect 24504 16590 24532 17682
rect 24872 17134 24900 19654
rect 25228 17196 25280 17202
rect 25228 17138 25280 17144
rect 24860 17128 24912 17134
rect 24860 17070 24912 17076
rect 24492 16584 24544 16590
rect 24492 16526 24544 16532
rect 24032 16244 24084 16250
rect 24032 16186 24084 16192
rect 24216 15496 24268 15502
rect 24216 15438 24268 15444
rect 24032 15360 24084 15366
rect 24032 15302 24084 15308
rect 23848 15156 23900 15162
rect 23848 15098 23900 15104
rect 23756 15088 23808 15094
rect 23756 15030 23808 15036
rect 24044 15026 24072 15302
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 24032 15020 24084 15026
rect 24032 14962 24084 14968
rect 23572 14884 23624 14890
rect 23572 14826 23624 14832
rect 23388 14816 23440 14822
rect 23388 14758 23440 14764
rect 23308 14606 23428 14634
rect 23296 14544 23348 14550
rect 23296 14486 23348 14492
rect 23308 13938 23336 14486
rect 23400 14346 23428 14606
rect 23756 14612 23808 14618
rect 23756 14554 23808 14560
rect 23664 14476 23716 14482
rect 23664 14418 23716 14424
rect 23388 14340 23440 14346
rect 23388 14282 23440 14288
rect 23400 13938 23428 14282
rect 23572 14272 23624 14278
rect 23572 14214 23624 14220
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23296 13932 23348 13938
rect 23296 13874 23348 13880
rect 23388 13932 23440 13938
rect 23388 13874 23440 13880
rect 23388 13796 23440 13802
rect 23388 13738 23440 13744
rect 23296 12980 23348 12986
rect 23296 12922 23348 12928
rect 23204 12164 23256 12170
rect 23204 12106 23256 12112
rect 23112 12096 23164 12102
rect 23112 12038 23164 12044
rect 23020 11552 23072 11558
rect 23020 11494 23072 11500
rect 23124 11286 23152 12038
rect 23308 11898 23336 12922
rect 23296 11892 23348 11898
rect 23296 11834 23348 11840
rect 23204 11756 23256 11762
rect 23204 11698 23256 11704
rect 23296 11756 23348 11762
rect 23296 11698 23348 11704
rect 23020 11280 23072 11286
rect 23020 11222 23072 11228
rect 23112 11280 23164 11286
rect 23112 11222 23164 11228
rect 23032 11150 23060 11222
rect 23020 11144 23072 11150
rect 23216 11132 23244 11698
rect 23020 11086 23072 11092
rect 23124 11104 23244 11132
rect 23020 11008 23072 11014
rect 23020 10950 23072 10956
rect 23032 10470 23060 10950
rect 23124 10742 23152 11104
rect 23308 11014 23336 11698
rect 23296 11008 23348 11014
rect 23296 10950 23348 10956
rect 23400 10826 23428 13738
rect 23492 13394 23520 14010
rect 23584 14006 23612 14214
rect 23572 14000 23624 14006
rect 23572 13942 23624 13948
rect 23572 13864 23624 13870
rect 23572 13806 23624 13812
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 23480 12708 23532 12714
rect 23480 12650 23532 12656
rect 23492 11898 23520 12650
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23480 11756 23532 11762
rect 23480 11698 23532 11704
rect 23492 11354 23520 11698
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23584 10826 23612 13806
rect 23676 11626 23704 14418
rect 23768 14414 23796 14554
rect 23952 14550 23980 14962
rect 23940 14544 23992 14550
rect 23940 14486 23992 14492
rect 23756 14408 23808 14414
rect 23756 14350 23808 14356
rect 23940 14408 23992 14414
rect 23940 14350 23992 14356
rect 23952 13462 23980 14350
rect 23940 13456 23992 13462
rect 23940 13398 23992 13404
rect 24044 13394 24072 14962
rect 24228 14958 24256 15438
rect 24216 14952 24268 14958
rect 24216 14894 24268 14900
rect 24228 14414 24256 14894
rect 24216 14408 24268 14414
rect 24216 14350 24268 14356
rect 24228 13870 24256 14350
rect 24504 14346 24532 16526
rect 24872 16522 24900 17070
rect 24860 16516 24912 16522
rect 24860 16458 24912 16464
rect 24768 15700 24820 15706
rect 24768 15642 24820 15648
rect 24780 14550 24808 15642
rect 24872 15570 24900 16458
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24768 14544 24820 14550
rect 24768 14486 24820 14492
rect 24492 14340 24544 14346
rect 24492 14282 24544 14288
rect 24216 13864 24268 13870
rect 24216 13806 24268 13812
rect 24032 13388 24084 13394
rect 24032 13330 24084 13336
rect 24032 11688 24084 11694
rect 24032 11630 24084 11636
rect 23664 11620 23716 11626
rect 23664 11562 23716 11568
rect 23664 11348 23716 11354
rect 23664 11290 23716 11296
rect 23308 10798 23428 10826
rect 23492 10798 23612 10826
rect 23676 10810 23704 11290
rect 24044 11218 24072 11630
rect 24504 11286 24532 14282
rect 24780 14074 24808 14486
rect 25134 14240 25190 14249
rect 25134 14175 25190 14184
rect 24768 14068 24820 14074
rect 24768 14010 24820 14016
rect 24780 13326 24808 14010
rect 25148 14006 25176 14175
rect 25136 14000 25188 14006
rect 25136 13942 25188 13948
rect 24952 13932 25004 13938
rect 24952 13874 25004 13880
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24492 11280 24544 11286
rect 24492 11222 24544 11228
rect 23940 11212 23992 11218
rect 23940 11154 23992 11160
rect 24032 11212 24084 11218
rect 24032 11154 24084 11160
rect 23952 11082 23980 11154
rect 23756 11076 23808 11082
rect 23756 11018 23808 11024
rect 23848 11076 23900 11082
rect 23848 11018 23900 11024
rect 23940 11076 23992 11082
rect 23940 11018 23992 11024
rect 23112 10736 23164 10742
rect 23112 10678 23164 10684
rect 23020 10464 23072 10470
rect 23020 10406 23072 10412
rect 23308 9586 23336 10798
rect 23492 10742 23520 10798
rect 23480 10736 23532 10742
rect 23480 10678 23532 10684
rect 23584 10198 23612 10798
rect 23664 10804 23716 10810
rect 23664 10746 23716 10752
rect 23664 10260 23716 10266
rect 23664 10202 23716 10208
rect 23572 10192 23624 10198
rect 23572 10134 23624 10140
rect 23572 9920 23624 9926
rect 23572 9862 23624 9868
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 23480 9376 23532 9382
rect 23480 9318 23532 9324
rect 23492 8974 23520 9318
rect 23480 8968 23532 8974
rect 23480 8910 23532 8916
rect 23296 8832 23348 8838
rect 23296 8774 23348 8780
rect 22928 8628 22980 8634
rect 22928 8570 22980 8576
rect 23308 8566 23336 8774
rect 23296 8560 23348 8566
rect 23296 8502 23348 8508
rect 23584 8498 23612 9862
rect 23676 8974 23704 10202
rect 23768 10130 23796 11018
rect 23860 10810 23888 11018
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 23756 10124 23808 10130
rect 23756 10066 23808 10072
rect 23860 9382 23888 10746
rect 23952 10266 23980 11018
rect 24044 10742 24072 11154
rect 24032 10736 24084 10742
rect 24032 10678 24084 10684
rect 24584 10532 24636 10538
rect 24504 10492 24584 10520
rect 24504 10418 24532 10492
rect 24584 10474 24636 10480
rect 24768 10532 24820 10538
rect 24768 10474 24820 10480
rect 24320 10390 24532 10418
rect 24676 10464 24728 10470
rect 24676 10406 24728 10412
rect 23940 10260 23992 10266
rect 23940 10202 23992 10208
rect 24320 10130 24348 10390
rect 24688 10130 24716 10406
rect 24308 10124 24360 10130
rect 24308 10066 24360 10072
rect 24400 10124 24452 10130
rect 24400 10066 24452 10072
rect 24676 10124 24728 10130
rect 24676 10066 24728 10072
rect 24216 9920 24268 9926
rect 24216 9862 24268 9868
rect 24228 9586 24256 9862
rect 24216 9580 24268 9586
rect 24216 9522 24268 9528
rect 23848 9376 23900 9382
rect 23848 9318 23900 9324
rect 24228 9058 24256 9522
rect 24136 9030 24256 9058
rect 23664 8968 23716 8974
rect 23664 8910 23716 8916
rect 23940 8832 23992 8838
rect 23940 8774 23992 8780
rect 23952 8498 23980 8774
rect 24136 8634 24164 9030
rect 24308 8900 24360 8906
rect 24308 8842 24360 8848
rect 24124 8628 24176 8634
rect 24124 8570 24176 8576
rect 23388 8492 23440 8498
rect 23388 8434 23440 8440
rect 23572 8492 23624 8498
rect 23572 8434 23624 8440
rect 23848 8492 23900 8498
rect 23848 8434 23900 8440
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 22928 8016 22980 8022
rect 22928 7958 22980 7964
rect 22744 7880 22796 7886
rect 22744 7822 22796 7828
rect 22652 7812 22704 7818
rect 22652 7754 22704 7760
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 22560 7404 22612 7410
rect 22560 7346 22612 7352
rect 22664 7290 22692 7754
rect 22756 7478 22784 7822
rect 22940 7478 22968 7958
rect 23400 7886 23428 8434
rect 23756 8356 23808 8362
rect 23756 8298 23808 8304
rect 23768 7993 23796 8298
rect 23754 7984 23810 7993
rect 23754 7919 23810 7928
rect 23860 7886 23888 8434
rect 24032 8424 24084 8430
rect 24032 8366 24084 8372
rect 24044 8090 24072 8366
rect 24136 8294 24164 8570
rect 24320 8498 24348 8842
rect 24308 8492 24360 8498
rect 24308 8434 24360 8440
rect 24308 8356 24360 8362
rect 24308 8298 24360 8304
rect 24124 8288 24176 8294
rect 24124 8230 24176 8236
rect 24216 8288 24268 8294
rect 24216 8230 24268 8236
rect 24032 8084 24084 8090
rect 24032 8026 24084 8032
rect 23388 7880 23440 7886
rect 23388 7822 23440 7828
rect 23848 7880 23900 7886
rect 23848 7822 23900 7828
rect 24124 7880 24176 7886
rect 24124 7822 24176 7828
rect 23020 7744 23072 7750
rect 23020 7686 23072 7692
rect 22744 7472 22796 7478
rect 22744 7414 22796 7420
rect 22928 7472 22980 7478
rect 22928 7414 22980 7420
rect 22572 7274 22692 7290
rect 22560 7268 22692 7274
rect 22612 7262 22692 7268
rect 22560 7210 22612 7216
rect 21548 6996 21600 7002
rect 21548 6938 21600 6944
rect 21732 6996 21784 7002
rect 21732 6938 21784 6944
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 21560 6322 21588 6938
rect 22008 6792 22060 6798
rect 22008 6734 22060 6740
rect 22020 6458 22048 6734
rect 22008 6452 22060 6458
rect 22008 6394 22060 6400
rect 23032 6322 23060 7686
rect 23400 7342 23428 7822
rect 23480 7744 23532 7750
rect 23480 7686 23532 7692
rect 23388 7336 23440 7342
rect 23388 7278 23440 7284
rect 23492 7002 23520 7686
rect 24136 7342 24164 7822
rect 24228 7546 24256 8230
rect 24216 7540 24268 7546
rect 24216 7482 24268 7488
rect 24228 7410 24256 7482
rect 24320 7410 24348 8298
rect 24412 7954 24440 10066
rect 24780 8838 24808 10474
rect 24964 9994 24992 13874
rect 25240 11082 25268 17138
rect 25792 14074 25820 21984
rect 25872 21966 25924 21972
rect 25976 21962 26004 22578
rect 26068 22522 26096 22646
rect 27080 22642 27108 24006
rect 27448 23118 27476 25162
rect 27540 24410 27568 25230
rect 27710 25191 27766 25200
rect 27724 25158 27752 25191
rect 27712 25152 27764 25158
rect 27712 25094 27764 25100
rect 27712 24608 27764 24614
rect 27710 24576 27712 24585
rect 27764 24576 27766 24585
rect 27710 24511 27766 24520
rect 27528 24404 27580 24410
rect 27528 24346 27580 24352
rect 27712 24064 27764 24070
rect 27712 24006 27764 24012
rect 27724 23905 27752 24006
rect 27710 23896 27766 23905
rect 27710 23831 27766 23840
rect 27528 23520 27580 23526
rect 27528 23462 27580 23468
rect 27540 23225 27568 23462
rect 27526 23216 27582 23225
rect 27526 23151 27582 23160
rect 27436 23112 27488 23118
rect 27436 23054 27488 23060
rect 27160 23044 27212 23050
rect 27160 22986 27212 22992
rect 27172 22778 27200 22986
rect 27344 22976 27396 22982
rect 27344 22918 27396 22924
rect 27160 22772 27212 22778
rect 27160 22714 27212 22720
rect 27356 22642 27384 22918
rect 27068 22636 27120 22642
rect 27068 22578 27120 22584
rect 27344 22636 27396 22642
rect 27344 22578 27396 22584
rect 26148 22568 26200 22574
rect 26068 22516 26148 22522
rect 26068 22510 26200 22516
rect 26068 22494 26188 22510
rect 26056 22432 26108 22438
rect 26056 22374 26108 22380
rect 25964 21956 26016 21962
rect 25964 21898 26016 21904
rect 25872 21888 25924 21894
rect 25872 21830 25924 21836
rect 25884 21350 25912 21830
rect 26068 21486 26096 22374
rect 26160 22094 26188 22494
rect 26160 22066 26280 22094
rect 26252 22030 26280 22066
rect 26240 22024 26292 22030
rect 26240 21966 26292 21972
rect 27448 21690 27476 23054
rect 27528 22976 27580 22982
rect 27528 22918 27580 22924
rect 27540 22778 27568 22918
rect 27528 22772 27580 22778
rect 27528 22714 27580 22720
rect 27710 22536 27766 22545
rect 27710 22471 27712 22480
rect 27764 22471 27766 22480
rect 27712 22442 27764 22448
rect 27528 22432 27580 22438
rect 27528 22374 27580 22380
rect 27540 22030 27568 22374
rect 27528 22024 27580 22030
rect 27528 21966 27580 21972
rect 27712 21888 27764 21894
rect 27710 21856 27712 21865
rect 27764 21856 27766 21865
rect 27710 21791 27766 21800
rect 27436 21684 27488 21690
rect 27436 21626 27488 21632
rect 27804 21548 27856 21554
rect 27804 21490 27856 21496
rect 26056 21480 26108 21486
rect 26056 21422 26108 21428
rect 25872 21344 25924 21350
rect 25872 21286 25924 21292
rect 27620 21344 27672 21350
rect 27620 21286 27672 21292
rect 27632 21185 27660 21286
rect 27618 21176 27674 21185
rect 27618 21111 27674 21120
rect 26424 20800 26476 20806
rect 26424 20742 26476 20748
rect 26436 20534 26464 20742
rect 26424 20528 26476 20534
rect 26424 20470 26476 20476
rect 27816 20058 27844 21490
rect 27804 20052 27856 20058
rect 27804 19994 27856 20000
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 25792 12850 25820 14010
rect 27528 13932 27580 13938
rect 27528 13874 27580 13880
rect 27540 13705 27568 13874
rect 27526 13696 27582 13705
rect 27526 13631 27582 13640
rect 25780 12844 25832 12850
rect 25780 12786 25832 12792
rect 25228 11076 25280 11082
rect 25228 11018 25280 11024
rect 24952 9988 25004 9994
rect 24952 9930 25004 9936
rect 25136 9988 25188 9994
rect 25136 9930 25188 9936
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 24768 8832 24820 8838
rect 24768 8774 24820 8780
rect 24780 8634 24808 8774
rect 24676 8628 24728 8634
rect 24676 8570 24728 8576
rect 24768 8628 24820 8634
rect 24768 8570 24820 8576
rect 24688 8430 24716 8570
rect 25056 8566 25084 8910
rect 25044 8560 25096 8566
rect 25044 8502 25096 8508
rect 24676 8424 24728 8430
rect 24676 8366 24728 8372
rect 24676 8288 24728 8294
rect 24676 8230 24728 8236
rect 24688 7954 24716 8230
rect 25056 8090 25084 8502
rect 25148 8362 25176 9930
rect 25240 8498 25268 11018
rect 25320 11008 25372 11014
rect 25320 10950 25372 10956
rect 25332 10674 25360 10950
rect 25320 10668 25372 10674
rect 25320 10610 25372 10616
rect 25228 8492 25280 8498
rect 25228 8434 25280 8440
rect 27712 8492 27764 8498
rect 27712 8434 27764 8440
rect 25136 8356 25188 8362
rect 25136 8298 25188 8304
rect 25044 8084 25096 8090
rect 25044 8026 25096 8032
rect 24400 7948 24452 7954
rect 24400 7890 24452 7896
rect 24676 7948 24728 7954
rect 24676 7890 24728 7896
rect 24216 7404 24268 7410
rect 24216 7346 24268 7352
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 24124 7336 24176 7342
rect 24124 7278 24176 7284
rect 24032 7200 24084 7206
rect 24032 7142 24084 7148
rect 23480 6996 23532 7002
rect 23480 6938 23532 6944
rect 21548 6316 21600 6322
rect 21548 6258 21600 6264
rect 23020 6316 23072 6322
rect 23020 6258 23072 6264
rect 23032 6118 23060 6258
rect 24044 6254 24072 7142
rect 24320 7002 24348 7346
rect 24308 6996 24360 7002
rect 24308 6938 24360 6944
rect 24412 6866 24440 7890
rect 25148 7818 25176 8298
rect 25136 7812 25188 7818
rect 25136 7754 25188 7760
rect 24400 6860 24452 6866
rect 24400 6802 24452 6808
rect 25148 6730 25176 7754
rect 27620 7268 27672 7274
rect 27620 7210 27672 7216
rect 25136 6724 25188 6730
rect 25136 6666 25188 6672
rect 27632 6458 27660 7210
rect 27620 6452 27672 6458
rect 27620 6394 27672 6400
rect 24032 6248 24084 6254
rect 24032 6190 24084 6196
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 23020 6112 23072 6118
rect 23020 6054 23072 6060
rect 27724 5914 27752 8434
rect 27804 6316 27856 6322
rect 27804 6258 27856 6264
rect 27816 6225 27844 6258
rect 27802 6216 27858 6225
rect 27802 6151 27858 6160
rect 27712 5908 27764 5914
rect 27712 5850 27764 5856
rect 27528 5704 27580 5710
rect 27528 5646 27580 5652
rect 14372 5636 14424 5642
rect 14372 5578 14424 5584
rect 16764 5636 16816 5642
rect 16764 5578 16816 5584
rect 17868 5636 17920 5642
rect 17868 5578 17920 5584
rect 15660 5568 15712 5574
rect 27540 5545 27568 5646
rect 15660 5510 15712 5516
rect 27526 5536 27582 5545
rect 13268 5364 13320 5370
rect 13268 5306 13320 5312
rect 15672 5302 15700 5510
rect 27526 5471 27582 5480
rect 13084 5296 13136 5302
rect 13084 5238 13136 5244
rect 15660 5296 15712 5302
rect 15660 5238 15712 5244
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5828 800 5856 2382
rect 8404 800 8432 2382
rect 5814 0 5870 800
rect 8390 0 8446 800
<< via2 >>
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 846 24656 902 24712
rect 846 23976 902 24032
rect 846 23060 848 23080
rect 848 23060 900 23080
rect 900 23060 902 23080
rect 846 23024 902 23060
rect 1398 22480 1454 22536
rect 1306 21120 1362 21176
rect 1398 20440 1454 20496
rect 846 19896 902 19952
rect 2870 22344 2926 22400
rect 2778 22072 2834 22128
rect 1490 17720 1546 17776
rect 846 15816 902 15872
rect 1398 13640 1454 13696
rect 846 11756 902 11792
rect 846 11736 848 11756
rect 848 11736 900 11756
rect 900 11736 902 11756
rect 2870 21800 2926 21856
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 10322 27548 10324 27568
rect 10324 27548 10376 27568
rect 10376 27548 10378 27568
rect 10322 27512 10378 27548
rect 10782 27532 10838 27568
rect 10782 27512 10784 27532
rect 10784 27512 10836 27532
rect 10836 27512 10838 27532
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 11794 27512 11850 27568
rect 14646 27648 14702 27704
rect 18970 27376 19026 27432
rect 19338 26868 19340 26888
rect 19340 26868 19392 26888
rect 19392 26868 19394 26888
rect 19338 26832 19394 26868
rect 19522 27240 19578 27296
rect 19982 27548 19984 27568
rect 19984 27548 20036 27568
rect 20036 27548 20038 27568
rect 19982 27512 20038 27548
rect 20166 27376 20222 27432
rect 20258 27276 20260 27296
rect 20260 27276 20312 27296
rect 20312 27276 20314 27296
rect 20258 27240 20314 27276
rect 20074 26852 20130 26888
rect 20074 26832 20076 26852
rect 20076 26832 20128 26852
rect 20128 26832 20130 26852
rect 20994 27240 21050 27296
rect 13542 20304 13598 20360
rect 14002 20848 14058 20904
rect 13910 20440 13966 20496
rect 12162 17720 12218 17776
rect 10690 13912 10746 13968
rect 9770 12144 9826 12200
rect 10874 12008 10930 12064
rect 10230 11348 10286 11384
rect 10230 11328 10232 11348
rect 10232 11328 10284 11348
rect 10284 11328 10286 11348
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 10598 11192 10654 11248
rect 9586 9868 9588 9888
rect 9588 9868 9640 9888
rect 9640 9868 9642 9888
rect 9586 9832 9642 9868
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 11334 10920 11390 10976
rect 12898 17720 12954 17776
rect 11978 11756 12034 11792
rect 11978 11736 11980 11756
rect 11980 11736 12032 11756
rect 12032 11736 12034 11756
rect 11702 11600 11758 11656
rect 11610 11056 11666 11112
rect 11610 9968 11666 10024
rect 12254 11192 12310 11248
rect 14554 20440 14610 20496
rect 15106 20984 15162 21040
rect 15474 20304 15530 20360
rect 12438 12300 12494 12336
rect 12438 12280 12440 12300
rect 12440 12280 12492 12300
rect 12492 12280 12494 12300
rect 13358 12280 13414 12336
rect 11794 6976 11850 7032
rect 11426 6840 11482 6896
rect 11610 6432 11666 6488
rect 13082 10920 13138 10976
rect 12622 6860 12678 6896
rect 12622 6840 12624 6860
rect 12624 6840 12676 6860
rect 12676 6840 12678 6860
rect 12346 6568 12402 6624
rect 12346 6060 12348 6080
rect 12348 6060 12400 6080
rect 12400 6060 12402 6080
rect 12346 6024 12402 6060
rect 13082 6976 13138 7032
rect 13542 11736 13598 11792
rect 13358 9560 13414 9616
rect 13266 7928 13322 7984
rect 12898 6160 12954 6216
rect 14278 15020 14334 15056
rect 14278 15000 14280 15020
rect 14280 15000 14332 15020
rect 14332 15000 14334 15020
rect 22282 26560 22338 26616
rect 22650 27276 22652 27296
rect 22652 27276 22704 27296
rect 22704 27276 22706 27296
rect 22650 27240 22706 27276
rect 23110 27240 23166 27296
rect 22558 26696 22614 26752
rect 23018 26560 23074 26616
rect 16486 20868 16542 20904
rect 16486 20848 16488 20868
rect 16488 20848 16540 20868
rect 16540 20848 16542 20868
rect 14094 11056 14150 11112
rect 15198 13776 15254 13832
rect 15198 12724 15200 12744
rect 15200 12724 15252 12744
rect 15252 12724 15254 12744
rect 15198 12688 15254 12724
rect 14830 11056 14886 11112
rect 15566 11756 15622 11792
rect 15566 11736 15568 11756
rect 15568 11736 15620 11756
rect 15620 11736 15622 11756
rect 15566 11464 15622 11520
rect 13542 6976 13598 7032
rect 13634 6568 13690 6624
rect 13450 6432 13506 6488
rect 14738 6568 14794 6624
rect 16118 13912 16174 13968
rect 15842 11600 15898 11656
rect 16118 12008 16174 12064
rect 16670 15272 16726 15328
rect 16394 12008 16450 12064
rect 16210 11600 16266 11656
rect 16118 11464 16174 11520
rect 15750 9968 15806 10024
rect 16026 9832 16082 9888
rect 15842 8084 15898 8120
rect 15842 8064 15844 8084
rect 15844 8064 15896 8084
rect 15896 8064 15898 8084
rect 15658 6976 15714 7032
rect 15106 6704 15162 6760
rect 14646 6060 14648 6080
rect 14648 6060 14700 6080
rect 14700 6060 14702 6080
rect 14646 6024 14702 6060
rect 18418 22480 18474 22536
rect 16854 11076 16910 11112
rect 16854 11056 16856 11076
rect 16856 11056 16908 11076
rect 16908 11056 16910 11076
rect 17682 13776 17738 13832
rect 18694 22652 18696 22672
rect 18696 22652 18748 22672
rect 18748 22652 18750 22672
rect 18694 22616 18750 22652
rect 18970 22636 19026 22672
rect 18970 22616 18972 22636
rect 18972 22616 19024 22636
rect 19024 22616 19026 22636
rect 17222 12008 17278 12064
rect 16762 9832 16818 9888
rect 16578 9560 16634 9616
rect 17038 6740 17040 6760
rect 17040 6740 17092 6760
rect 17092 6740 17094 6760
rect 17038 6704 17094 6740
rect 17774 11056 17830 11112
rect 18050 12180 18052 12200
rect 18052 12180 18104 12200
rect 18104 12180 18106 12200
rect 18050 12144 18106 12180
rect 18050 11092 18052 11112
rect 18052 11092 18104 11112
rect 18104 11092 18106 11112
rect 18050 11056 18106 11092
rect 21270 24148 21272 24168
rect 21272 24148 21324 24168
rect 21324 24148 21326 24168
rect 21270 24112 21326 24148
rect 23570 26288 23626 26344
rect 19246 22480 19302 22536
rect 18234 12144 18290 12200
rect 19890 21020 19892 21040
rect 19892 21020 19944 21040
rect 19944 21020 19946 21040
rect 19890 20984 19946 21020
rect 20442 21020 20444 21040
rect 20444 21020 20496 21040
rect 20496 21020 20498 21040
rect 20442 20984 20498 21020
rect 20534 20304 20590 20360
rect 19798 19760 19854 19816
rect 18786 12688 18842 12744
rect 18510 12144 18566 12200
rect 18510 11328 18566 11384
rect 20626 20204 20628 20224
rect 20628 20204 20680 20224
rect 20680 20204 20682 20224
rect 20626 20168 20682 20204
rect 21362 20304 21418 20360
rect 21638 20168 21694 20224
rect 20902 19352 20958 19408
rect 19338 12300 19394 12336
rect 19338 12280 19340 12300
rect 19340 12280 19392 12300
rect 19392 12280 19394 12300
rect 21638 19508 21694 19544
rect 21638 19488 21640 19508
rect 21640 19488 21692 19508
rect 21692 19488 21694 19508
rect 20718 16496 20774 16552
rect 19982 13776 20038 13832
rect 19982 13232 20038 13288
rect 20534 12300 20590 12336
rect 20534 12280 20536 12300
rect 20536 12280 20588 12300
rect 20588 12280 20590 12300
rect 22374 19796 22376 19816
rect 22376 19796 22428 19816
rect 22428 19796 22430 19816
rect 22374 19760 22430 19796
rect 24306 26732 24308 26752
rect 24308 26732 24360 26752
rect 24360 26732 24362 26752
rect 24306 26696 24362 26732
rect 22926 24112 22982 24168
rect 22558 19488 22614 19544
rect 21454 16516 21510 16552
rect 21454 16496 21456 16516
rect 21456 16496 21508 16516
rect 21508 16496 21510 16516
rect 22098 13640 22154 13696
rect 21822 13096 21878 13152
rect 18142 7828 18144 7848
rect 18144 7828 18196 7848
rect 18196 7828 18198 7848
rect 18142 7792 18198 7828
rect 17958 7404 18014 7440
rect 17958 7384 17960 7404
rect 17960 7384 18012 7404
rect 18012 7384 18014 7404
rect 18326 7384 18382 7440
rect 22282 13640 22338 13696
rect 22190 13096 22246 13152
rect 21362 11056 21418 11112
rect 20350 7404 20406 7440
rect 20534 7656 20590 7712
rect 20350 7384 20352 7404
rect 20352 7384 20404 7404
rect 20404 7384 20406 7404
rect 17682 6196 17684 6216
rect 17684 6196 17736 6216
rect 17736 6196 17738 6216
rect 17682 6160 17738 6196
rect 18694 6704 18750 6760
rect 20810 7828 20812 7848
rect 20812 7828 20864 7848
rect 20864 7828 20866 7848
rect 20810 7792 20866 7828
rect 21086 7540 21142 7576
rect 21086 7520 21088 7540
rect 21088 7520 21140 7540
rect 21140 7520 21142 7540
rect 21270 7792 21326 7848
rect 21178 7384 21234 7440
rect 22650 14184 22706 14240
rect 21914 7656 21970 7712
rect 27710 26560 27766 26616
rect 27342 26288 27398 26344
rect 27526 25880 27582 25936
rect 23110 15544 23166 15600
rect 25134 14184 25190 14240
rect 23754 7928 23810 7984
rect 27710 25200 27766 25256
rect 27710 24556 27712 24576
rect 27712 24556 27764 24576
rect 27764 24556 27766 24576
rect 27710 24520 27766 24556
rect 27710 23840 27766 23896
rect 27526 23160 27582 23216
rect 27710 22500 27766 22536
rect 27710 22480 27712 22500
rect 27712 22480 27764 22500
rect 27764 22480 27766 22500
rect 27710 21836 27712 21856
rect 27712 21836 27764 21856
rect 27764 21836 27766 21856
rect 27710 21800 27766 21836
rect 27618 21120 27674 21176
rect 27526 13640 27582 13696
rect 27802 6160 27858 6216
rect 27526 5480 27582 5536
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 14641 27706 14707 27709
rect 14641 27704 19442 27706
rect 14641 27648 14646 27704
rect 14702 27648 19442 27704
rect 14641 27646 19442 27648
rect 14641 27643 14707 27646
rect 10317 27570 10383 27573
rect 10777 27570 10843 27573
rect 11789 27570 11855 27573
rect 10317 27568 11855 27570
rect 10317 27512 10322 27568
rect 10378 27512 10782 27568
rect 10838 27512 11794 27568
rect 11850 27512 11855 27568
rect 10317 27510 11855 27512
rect 19382 27570 19442 27646
rect 19977 27570 20043 27573
rect 19382 27568 20043 27570
rect 19382 27512 19982 27568
rect 20038 27512 20043 27568
rect 19382 27510 20043 27512
rect 10317 27507 10383 27510
rect 10777 27507 10843 27510
rect 11789 27507 11855 27510
rect 19977 27507 20043 27510
rect 18965 27434 19031 27437
rect 20161 27434 20227 27437
rect 18965 27432 20227 27434
rect 18965 27376 18970 27432
rect 19026 27376 20166 27432
rect 20222 27376 20227 27432
rect 18965 27374 20227 27376
rect 18965 27371 19031 27374
rect 20161 27371 20227 27374
rect 19517 27298 19583 27301
rect 20253 27298 20319 27301
rect 20989 27298 21055 27301
rect 19517 27296 21055 27298
rect 19517 27240 19522 27296
rect 19578 27240 20258 27296
rect 20314 27240 20994 27296
rect 21050 27240 21055 27296
rect 19517 27238 21055 27240
rect 19517 27235 19583 27238
rect 20253 27235 20319 27238
rect 20989 27235 21055 27238
rect 22645 27298 22711 27301
rect 23105 27298 23171 27301
rect 22645 27296 23171 27298
rect 22645 27240 22650 27296
rect 22706 27240 23110 27296
rect 23166 27240 23171 27296
rect 22645 27238 23171 27240
rect 22645 27235 22711 27238
rect 23105 27235 23171 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 19333 26890 19399 26893
rect 20069 26890 20135 26893
rect 19333 26888 20135 26890
rect 19333 26832 19338 26888
rect 19394 26832 20074 26888
rect 20130 26832 20135 26888
rect 19333 26830 20135 26832
rect 19333 26827 19399 26830
rect 20069 26827 20135 26830
rect 22553 26754 22619 26757
rect 24301 26754 24367 26757
rect 22553 26752 24367 26754
rect 22553 26696 22558 26752
rect 22614 26696 24306 26752
rect 24362 26696 24367 26752
rect 22553 26694 24367 26696
rect 22553 26691 22619 26694
rect 24301 26691 24367 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 22277 26618 22343 26621
rect 23013 26618 23079 26621
rect 22277 26616 23079 26618
rect 22277 26560 22282 26616
rect 22338 26560 23018 26616
rect 23074 26560 23079 26616
rect 22277 26558 23079 26560
rect 22277 26555 22343 26558
rect 23013 26555 23079 26558
rect 27705 26618 27771 26621
rect 28532 26618 29332 26648
rect 27705 26616 29332 26618
rect 27705 26560 27710 26616
rect 27766 26560 29332 26616
rect 27705 26558 29332 26560
rect 27705 26555 27771 26558
rect 28532 26528 29332 26558
rect 23565 26346 23631 26349
rect 27337 26346 27403 26349
rect 23565 26344 27403 26346
rect 23565 26288 23570 26344
rect 23626 26288 27342 26344
rect 27398 26288 27403 26344
rect 23565 26286 27403 26288
rect 23565 26283 23631 26286
rect 27337 26283 27403 26286
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 27521 25938 27587 25941
rect 28532 25938 29332 25968
rect 27521 25936 29332 25938
rect 27521 25880 27526 25936
rect 27582 25880 29332 25936
rect 27521 25878 29332 25880
rect 27521 25875 27587 25878
rect 28532 25848 29332 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 27705 25258 27771 25261
rect 28532 25258 29332 25288
rect 27705 25256 29332 25258
rect 27705 25200 27710 25256
rect 27766 25200 29332 25256
rect 27705 25198 29332 25200
rect 27705 25195 27771 25198
rect 28532 25168 29332 25198
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 841 24714 907 24717
rect 798 24712 907 24714
rect 798 24656 846 24712
rect 902 24656 907 24712
rect 798 24651 907 24656
rect 798 24608 858 24651
rect 0 24518 858 24608
rect 27705 24578 27771 24581
rect 28532 24578 29332 24608
rect 27705 24576 29332 24578
rect 27705 24520 27710 24576
rect 27766 24520 29332 24576
rect 27705 24518 29332 24520
rect 0 24488 800 24518
rect 27705 24515 27771 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 28532 24488 29332 24518
rect 4210 24447 4526 24448
rect 21265 24170 21331 24173
rect 22921 24170 22987 24173
rect 21265 24168 22987 24170
rect 21265 24112 21270 24168
rect 21326 24112 22926 24168
rect 22982 24112 22987 24168
rect 21265 24110 22987 24112
rect 21265 24107 21331 24110
rect 22921 24107 22987 24110
rect 841 24034 907 24037
rect 798 24032 907 24034
rect 798 23976 846 24032
rect 902 23976 907 24032
rect 798 23971 907 23976
rect 798 23928 858 23971
rect 0 23838 858 23928
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 27705 23898 27771 23901
rect 28532 23898 29332 23928
rect 27705 23896 29332 23898
rect 27705 23840 27710 23896
rect 27766 23840 29332 23896
rect 27705 23838 29332 23840
rect 0 23808 800 23838
rect 27705 23835 27771 23838
rect 28532 23808 29332 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 0 23218 800 23248
rect 27521 23218 27587 23221
rect 28532 23218 29332 23248
rect 0 23128 858 23218
rect 27521 23216 29332 23218
rect 27521 23160 27526 23216
rect 27582 23160 29332 23216
rect 27521 23158 29332 23160
rect 27521 23155 27587 23158
rect 28532 23128 29332 23158
rect 798 23085 858 23128
rect 798 23080 907 23085
rect 798 23024 846 23080
rect 902 23024 907 23080
rect 798 23022 907 23024
rect 841 23019 907 23022
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 18689 22674 18755 22677
rect 18965 22674 19031 22677
rect 18689 22672 19031 22674
rect 18689 22616 18694 22672
rect 18750 22616 18970 22672
rect 19026 22616 19031 22672
rect 18689 22614 19031 22616
rect 18689 22611 18755 22614
rect 18965 22611 19031 22614
rect 0 22538 800 22568
rect 1393 22538 1459 22541
rect 0 22536 1459 22538
rect 0 22480 1398 22536
rect 1454 22480 1459 22536
rect 0 22478 1459 22480
rect 0 22448 800 22478
rect 1393 22475 1459 22478
rect 18413 22538 18479 22541
rect 19241 22538 19307 22541
rect 18413 22536 19307 22538
rect 18413 22480 18418 22536
rect 18474 22480 19246 22536
rect 19302 22480 19307 22536
rect 18413 22478 19307 22480
rect 18413 22475 18479 22478
rect 19241 22475 19307 22478
rect 27705 22538 27771 22541
rect 28532 22538 29332 22568
rect 27705 22536 29332 22538
rect 27705 22480 27710 22536
rect 27766 22480 29332 22536
rect 27705 22478 29332 22480
rect 27705 22475 27771 22478
rect 28532 22448 29332 22478
rect 2865 22402 2931 22405
rect 2822 22400 2931 22402
rect 2822 22344 2870 22400
rect 2926 22344 2931 22400
rect 2822 22339 2931 22344
rect 2822 22133 2882 22339
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 2773 22128 2882 22133
rect 2773 22072 2778 22128
rect 2834 22072 2882 22128
rect 2773 22070 2882 22072
rect 2773 22067 2839 22070
rect 0 21858 800 21888
rect 2865 21858 2931 21861
rect 0 21856 2931 21858
rect 0 21800 2870 21856
rect 2926 21800 2931 21856
rect 0 21798 2931 21800
rect 0 21768 800 21798
rect 2865 21795 2931 21798
rect 27705 21858 27771 21861
rect 28532 21858 29332 21888
rect 27705 21856 29332 21858
rect 27705 21800 27710 21856
rect 27766 21800 29332 21856
rect 27705 21798 29332 21800
rect 27705 21795 27771 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 28532 21768 29332 21798
rect 4870 21727 5186 21728
rect 4210 21248 4526 21249
rect 0 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 1301 21178 1367 21181
rect 0 21176 1367 21178
rect 0 21120 1306 21176
rect 1362 21120 1367 21176
rect 0 21118 1367 21120
rect 0 21088 800 21118
rect 1301 21115 1367 21118
rect 27613 21178 27679 21181
rect 28532 21178 29332 21208
rect 27613 21176 29332 21178
rect 27613 21120 27618 21176
rect 27674 21120 29332 21176
rect 27613 21118 29332 21120
rect 27613 21115 27679 21118
rect 28532 21088 29332 21118
rect 15101 21042 15167 21045
rect 19885 21042 19951 21045
rect 20437 21042 20503 21045
rect 15101 21040 20503 21042
rect 15101 20984 15106 21040
rect 15162 20984 19890 21040
rect 19946 20984 20442 21040
rect 20498 20984 20503 21040
rect 15101 20982 20503 20984
rect 15101 20979 15167 20982
rect 19885 20979 19951 20982
rect 20437 20979 20503 20982
rect 13997 20906 14063 20909
rect 16481 20906 16547 20909
rect 13997 20904 16547 20906
rect 13997 20848 14002 20904
rect 14058 20848 16486 20904
rect 16542 20848 16547 20904
rect 13997 20846 16547 20848
rect 13997 20843 14063 20846
rect 16481 20843 16547 20846
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 0 20498 800 20528
rect 1393 20498 1459 20501
rect 0 20496 1459 20498
rect 0 20440 1398 20496
rect 1454 20440 1459 20496
rect 0 20438 1459 20440
rect 0 20408 800 20438
rect 1393 20435 1459 20438
rect 13905 20498 13971 20501
rect 14549 20498 14615 20501
rect 13905 20496 14615 20498
rect 13905 20440 13910 20496
rect 13966 20440 14554 20496
rect 14610 20440 14615 20496
rect 13905 20438 14615 20440
rect 13905 20435 13971 20438
rect 14549 20435 14615 20438
rect 13537 20362 13603 20365
rect 15469 20362 15535 20365
rect 13537 20360 15535 20362
rect 13537 20304 13542 20360
rect 13598 20304 15474 20360
rect 15530 20304 15535 20360
rect 13537 20302 15535 20304
rect 13537 20299 13603 20302
rect 15469 20299 15535 20302
rect 20529 20362 20595 20365
rect 21357 20362 21423 20365
rect 22502 20362 22508 20364
rect 20529 20360 22508 20362
rect 20529 20304 20534 20360
rect 20590 20304 21362 20360
rect 21418 20304 22508 20360
rect 20529 20302 22508 20304
rect 20529 20299 20595 20302
rect 21357 20299 21423 20302
rect 22502 20300 22508 20302
rect 22572 20300 22578 20364
rect 20621 20226 20687 20229
rect 21633 20226 21699 20229
rect 20621 20224 21699 20226
rect 20621 20168 20626 20224
rect 20682 20168 21638 20224
rect 21694 20168 21699 20224
rect 20621 20166 21699 20168
rect 20621 20163 20687 20166
rect 21633 20163 21699 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 841 19954 907 19957
rect 798 19952 907 19954
rect 798 19896 846 19952
rect 902 19896 907 19952
rect 798 19891 907 19896
rect 798 19848 858 19891
rect 0 19758 858 19848
rect 19793 19818 19859 19821
rect 22369 19818 22435 19821
rect 23054 19818 23060 19820
rect 19793 19816 23060 19818
rect 19793 19760 19798 19816
rect 19854 19760 22374 19816
rect 22430 19760 23060 19816
rect 19793 19758 23060 19760
rect 0 19728 800 19758
rect 19793 19755 19859 19758
rect 22369 19755 22435 19758
rect 23054 19756 23060 19758
rect 23124 19756 23130 19820
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 21633 19546 21699 19549
rect 22553 19546 22619 19549
rect 21633 19544 22619 19546
rect 21633 19488 21638 19544
rect 21694 19488 22558 19544
rect 22614 19488 22619 19544
rect 21633 19486 22619 19488
rect 21633 19483 21699 19486
rect 22553 19483 22619 19486
rect 20662 19348 20668 19412
rect 20732 19410 20738 19412
rect 20897 19410 20963 19413
rect 20732 19408 20963 19410
rect 20732 19352 20902 19408
rect 20958 19352 20963 19408
rect 20732 19350 20963 19352
rect 20732 19348 20738 19350
rect 20897 19347 20963 19350
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 0 17778 800 17808
rect 1485 17778 1551 17781
rect 0 17776 1551 17778
rect 0 17720 1490 17776
rect 1546 17720 1551 17776
rect 0 17718 1551 17720
rect 0 17688 800 17718
rect 1485 17715 1551 17718
rect 12157 17778 12223 17781
rect 12893 17778 12959 17781
rect 12157 17776 12959 17778
rect 12157 17720 12162 17776
rect 12218 17720 12898 17776
rect 12954 17720 12959 17776
rect 12157 17718 12959 17720
rect 12157 17715 12223 17718
rect 12893 17715 12959 17718
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 20713 16554 20779 16557
rect 21449 16554 21515 16557
rect 20713 16552 21515 16554
rect 20713 16496 20718 16552
rect 20774 16496 21454 16552
rect 21510 16496 21515 16552
rect 20713 16494 21515 16496
rect 20713 16491 20779 16494
rect 21449 16491 21515 16494
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 841 15874 907 15877
rect 798 15872 907 15874
rect 798 15816 846 15872
rect 902 15816 907 15872
rect 798 15811 907 15816
rect 798 15768 858 15811
rect 0 15678 858 15768
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 0 15648 800 15678
rect 23105 15604 23171 15605
rect 23054 15540 23060 15604
rect 23124 15602 23171 15604
rect 23124 15600 23216 15602
rect 23166 15544 23216 15600
rect 23124 15542 23216 15544
rect 23124 15540 23171 15542
rect 23105 15539 23171 15540
rect 16665 15332 16731 15333
rect 16614 15330 16620 15332
rect 16574 15270 16620 15330
rect 16684 15328 16731 15332
rect 16726 15272 16731 15328
rect 16614 15268 16620 15270
rect 16684 15268 16731 15272
rect 16665 15267 16731 15268
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 14273 15058 14339 15061
rect 20662 15058 20668 15060
rect 14273 15056 20668 15058
rect 14273 15000 14278 15056
rect 14334 15000 20668 15056
rect 14273 14998 20668 15000
rect 14273 14995 14339 14998
rect 20662 14996 20668 14998
rect 20732 14996 20738 15060
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 22502 14180 22508 14244
rect 22572 14242 22578 14244
rect 22645 14242 22711 14245
rect 25129 14242 25195 14245
rect 22572 14240 25195 14242
rect 22572 14184 22650 14240
rect 22706 14184 25134 14240
rect 25190 14184 25195 14240
rect 22572 14182 25195 14184
rect 22572 14180 22578 14182
rect 22645 14179 22711 14182
rect 25129 14179 25195 14182
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 10685 13970 10751 13973
rect 16113 13970 16179 13973
rect 10685 13968 16179 13970
rect 10685 13912 10690 13968
rect 10746 13912 16118 13968
rect 16174 13912 16179 13968
rect 10685 13910 16179 13912
rect 10685 13907 10751 13910
rect 16113 13907 16179 13910
rect 15193 13834 15259 13837
rect 15326 13834 15332 13836
rect 15193 13832 15332 13834
rect 15193 13776 15198 13832
rect 15254 13776 15332 13832
rect 15193 13774 15332 13776
rect 15193 13771 15259 13774
rect 15326 13772 15332 13774
rect 15396 13772 15402 13836
rect 17677 13834 17743 13837
rect 17902 13834 17908 13836
rect 17677 13832 17908 13834
rect 17677 13776 17682 13832
rect 17738 13776 17908 13832
rect 17677 13774 17908 13776
rect 17677 13771 17743 13774
rect 17902 13772 17908 13774
rect 17972 13772 17978 13836
rect 19977 13834 20043 13837
rect 20110 13834 20116 13836
rect 19977 13832 20116 13834
rect 19977 13776 19982 13832
rect 20038 13776 20116 13832
rect 19977 13774 20116 13776
rect 19977 13771 20043 13774
rect 20110 13772 20116 13774
rect 20180 13772 20186 13836
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 22093 13698 22159 13701
rect 22277 13698 22343 13701
rect 22093 13696 22343 13698
rect 22093 13640 22098 13696
rect 22154 13640 22282 13696
rect 22338 13640 22343 13696
rect 22093 13638 22343 13640
rect 22093 13635 22159 13638
rect 22277 13635 22343 13638
rect 27521 13698 27587 13701
rect 28532 13698 29332 13728
rect 27521 13696 29332 13698
rect 27521 13640 27526 13696
rect 27582 13640 29332 13696
rect 27521 13638 29332 13640
rect 27521 13635 27587 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 28532 13608 29332 13638
rect 4210 13567 4526 13568
rect 19977 13292 20043 13293
rect 19926 13290 19932 13292
rect 19886 13230 19932 13290
rect 19996 13288 20043 13292
rect 20038 13232 20043 13288
rect 19926 13228 19932 13230
rect 19996 13228 20043 13232
rect 19977 13227 20043 13228
rect 21817 13154 21883 13157
rect 22185 13154 22251 13157
rect 21817 13152 22251 13154
rect 21817 13096 21822 13152
rect 21878 13096 22190 13152
rect 22246 13096 22251 13152
rect 21817 13094 22251 13096
rect 21817 13091 21883 13094
rect 22185 13091 22251 13094
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 15193 12746 15259 12749
rect 18781 12746 18847 12749
rect 15193 12744 18847 12746
rect 15193 12688 15198 12744
rect 15254 12688 18786 12744
rect 18842 12688 18847 12744
rect 15193 12686 18847 12688
rect 15193 12683 15259 12686
rect 18781 12683 18847 12686
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 12433 12338 12499 12341
rect 13353 12338 13419 12341
rect 12433 12336 13419 12338
rect 12433 12280 12438 12336
rect 12494 12280 13358 12336
rect 13414 12280 13419 12336
rect 12433 12278 13419 12280
rect 12433 12275 12499 12278
rect 13353 12275 13419 12278
rect 19333 12338 19399 12341
rect 20529 12338 20595 12341
rect 19333 12336 20595 12338
rect 19333 12280 19338 12336
rect 19394 12280 20534 12336
rect 20590 12280 20595 12336
rect 19333 12278 20595 12280
rect 19333 12275 19399 12278
rect 20529 12275 20595 12278
rect 9765 12202 9831 12205
rect 18045 12202 18111 12205
rect 9765 12200 18111 12202
rect 9765 12144 9770 12200
rect 9826 12144 18050 12200
rect 18106 12144 18111 12200
rect 9765 12142 18111 12144
rect 9765 12139 9831 12142
rect 18045 12139 18111 12142
rect 18229 12202 18295 12205
rect 18505 12202 18571 12205
rect 18229 12200 18571 12202
rect 18229 12144 18234 12200
rect 18290 12144 18510 12200
rect 18566 12144 18571 12200
rect 18229 12142 18571 12144
rect 18229 12139 18295 12142
rect 18505 12139 18571 12142
rect 10869 12066 10935 12069
rect 16113 12066 16179 12069
rect 16389 12066 16455 12069
rect 17217 12066 17283 12069
rect 10869 12064 17283 12066
rect 10869 12008 10874 12064
rect 10930 12008 16118 12064
rect 16174 12008 16394 12064
rect 16450 12008 17222 12064
rect 17278 12008 17283 12064
rect 10869 12006 17283 12008
rect 10869 12003 10935 12006
rect 16113 12003 16179 12006
rect 16389 12003 16455 12006
rect 17217 12003 17283 12006
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 841 11794 907 11797
rect 798 11792 907 11794
rect 798 11736 846 11792
rect 902 11736 907 11792
rect 798 11731 907 11736
rect 11973 11794 12039 11797
rect 13537 11794 13603 11797
rect 15561 11794 15627 11797
rect 11973 11792 15627 11794
rect 11973 11736 11978 11792
rect 12034 11736 13542 11792
rect 13598 11736 15566 11792
rect 15622 11736 15627 11792
rect 11973 11734 15627 11736
rect 11973 11731 12039 11734
rect 13537 11731 13603 11734
rect 15561 11731 15627 11734
rect 798 11688 858 11731
rect 0 11598 858 11688
rect 11697 11658 11763 11661
rect 15837 11658 15903 11661
rect 16205 11658 16271 11661
rect 11697 11656 16271 11658
rect 11697 11600 11702 11656
rect 11758 11600 15842 11656
rect 15898 11600 16210 11656
rect 16266 11600 16271 11656
rect 11697 11598 16271 11600
rect 0 11568 800 11598
rect 11697 11595 11763 11598
rect 15837 11595 15903 11598
rect 16205 11595 16271 11598
rect 15561 11522 15627 11525
rect 16113 11522 16179 11525
rect 15561 11520 16179 11522
rect 15561 11464 15566 11520
rect 15622 11464 16118 11520
rect 16174 11464 16179 11520
rect 15561 11462 16179 11464
rect 15561 11459 15627 11462
rect 16113 11459 16179 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 10225 11386 10291 11389
rect 18505 11386 18571 11389
rect 10225 11384 18571 11386
rect 10225 11328 10230 11384
rect 10286 11328 18510 11384
rect 18566 11328 18571 11384
rect 10225 11326 18571 11328
rect 10225 11323 10291 11326
rect 18505 11323 18571 11326
rect 10593 11250 10659 11253
rect 12249 11250 12315 11253
rect 10593 11248 12315 11250
rect 10593 11192 10598 11248
rect 10654 11192 12254 11248
rect 12310 11192 12315 11248
rect 10593 11190 12315 11192
rect 10593 11187 10659 11190
rect 12249 11187 12315 11190
rect 11605 11114 11671 11117
rect 14089 11114 14155 11117
rect 11605 11112 14155 11114
rect 11605 11056 11610 11112
rect 11666 11056 14094 11112
rect 14150 11056 14155 11112
rect 11605 11054 14155 11056
rect 11605 11051 11671 11054
rect 14089 11051 14155 11054
rect 14825 11114 14891 11117
rect 16849 11114 16915 11117
rect 17769 11114 17835 11117
rect 14825 11112 17835 11114
rect 14825 11056 14830 11112
rect 14886 11056 16854 11112
rect 16910 11056 17774 11112
rect 17830 11056 17835 11112
rect 14825 11054 17835 11056
rect 14825 11051 14891 11054
rect 16849 11051 16915 11054
rect 17769 11051 17835 11054
rect 18045 11114 18111 11117
rect 21357 11114 21423 11117
rect 18045 11112 21423 11114
rect 18045 11056 18050 11112
rect 18106 11056 21362 11112
rect 21418 11056 21423 11112
rect 18045 11054 21423 11056
rect 18045 11051 18111 11054
rect 21357 11051 21423 11054
rect 11329 10978 11395 10981
rect 13077 10978 13143 10981
rect 11329 10976 13143 10978
rect 11329 10920 11334 10976
rect 11390 10920 13082 10976
rect 13138 10920 13143 10976
rect 11329 10918 13143 10920
rect 11329 10915 11395 10918
rect 13077 10915 13143 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 11605 10026 11671 10029
rect 15745 10026 15811 10029
rect 11605 10024 15811 10026
rect 11605 9968 11610 10024
rect 11666 9968 15750 10024
rect 15806 9968 15811 10024
rect 11605 9966 15811 9968
rect 11605 9963 11671 9966
rect 15745 9963 15811 9966
rect 9581 9890 9647 9893
rect 16021 9890 16087 9893
rect 16757 9890 16823 9893
rect 9581 9888 16823 9890
rect 9581 9832 9586 9888
rect 9642 9832 16026 9888
rect 16082 9832 16762 9888
rect 16818 9832 16823 9888
rect 9581 9830 16823 9832
rect 9581 9827 9647 9830
rect 16021 9827 16087 9830
rect 16757 9827 16823 9830
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 13353 9618 13419 9621
rect 16573 9618 16639 9621
rect 13353 9616 16639 9618
rect 13353 9560 13358 9616
rect 13414 9560 16578 9616
rect 16634 9560 16639 9616
rect 13353 9558 16639 9560
rect 13353 9555 13419 9558
rect 16573 9555 16639 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 15837 8122 15903 8125
rect 16614 8122 16620 8124
rect 15837 8120 16620 8122
rect 15837 8064 15842 8120
rect 15898 8064 16620 8120
rect 15837 8062 16620 8064
rect 15837 8059 15903 8062
rect 16614 8060 16620 8062
rect 16684 8060 16690 8124
rect 13261 7986 13327 7989
rect 23749 7986 23815 7989
rect 13261 7984 23815 7986
rect 13261 7928 13266 7984
rect 13322 7928 23754 7984
rect 23810 7928 23815 7984
rect 13261 7926 23815 7928
rect 13261 7923 13327 7926
rect 23749 7923 23815 7926
rect 18137 7850 18203 7853
rect 20805 7850 20871 7853
rect 21265 7850 21331 7853
rect 18137 7848 21331 7850
rect 18137 7792 18142 7848
rect 18198 7792 20810 7848
rect 20866 7792 21270 7848
rect 21326 7792 21331 7848
rect 18137 7790 21331 7792
rect 18137 7787 18203 7790
rect 20805 7787 20871 7790
rect 21265 7787 21331 7790
rect 20529 7714 20595 7717
rect 21909 7714 21975 7717
rect 20529 7712 21975 7714
rect 20529 7656 20534 7712
rect 20590 7656 21914 7712
rect 21970 7656 21975 7712
rect 20529 7654 21975 7656
rect 20529 7651 20595 7654
rect 21909 7651 21975 7654
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 17902 7516 17908 7580
rect 17972 7578 17978 7580
rect 21081 7578 21147 7581
rect 17972 7576 21147 7578
rect 17972 7520 21086 7576
rect 21142 7520 21147 7576
rect 17972 7518 21147 7520
rect 17972 7516 17978 7518
rect 21081 7515 21147 7518
rect 17953 7442 18019 7445
rect 18321 7442 18387 7445
rect 19926 7442 19932 7444
rect 17953 7440 19932 7442
rect 17953 7384 17958 7440
rect 18014 7384 18326 7440
rect 18382 7384 19932 7440
rect 17953 7382 19932 7384
rect 17953 7379 18019 7382
rect 18321 7379 18387 7382
rect 19926 7380 19932 7382
rect 19996 7380 20002 7444
rect 20345 7442 20411 7445
rect 21173 7442 21239 7445
rect 20345 7440 21239 7442
rect 20345 7384 20350 7440
rect 20406 7384 21178 7440
rect 21234 7384 21239 7440
rect 20345 7382 21239 7384
rect 20345 7379 20411 7382
rect 21173 7379 21239 7382
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 11789 7034 11855 7037
rect 13077 7034 13143 7037
rect 13537 7034 13603 7037
rect 15653 7034 15719 7037
rect 11789 7032 15719 7034
rect 11789 6976 11794 7032
rect 11850 6976 13082 7032
rect 13138 6976 13542 7032
rect 13598 6976 15658 7032
rect 15714 6976 15719 7032
rect 11789 6974 15719 6976
rect 11789 6971 11855 6974
rect 13077 6971 13143 6974
rect 13537 6971 13603 6974
rect 15653 6971 15719 6974
rect 11421 6898 11487 6901
rect 12617 6898 12683 6901
rect 11421 6896 12683 6898
rect 11421 6840 11426 6896
rect 11482 6840 12622 6896
rect 12678 6840 12683 6896
rect 11421 6838 12683 6840
rect 11421 6835 11487 6838
rect 12617 6835 12683 6838
rect 15101 6762 15167 6765
rect 15326 6762 15332 6764
rect 15101 6760 15332 6762
rect 15101 6704 15106 6760
rect 15162 6704 15332 6760
rect 15101 6702 15332 6704
rect 15101 6699 15167 6702
rect 15326 6700 15332 6702
rect 15396 6700 15402 6764
rect 17033 6762 17099 6765
rect 18689 6762 18755 6765
rect 15518 6760 18755 6762
rect 15518 6704 17038 6760
rect 17094 6704 18694 6760
rect 18750 6704 18755 6760
rect 15518 6702 18755 6704
rect 12341 6626 12407 6629
rect 13629 6626 13695 6629
rect 12341 6624 13695 6626
rect 12341 6568 12346 6624
rect 12402 6568 13634 6624
rect 13690 6568 13695 6624
rect 12341 6566 13695 6568
rect 12341 6563 12407 6566
rect 13629 6563 13695 6566
rect 14733 6626 14799 6629
rect 15518 6626 15578 6702
rect 17033 6699 17099 6702
rect 18689 6699 18755 6702
rect 14733 6624 15578 6626
rect 14733 6568 14738 6624
rect 14794 6568 15578 6624
rect 14733 6566 15578 6568
rect 14733 6563 14799 6566
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 11605 6490 11671 6493
rect 13445 6490 13511 6493
rect 11605 6488 13511 6490
rect 11605 6432 11610 6488
rect 11666 6432 13450 6488
rect 13506 6432 13511 6488
rect 11605 6430 13511 6432
rect 11605 6427 11671 6430
rect 13445 6427 13511 6430
rect 12893 6218 12959 6221
rect 17677 6218 17743 6221
rect 12893 6216 17743 6218
rect 12893 6160 12898 6216
rect 12954 6160 17682 6216
rect 17738 6160 17743 6216
rect 12893 6158 17743 6160
rect 12893 6155 12959 6158
rect 17677 6155 17743 6158
rect 27797 6218 27863 6221
rect 28532 6218 29332 6248
rect 27797 6216 29332 6218
rect 27797 6160 27802 6216
rect 27858 6160 29332 6216
rect 27797 6158 29332 6160
rect 27797 6155 27863 6158
rect 28532 6128 29332 6158
rect 12341 6082 12407 6085
rect 14641 6082 14707 6085
rect 12341 6080 14707 6082
rect 12341 6024 12346 6080
rect 12402 6024 14646 6080
rect 14702 6024 14707 6080
rect 12341 6022 14707 6024
rect 12341 6019 12407 6022
rect 14641 6019 14707 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 27521 5538 27587 5541
rect 28532 5538 29332 5568
rect 27521 5536 29332 5538
rect 27521 5480 27526 5536
rect 27582 5480 29332 5536
rect 27521 5478 29332 5480
rect 27521 5475 27587 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 28532 5448 29332 5478
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 20110 4796 20116 4860
rect 20180 4858 20186 4860
rect 28532 4858 29332 4888
rect 20180 4798 29332 4858
rect 20180 4796 20186 4798
rect 28532 4768 29332 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 22508 20300 22572 20364
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 23060 19756 23124 19820
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 20668 19348 20732 19412
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 23060 15600 23124 15604
rect 23060 15544 23110 15600
rect 23110 15544 23124 15600
rect 23060 15540 23124 15544
rect 16620 15328 16684 15332
rect 16620 15272 16670 15328
rect 16670 15272 16684 15328
rect 16620 15268 16684 15272
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 20668 14996 20732 15060
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 22508 14180 22572 14244
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 15332 13772 15396 13836
rect 17908 13772 17972 13836
rect 20116 13772 20180 13836
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 19932 13288 19996 13292
rect 19932 13232 19982 13288
rect 19982 13232 19996 13288
rect 19932 13228 19996 13232
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 16620 8060 16684 8124
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 17908 7516 17972 7580
rect 19932 7380 19996 7444
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 15332 6700 15396 6764
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 20116 4796 20180 4860
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 28864 4528 28880
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 28320 5188 28880
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 22507 20364 22573 20365
rect 22507 20300 22508 20364
rect 22572 20300 22573 20364
rect 22507 20299 22573 20300
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 20667 19412 20733 19413
rect 20667 19348 20668 19412
rect 20732 19348 20733 19412
rect 20667 19347 20733 19348
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 16619 15332 16685 15333
rect 16619 15268 16620 15332
rect 16684 15268 16685 15332
rect 16619 15267 16685 15268
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 15331 13836 15397 13837
rect 15331 13772 15332 13836
rect 15396 13772 15397 13836
rect 15331 13771 15397 13772
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 15334 6765 15394 13771
rect 16622 8125 16682 15267
rect 20670 15061 20730 19347
rect 20667 15060 20733 15061
rect 20667 14996 20668 15060
rect 20732 14996 20733 15060
rect 20667 14995 20733 14996
rect 22510 14245 22570 20299
rect 23059 19820 23125 19821
rect 23059 19756 23060 19820
rect 23124 19756 23125 19820
rect 23059 19755 23125 19756
rect 23062 15605 23122 19755
rect 23059 15604 23125 15605
rect 23059 15540 23060 15604
rect 23124 15540 23125 15604
rect 23059 15539 23125 15540
rect 22507 14244 22573 14245
rect 22507 14180 22508 14244
rect 22572 14180 22573 14244
rect 22507 14179 22573 14180
rect 17907 13836 17973 13837
rect 17907 13772 17908 13836
rect 17972 13772 17973 13836
rect 17907 13771 17973 13772
rect 20115 13836 20181 13837
rect 20115 13772 20116 13836
rect 20180 13772 20181 13836
rect 20115 13771 20181 13772
rect 16619 8124 16685 8125
rect 16619 8060 16620 8124
rect 16684 8060 16685 8124
rect 16619 8059 16685 8060
rect 17910 7581 17970 13771
rect 19931 13292 19997 13293
rect 19931 13228 19932 13292
rect 19996 13228 19997 13292
rect 19931 13227 19997 13228
rect 17907 7580 17973 7581
rect 17907 7516 17908 7580
rect 17972 7516 17973 7580
rect 17907 7515 17973 7516
rect 19934 7445 19994 13227
rect 19931 7444 19997 7445
rect 19931 7380 19932 7444
rect 19996 7380 19997 7444
rect 19931 7379 19997 7380
rect 15331 6764 15397 6765
rect 15331 6700 15332 6764
rect 15396 6700 15397 6764
rect 15331 6699 15397 6700
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 20118 4861 20178 13771
rect 20115 4860 20181 4861
rect 20115 4796 20116 4860
rect 20180 4796 20181 4860
rect 20115 4795 20181 4796
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 18001
transform 1 0 20424 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 18001
transform -1 0 24104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 18001
transform 1 0 12696 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 18001
transform 1 0 11960 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 18001
transform 1 0 6808 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 18001
transform 1 0 5336 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 18001
transform 1 0 4324 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 18001
transform 1 0 4416 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 18001
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0630_
timestamp 18001
transform 1 0 3128 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 18001
transform 1 0 10580 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 18001
transform 1 0 10028 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 18001
transform 1 0 10028 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 18001
transform 1 0 14168 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0635_
timestamp 18001
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0636_
timestamp 18001
transform -1 0 12420 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 18001
transform 1 0 15548 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 18001
transform 1 0 16744 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 18001
transform 1 0 19044 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 18001
transform -1 0 20608 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 18001
transform -1 0 22724 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0642_
timestamp 18001
transform -1 0 18952 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 18001
transform -1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0644_
timestamp 18001
transform -1 0 23368 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 18001
transform -1 0 23552 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 18001
transform -1 0 20608 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 18001
transform -1 0 21528 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0648_
timestamp 18001
transform -1 0 21160 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0649_
timestamp 18001
transform -1 0 18952 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 18001
transform 1 0 17388 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0651_
timestamp 18001
transform 1 0 18400 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 18001
transform 1 0 15732 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0653_
timestamp 18001
transform -1 0 13064 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0654_
timestamp 18001
transform 1 0 12512 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 18001
transform -1 0 12696 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 18001
transform -1 0 12052 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 18001
transform 1 0 15824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 18001
transform 1 0 24196 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 18001
transform 1 0 22908 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0660_
timestamp 18001
transform 1 0 22632 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 18001
transform -1 0 22540 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _0662_
timestamp 18001
transform -1 0 26312 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0663_
timestamp 18001
transform -1 0 26404 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0664_
timestamp 18001
transform -1 0 25760 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0665_
timestamp 18001
transform -1 0 25668 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0666_
timestamp 18001
transform -1 0 26496 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0667_
timestamp 18001
transform 1 0 23828 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0668_
timestamp 18001
transform -1 0 25300 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _0669_
timestamp 18001
transform 1 0 25760 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0670_
timestamp 18001
transform -1 0 25116 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0671_
timestamp 18001
transform -1 0 25024 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0672_
timestamp 18001
transform -1 0 20792 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0673_
timestamp 18001
transform 1 0 22908 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _0674_
timestamp 18001
transform 1 0 24472 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0675_
timestamp 18001
transform 1 0 24380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0676_
timestamp 18001
transform -1 0 24196 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0677_
timestamp 18001
transform 1 0 12604 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0678_
timestamp 18001
transform -1 0 5152 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0679_
timestamp 18001
transform 1 0 1656 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0680_
timestamp 18001
transform 1 0 2484 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0681_
timestamp 18001
transform 1 0 1748 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0682_
timestamp 18001
transform -1 0 3588 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0683_
timestamp 18001
transform -1 0 3036 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0684_
timestamp 18001
transform 1 0 4416 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0685_
timestamp 18001
transform 1 0 3036 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _0686_
timestamp 18001
transform -1 0 4784 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0687_
timestamp 18001
transform 1 0 4968 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0688_
timestamp 18001
transform 1 0 2208 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0689_
timestamp 18001
transform -1 0 3956 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0690_
timestamp 18001
transform 1 0 3128 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0691_
timestamp 18001
transform -1 0 4048 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0692_
timestamp 18001
transform 1 0 3956 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0693_
timestamp 18001
transform -1 0 5336 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0694_
timestamp 18001
transform 1 0 4784 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_2  _0695_
timestamp 18001
transform -1 0 6256 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _0696_
timestamp 18001
transform 1 0 3956 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0697_
timestamp 18001
transform -1 0 6716 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0698_
timestamp 18001
transform -1 0 7084 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0699_
timestamp 18001
transform -1 0 6348 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0700_
timestamp 18001
transform -1 0 5428 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0701_
timestamp 18001
transform 1 0 4784 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0702_
timestamp 18001
transform 1 0 5428 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0703_
timestamp 18001
transform -1 0 5612 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _0704_
timestamp 18001
transform 1 0 5704 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0705_
timestamp 18001
transform 1 0 6716 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _0706_
timestamp 18001
transform 1 0 6348 0 1 22848
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0707_
timestamp 18001
transform -1 0 7728 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0708_
timestamp 18001
transform -1 0 6072 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0709_
timestamp 18001
transform 1 0 6440 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0710_
timestamp 18001
transform 1 0 6164 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0711_
timestamp 18001
transform 1 0 7176 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0712_
timestamp 18001
transform 1 0 6532 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0713_
timestamp 18001
transform 1 0 7452 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0714_
timestamp 18001
transform 1 0 7084 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0715_
timestamp 18001
transform -1 0 8188 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 18001
transform 1 0 9568 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0717_
timestamp 18001
transform 1 0 8372 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0718_
timestamp 18001
transform 1 0 8832 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0719_
timestamp 18001
transform 1 0 5060 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0720_
timestamp 18001
transform 1 0 1656 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0721_
timestamp 18001
transform 1 0 2300 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0722_
timestamp 18001
transform -1 0 8096 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0723_
timestamp 18001
transform -1 0 4048 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0724_
timestamp 18001
transform 1 0 1656 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0725_
timestamp 18001
transform 1 0 2300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0726_
timestamp 18001
transform 1 0 1748 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0727_
timestamp 18001
transform -1 0 3128 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0728_
timestamp 18001
transform -1 0 3772 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0729_
timestamp 18001
transform 1 0 2116 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0730_
timestamp 18001
transform -1 0 3772 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0731_
timestamp 18001
transform -1 0 3404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0732_
timestamp 18001
transform -1 0 3864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0733_
timestamp 18001
transform 1 0 1380 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0734_
timestamp 18001
transform 1 0 2300 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0735_
timestamp 18001
transform 1 0 1656 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0736_
timestamp 18001
transform -1 0 2760 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0737_
timestamp 18001
transform 1 0 2024 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0738_
timestamp 18001
transform 1 0 2484 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0739_
timestamp 18001
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0740_
timestamp 18001
transform 1 0 3036 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_2  _0741_
timestamp 18001
transform -1 0 5152 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0742_
timestamp 18001
transform -1 0 3404 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0743_
timestamp 18001
transform 1 0 2852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0744_
timestamp 18001
transform 1 0 4876 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0745_
timestamp 18001
transform -1 0 2852 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0746_
timestamp 18001
transform 1 0 2024 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0747_
timestamp 18001
transform 1 0 1656 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0748_
timestamp 18001
transform 1 0 3220 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0749_
timestamp 18001
transform 1 0 2024 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0750_
timestamp 18001
transform 1 0 2392 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0751_
timestamp 18001
transform 1 0 4140 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0752_
timestamp 18001
transform 1 0 2944 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0753_
timestamp 18001
transform 1 0 4048 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0754_
timestamp 18001
transform -1 0 5704 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0755_
timestamp 18001
transform 1 0 5060 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0756_
timestamp 18001
transform 1 0 6440 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0757_
timestamp 18001
transform -1 0 4416 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0758_
timestamp 18001
transform 1 0 2760 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0759_
timestamp 18001
transform 1 0 4968 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _0760_
timestamp 18001
transform -1 0 2852 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0761_
timestamp 18001
transform 1 0 2760 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0762_
timestamp 18001
transform 1 0 1380 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0763_
timestamp 18001
transform 1 0 3496 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0764_
timestamp 18001
transform 1 0 2300 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0765_
timestamp 18001
transform 1 0 3036 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _0766_
timestamp 18001
transform -1 0 3496 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0767_
timestamp 18001
transform 1 0 4600 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0768_
timestamp 18001
transform 1 0 3404 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0769_
timestamp 18001
transform 1 0 4140 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0770_
timestamp 18001
transform 1 0 5244 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0771_
timestamp 18001
transform 1 0 4968 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0772_
timestamp 18001
transform 1 0 6348 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0773_
timestamp 18001
transform -1 0 7912 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0774_
timestamp 18001
transform 1 0 5336 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0775_
timestamp 18001
transform 1 0 3036 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0776_
timestamp 18001
transform -1 0 4048 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0777_
timestamp 18001
transform 1 0 2024 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0778_
timestamp 18001
transform 1 0 3496 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0779_
timestamp 18001
transform 1 0 4140 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0780_
timestamp 18001
transform 1 0 2852 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0781_
timestamp 18001
transform -1 0 4508 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0782_
timestamp 18001
transform 1 0 2852 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0783_
timestamp 18001
transform 1 0 4508 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0784_
timestamp 18001
transform 1 0 3864 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0785_
timestamp 18001
transform -1 0 5612 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0786_
timestamp 18001
transform 1 0 4416 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0787_
timestamp 18001
transform 1 0 6348 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0788_
timestamp 18001
transform 1 0 5428 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_2  _0789_
timestamp 18001
transform 1 0 6532 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _0790_
timestamp 18001
transform 1 0 6072 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0791_
timestamp 18001
transform -1 0 7820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0792_
timestamp 18001
transform 1 0 7268 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0793_
timestamp 18001
transform 1 0 6808 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0794_
timestamp 18001
transform 1 0 4416 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0795_
timestamp 18001
transform 1 0 3772 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0796_
timestamp 18001
transform 1 0 7360 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0797_
timestamp 18001
transform 1 0 6348 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0798_
timestamp 18001
transform -1 0 7176 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0799_
timestamp 18001
transform -1 0 6992 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0800_
timestamp 18001
transform -1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0801_
timestamp 18001
transform 1 0 5704 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0802_
timestamp 18001
transform -1 0 6716 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0803_
timestamp 18001
transform 1 0 5152 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0804_
timestamp 18001
transform 1 0 5612 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0805_
timestamp 18001
transform -1 0 6992 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0806_
timestamp 18001
transform 1 0 5060 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0807_
timestamp 18001
transform 1 0 7820 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0808_
timestamp 18001
transform 1 0 6808 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0809_
timestamp 18001
transform 1 0 6808 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0810_
timestamp 18001
transform 1 0 7084 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0811_
timestamp 18001
transform -1 0 7544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0812_
timestamp 18001
transform 1 0 7544 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0813_
timestamp 18001
transform 1 0 7544 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0814_
timestamp 18001
transform -1 0 8188 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0815_
timestamp 18001
transform 1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0816_
timestamp 18001
transform -1 0 8740 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0817_
timestamp 18001
transform -1 0 8648 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0818_
timestamp 18001
transform -1 0 8648 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0819_
timestamp 18001
transform -1 0 8556 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _0820_
timestamp 18001
transform -1 0 7544 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _0821_
timestamp 18001
transform -1 0 8832 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _0822_
timestamp 18001
transform 1 0 8648 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _0823_
timestamp 18001
transform 1 0 6072 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__o31ai_4  _0824_
timestamp 18001
transform 1 0 3864 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__a31o_1  _0825_
timestamp 18001
transform -1 0 3680 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 18001
transform -1 0 4232 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0827_
timestamp 18001
transform 1 0 1932 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0828_
timestamp 18001
transform -1 0 3312 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0829_
timestamp 18001
transform 1 0 2576 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0830_
timestamp 18001
transform 1 0 3496 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0831_
timestamp 18001
transform 1 0 5336 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0832_
timestamp 18001
transform 1 0 4140 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0833_
timestamp 18001
transform 1 0 4600 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0834_
timestamp 18001
transform 1 0 5612 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _0835_
timestamp 18001
transform 1 0 4416 0 1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _0836_
timestamp 18001
transform 1 0 6440 0 1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_1  _0837_
timestamp 18001
transform 1 0 8188 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _0838_
timestamp 18001
transform 1 0 6808 0 1 15232
box -38 -48 2062 592
use sky130_fd_sc_hd__o31ai_4  _0839_
timestamp 18001
transform 1 0 4692 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__a31o_2  _0840_
timestamp 18001
transform -1 0 4416 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0841_
timestamp 18001
transform 1 0 4048 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0842_
timestamp 18001
transform -1 0 5152 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _0843_
timestamp 18001
transform 1 0 4600 0 1 21760
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_4  _0844_
timestamp 18001
transform 1 0 5428 0 1 20672
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0845_
timestamp 18001
transform -1 0 6624 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _0846_
timestamp 18001
transform 1 0 5796 0 1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _0847_
timestamp 18001
transform 1 0 6532 0 1 17408
box -38 -48 2062 592
use sky130_fd_sc_hd__a21boi_4  _0848_
timestamp 18001
transform 1 0 6348 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__xnor2_4  _0849_
timestamp 18001
transform 1 0 7544 0 -1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _0850_
timestamp 18001
transform 1 0 10212 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0851_
timestamp 18001
transform 1 0 5336 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _0852_
timestamp 18001
transform 1 0 5152 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0853_
timestamp 18001
transform 1 0 6716 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0854_
timestamp 18001
transform 1 0 7452 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0855_
timestamp 18001
transform 1 0 7452 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_2  _0856_
timestamp 18001
transform 1 0 6716 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0857_
timestamp 18001
transform -1 0 9844 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0858_
timestamp 18001
transform 1 0 8924 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 18001
transform 1 0 10120 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_4  _0860_
timestamp 18001
transform 1 0 7176 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__xnor2_4  _0861_
timestamp 18001
transform 1 0 7268 0 -1 21760
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _0862_
timestamp 18001
transform 1 0 8280 0 -1 19584
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _0863_
timestamp 18001
transform -1 0 9476 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0864_
timestamp 18001
transform -1 0 7544 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0865_
timestamp 18001
transform 1 0 7544 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0866_
timestamp 18001
transform 1 0 9200 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0867_
timestamp 18001
transform 1 0 8188 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0868_
timestamp 18001
transform -1 0 8280 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a41oi_4  _0869_
timestamp 18001
transform 1 0 8924 0 1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0870_
timestamp 18001
transform 1 0 9384 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0871_
timestamp 18001
transform -1 0 10120 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0872_
timestamp 18001
transform 1 0 7360 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0873_
timestamp 18001
transform 1 0 6716 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0874_
timestamp 18001
transform 1 0 7452 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _0875_
timestamp 18001
transform 1 0 6900 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0876_
timestamp 18001
transform 1 0 8004 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0877_
timestamp 18001
transform 1 0 8188 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0878_
timestamp 18001
transform -1 0 8188 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0879_
timestamp 18001
transform 1 0 8648 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0880_
timestamp 18001
transform -1 0 8924 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _0881_
timestamp 18001
transform -1 0 9476 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0882_
timestamp 18001
transform 1 0 9384 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0883_
timestamp 18001
transform -1 0 11960 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0884_
timestamp 18001
transform -1 0 12972 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0885_
timestamp 18001
transform -1 0 12512 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_2  _0886_
timestamp 18001
transform -1 0 12052 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0887_
timestamp 18001
transform -1 0 11132 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0888_
timestamp 18001
transform -1 0 12144 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0889_
timestamp 18001
transform -1 0 12604 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0890_
timestamp 18001
transform 1 0 9936 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0891_
timestamp 18001
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0892_
timestamp 18001
transform -1 0 10764 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _0893_
timestamp 18001
transform 1 0 10580 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0894_
timestamp 18001
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0895_
timestamp 18001
transform 1 0 10672 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0896_
timestamp 18001
transform -1 0 9844 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0897_
timestamp 18001
transform -1 0 9568 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0898_
timestamp 18001
transform -1 0 9936 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0899_
timestamp 18001
transform 1 0 9660 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0900_
timestamp 18001
transform 1 0 10120 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0901_
timestamp 18001
transform 1 0 10028 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0902_
timestamp 18001
transform 1 0 9936 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0903_
timestamp 18001
transform -1 0 9384 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0904_
timestamp 18001
transform 1 0 9200 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0905_
timestamp 18001
transform 1 0 10212 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0906_
timestamp 18001
transform -1 0 11316 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0907_
timestamp 18001
transform -1 0 12788 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0908_
timestamp 18001
transform -1 0 13432 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0909_
timestamp 18001
transform 1 0 12604 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0910_
timestamp 18001
transform 1 0 12788 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0911_
timestamp 18001
transform 1 0 12052 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _0912_
timestamp 18001
transform -1 0 12788 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_1  _0913_
timestamp 18001
transform -1 0 12696 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0914_
timestamp 18001
transform 1 0 12696 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_4  _0915_
timestamp 18001
transform 1 0 11684 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__o21a_1  _0916_
timestamp 18001
transform -1 0 13064 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0917_
timestamp 18001
transform 1 0 13984 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0918_
timestamp 18001
transform -1 0 13892 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0919_
timestamp 18001
transform 1 0 13432 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0920_
timestamp 18001
transform -1 0 13524 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0921_
timestamp 18001
transform -1 0 14720 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0922_
timestamp 18001
transform 1 0 12144 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0923_
timestamp 18001
transform -1 0 11868 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0924_
timestamp 18001
transform 1 0 12420 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0925_
timestamp 18001
transform -1 0 12420 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0926_
timestamp 18001
transform 1 0 11776 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0927_
timestamp 18001
transform -1 0 13064 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0928_
timestamp 18001
transform 1 0 14076 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0929_
timestamp 18001
transform 1 0 14444 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor3b_1  _0930_
timestamp 18001
transform -1 0 17204 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0931_
timestamp 18001
transform 1 0 16652 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0932_
timestamp 18001
transform -1 0 10304 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0933_
timestamp 18001
transform -1 0 16468 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0934_
timestamp 18001
transform -1 0 15364 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _0935_
timestamp 18001
transform 1 0 15456 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0936_
timestamp 18001
transform 1 0 15364 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0937_
timestamp 18001
transform 1 0 15916 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0938_
timestamp 18001
transform -1 0 17848 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0939_
timestamp 18001
transform 1 0 16744 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0940_
timestamp 18001
transform 1 0 16836 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0941_
timestamp 18001
transform 1 0 10304 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0942_
timestamp 18001
transform 1 0 15088 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0943_
timestamp 18001
transform -1 0 18216 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0944_
timestamp 18001
transform -1 0 18768 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0945_
timestamp 18001
transform -1 0 11132 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0946_
timestamp 18001
transform 1 0 11132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0947_
timestamp 18001
transform -1 0 18400 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0948_
timestamp 18001
transform -1 0 19136 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _0949_
timestamp 18001
transform 1 0 18400 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _0950_
timestamp 18001
transform 1 0 9660 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0951_
timestamp 18001
transform 1 0 21160 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0952_
timestamp 18001
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a311oi_1  _0953_
timestamp 18001
transform 1 0 16652 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _0954_
timestamp 18001
transform -1 0 17848 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0955_
timestamp 18001
transform 1 0 16376 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_1  _0956_
timestamp 18001
transform -1 0 15088 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _0957_
timestamp 18001
transform -1 0 14444 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0958_
timestamp 18001
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _0959_
timestamp 18001
transform 1 0 13984 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0960_
timestamp 18001
transform -1 0 13984 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0961_
timestamp 18001
transform -1 0 21160 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0962_
timestamp 18001
transform -1 0 20424 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0963_
timestamp 18001
transform -1 0 19780 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0964_
timestamp 18001
transform -1 0 18308 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0965_
timestamp 18001
transform -1 0 9384 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _0966_
timestamp 18001
transform -1 0 10120 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _0967_
timestamp 18001
transform 1 0 9384 0 -1 17408
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 18001
transform -1 0 17480 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0969_
timestamp 18001
transform 1 0 9476 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0970_
timestamp 18001
transform 1 0 19872 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0971_
timestamp 18001
transform -1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0972_
timestamp 18001
transform -1 0 20056 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _0973_
timestamp 18001
transform -1 0 10212 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _0974_
timestamp 18001
transform 1 0 9108 0 1 15232
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0975_
timestamp 18001
transform -1 0 16192 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0976_
timestamp 18001
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0977_
timestamp 18001
transform 1 0 20884 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _0978_
timestamp 18001
transform 1 0 9108 0 -1 15232
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_1  _0979_
timestamp 18001
transform -1 0 21252 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0980_
timestamp 18001
transform -1 0 20792 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0981_
timestamp 18001
transform 1 0 8464 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0982_
timestamp 18001
transform 1 0 8924 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 18001
transform -1 0 18492 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0984_
timestamp 18001
transform -1 0 19136 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0985_
timestamp 18001
transform 1 0 18584 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0986_
timestamp 18001
transform 1 0 8556 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 18001
transform 1 0 18124 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0988_
timestamp 18001
transform -1 0 20700 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0989_
timestamp 18001
transform -1 0 20056 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0990_
timestamp 18001
transform 1 0 8924 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0991_
timestamp 18001
transform 1 0 9384 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0992_
timestamp 18001
transform 1 0 16100 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0993_
timestamp 18001
transform 1 0 8464 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0994_
timestamp 18001
transform 1 0 8924 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 18001
transform -1 0 16100 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0996_
timestamp 18001
transform 1 0 7912 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0997_
timestamp 18001
transform 1 0 8372 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 18001
transform 1 0 14168 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0999_
timestamp 18001
transform 1 0 14444 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1000_
timestamp 18001
transform 1 0 7544 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1001_
timestamp 18001
transform 1 0 8648 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1002_
timestamp 18001
transform 1 0 14076 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1003_
timestamp 18001
transform -1 0 12052 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1004_
timestamp 18001
transform -1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1005_
timestamp 18001
transform 1 0 11776 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1006_
timestamp 18001
transform -1 0 13156 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1007_
timestamp 18001
transform -1 0 12328 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1008_
timestamp 18001
transform -1 0 11408 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1009_
timestamp 18001
transform 1 0 10304 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1010_
timestamp 18001
transform 1 0 12328 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1011_
timestamp 18001
transform 1 0 11684 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _1012_
timestamp 18001
transform -1 0 13984 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1013_
timestamp 18001
transform 1 0 15732 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1014_
timestamp 18001
transform 1 0 8924 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1015_
timestamp 18001
transform -1 0 9384 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 18001
transform 1 0 19688 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1017_
timestamp 18001
transform 1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1018_
timestamp 18001
transform -1 0 19688 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1019_
timestamp 18001
transform 1 0 8924 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1020_
timestamp 18001
transform -1 0 9384 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1021_
timestamp 18001
transform 1 0 17664 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_1  _1022_
timestamp 18001
transform -1 0 18492 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1023_
timestamp 18001
transform 1 0 17940 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _1024_
timestamp 18001
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1025_
timestamp 18001
transform 1 0 18492 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1026_
timestamp 18001
transform -1 0 19412 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1027_
timestamp 18001
transform 1 0 19872 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1028_
timestamp 18001
transform -1 0 20884 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1029_
timestamp 18001
transform 1 0 20792 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1030_
timestamp 18001
transform 1 0 19780 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1031_
timestamp 18001
transform 1 0 19228 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a41oi_4  _1032_
timestamp 18001
transform 1 0 17296 0 -1 21760
box -38 -48 2062 592
use sky130_fd_sc_hd__a41o_1  _1033_
timestamp 18001
transform 1 0 17296 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1034_
timestamp 18001
transform 1 0 17756 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1035_
timestamp 18001
transform 1 0 23276 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1036_
timestamp 18001
transform -1 0 24288 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1037_
timestamp 18001
transform 1 0 12696 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1038_
timestamp 18001
transform 1 0 12328 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1039_
timestamp 18001
transform 1 0 15364 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1040_
timestamp 18001
transform 1 0 16468 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1041_
timestamp 18001
transform 1 0 18124 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1042_
timestamp 18001
transform -1 0 18124 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _1043_
timestamp 18001
transform -1 0 22448 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1044_
timestamp 18001
transform 1 0 8188 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1045_
timestamp 18001
transform 1 0 9384 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1046_
timestamp 18001
transform 1 0 9844 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1047_
timestamp 18001
transform 1 0 18860 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1048_
timestamp 18001
transform 1 0 21896 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _1049_
timestamp 18001
transform 1 0 23184 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1050_
timestamp 18001
transform -1 0 22448 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1051_
timestamp 18001
transform -1 0 22908 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _1052_
timestamp 18001
transform -1 0 23644 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1053_
timestamp 18001
transform -1 0 24104 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1054_
timestamp 18001
transform -1 0 25392 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1055_
timestamp 18001
transform 1 0 22816 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _1056_
timestamp 18001
transform -1 0 24012 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1057_
timestamp 18001
transform -1 0 25208 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1058_
timestamp 18001
transform 1 0 22724 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1059_
timestamp 18001
transform -1 0 24196 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1060_
timestamp 18001
transform 1 0 24288 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1061_
timestamp 18001
transform -1 0 24012 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1062_
timestamp 18001
transform -1 0 24472 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1063_
timestamp 18001
transform -1 0 23920 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1064_
timestamp 18001
transform 1 0 22816 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1065_
timestamp 18001
transform 1 0 21988 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1066_
timestamp 18001
transform -1 0 22816 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1067_
timestamp 18001
transform -1 0 23920 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1068_
timestamp 18001
transform -1 0 21528 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1069_
timestamp 18001
transform 1 0 21804 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1070_
timestamp 18001
transform 1 0 22908 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1071_
timestamp 18001
transform 1 0 22356 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1072_
timestamp 18001
transform 1 0 25300 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1073_
timestamp 18001
transform 1 0 15180 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1074_
timestamp 18001
transform 1 0 13616 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1075_
timestamp 18001
transform 1 0 14444 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1076_
timestamp 18001
transform 1 0 14904 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1077_
timestamp 18001
transform -1 0 14904 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1078_
timestamp 18001
transform 1 0 11316 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1079_
timestamp 18001
transform 1 0 12144 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1080_
timestamp 18001
transform 1 0 12604 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _1081_
timestamp 18001
transform 1 0 11776 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1082_
timestamp 18001
transform 1 0 10764 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1083_
timestamp 18001
transform 1 0 10396 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1084_
timestamp 18001
transform 1 0 11500 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1085_
timestamp 18001
transform 1 0 12696 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1086_
timestamp 18001
transform 1 0 12144 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _1087_
timestamp 18001
transform 1 0 11868 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1088_
timestamp 18001
transform -1 0 11408 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1089_
timestamp 18001
transform 1 0 11132 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 18001
transform -1 0 11224 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1091_
timestamp 18001
transform 1 0 12420 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1092_
timestamp 18001
transform 1 0 11868 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1093_
timestamp 18001
transform -1 0 12604 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1094_
timestamp 18001
transform -1 0 12696 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1095_
timestamp 18001
transform 1 0 12972 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1096_
timestamp 18001
transform 1 0 11868 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1097_
timestamp 18001
transform -1 0 11776 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1098_
timestamp 18001
transform -1 0 13708 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1099_
timestamp 18001
transform 1 0 12696 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1100_
timestamp 18001
transform -1 0 12788 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _1101_
timestamp 18001
transform 1 0 12512 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a221oi_2  _1102_
timestamp 18001
transform 1 0 11960 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _1103_
timestamp 18001
transform -1 0 15364 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1104_
timestamp 18001
transform -1 0 14720 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1105_
timestamp 18001
transform 1 0 14720 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1106_
timestamp 18001
transform -1 0 15732 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1107_
timestamp 18001
transform 1 0 15916 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1108_
timestamp 18001
transform 1 0 14352 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1109_
timestamp 18001
transform -1 0 16100 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1110_
timestamp 18001
transform 1 0 15088 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1111_
timestamp 18001
transform 1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1112_
timestamp 18001
transform 1 0 15180 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1113_
timestamp 18001
transform 1 0 16744 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1114_
timestamp 18001
transform 1 0 16100 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1115_
timestamp 18001
transform 1 0 17480 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1116_
timestamp 18001
transform 1 0 16652 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1117_
timestamp 18001
transform -1 0 17480 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1118_
timestamp 18001
transform -1 0 17296 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1119_
timestamp 18001
transform 1 0 18124 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_2  _1120_
timestamp 18001
transform -1 0 17480 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _1121_
timestamp 18001
transform -1 0 18676 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1122_
timestamp 18001
transform 1 0 19228 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1123_
timestamp 18001
transform -1 0 18952 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _1124_
timestamp 18001
transform 1 0 19596 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a221oi_4  _1125_
timestamp 18001
transform 1 0 17664 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__a211o_1  _1126_
timestamp 18001
transform 1 0 20332 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1127_
timestamp 18001
transform 1 0 21068 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1128_
timestamp 18001
transform 1 0 20976 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1129_
timestamp 18001
transform 1 0 21804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1130_
timestamp 18001
transform 1 0 19412 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1131_
timestamp 18001
transform 1 0 20608 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1132_
timestamp 18001
transform 1 0 20332 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1133_
timestamp 18001
transform -1 0 21068 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _1134_
timestamp 18001
transform 1 0 20792 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1135_
timestamp 18001
transform 1 0 20700 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1136_
timestamp 18001
transform 1 0 20056 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1137_
timestamp 18001
transform 1 0 19780 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1138_
timestamp 18001
transform 1 0 21252 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1139_
timestamp 18001
transform -1 0 21252 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1140_
timestamp 18001
transform 1 0 21804 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1141_
timestamp 18001
transform -1 0 20884 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1142_
timestamp 18001
transform 1 0 19504 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1143_
timestamp 18001
transform -1 0 19504 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1144_
timestamp 18001
transform -1 0 23092 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1145_
timestamp 18001
transform -1 0 25024 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1146_
timestamp 18001
transform 1 0 23552 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_2  _1147_
timestamp 18001
transform 1 0 22448 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_1  _1148_
timestamp 18001
transform -1 0 23092 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1149_
timestamp 18001
transform -1 0 24840 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1150_
timestamp 18001
transform 1 0 23736 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _1151_
timestamp 18001
transform -1 0 24012 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1152_
timestamp 18001
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1153_
timestamp 18001
transform 1 0 23092 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1154_
timestamp 18001
transform -1 0 22448 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1155_
timestamp 18001
transform -1 0 23460 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1156_
timestamp 18001
transform 1 0 23460 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1157_
timestamp 18001
transform -1 0 22816 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1158_
timestamp 18001
transform 1 0 20700 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_2  _1159_
timestamp 18001
transform 1 0 21528 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _1160_
timestamp 18001
transform -1 0 21896 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1161_
timestamp 18001
transform -1 0 18216 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1162_
timestamp 18001
transform 1 0 17664 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1163_
timestamp 18001
transform -1 0 17020 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1164_
timestamp 18001
transform 1 0 21528 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1165_
timestamp 18001
transform -1 0 22264 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1166_
timestamp 18001
transform 1 0 22264 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1167_
timestamp 18001
transform -1 0 22724 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1168_
timestamp 18001
transform 1 0 20516 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1169_
timestamp 18001
transform -1 0 22172 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1170_
timestamp 18001
transform 1 0 22172 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1171_
timestamp 18001
transform -1 0 19964 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1172_
timestamp 18001
transform -1 0 20884 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1173_
timestamp 18001
transform -1 0 19228 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o221ai_2  _1174_
timestamp 18001
transform -1 0 20332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _1175_
timestamp 18001
transform 1 0 18400 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1176_
timestamp 18001
transform 1 0 18492 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1177_
timestamp 18001
transform 1 0 18768 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1178_
timestamp 18001
transform 1 0 19320 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1179_
timestamp 18001
transform 1 0 19596 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1180_
timestamp 18001
transform 1 0 18584 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1181_
timestamp 18001
transform 1 0 18032 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1182_
timestamp 18001
transform 1 0 18768 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1183_
timestamp 18001
transform -1 0 17388 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1184_
timestamp 18001
transform -1 0 16560 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1185_
timestamp 18001
transform 1 0 17296 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o221ai_2  _1186_
timestamp 18001
transform -1 0 17756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _1187_
timestamp 18001
transform 1 0 16284 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1188_
timestamp 18001
transform -1 0 16376 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1189_
timestamp 18001
transform 1 0 14812 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1190_
timestamp 18001
transform -1 0 15548 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1191_
timestamp 18001
transform -1 0 15180 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1192_
timestamp 18001
transform -1 0 14628 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1193_
timestamp 18001
transform 1 0 15824 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1194_
timestamp 18001
transform 1 0 14628 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1195_
timestamp 18001
transform -1 0 14352 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1196_
timestamp 18001
transform 1 0 10764 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1197_
timestamp 18001
transform -1 0 12880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1198_
timestamp 18001
transform -1 0 12604 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a41oi_2  _1199_
timestamp 18001
transform 1 0 11500 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__a221oi_2  _1200_
timestamp 18001
transform -1 0 12144 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_1  _1201_
timestamp 18001
transform 1 0 12144 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1202_
timestamp 18001
transform -1 0 15272 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1203_
timestamp 18001
transform 1 0 15088 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1204_
timestamp 18001
transform -1 0 14628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _1205_
timestamp 18001
transform 1 0 11868 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1206_
timestamp 18001
transform 1 0 12512 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1207_
timestamp 18001
transform 1 0 12788 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _1208_
timestamp 18001
transform 1 0 11960 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1209_
timestamp 18001
transform 1 0 12052 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1210_
timestamp 18001
transform -1 0 23644 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1211_
timestamp 18001
transform -1 0 18676 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1212_
timestamp 18001
transform -1 0 23828 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1213_
timestamp 18001
transform 1 0 23000 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1214_
timestamp 18001
transform 1 0 22448 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1215_
timestamp 18001
transform 1 0 15272 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_1  _1216_
timestamp 18001
transform -1 0 15364 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1217_
timestamp 18001
transform 1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1218_
timestamp 18001
transform -1 0 11040 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1219_
timestamp 18001
transform 1 0 15364 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1220_
timestamp 18001
transform -1 0 21344 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1221_
timestamp 18001
transform -1 0 22172 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1222_
timestamp 18001
transform -1 0 19136 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o2111ai_1  _1223_
timestamp 18001
transform 1 0 19228 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1224_
timestamp 18001
transform -1 0 15088 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1225_
timestamp 18001
transform 1 0 13616 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1226_
timestamp 18001
transform -1 0 15180 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1227_
timestamp 18001
transform -1 0 15456 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1228_
timestamp 18001
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1229_
timestamp 18001
transform -1 0 18124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1230_
timestamp 18001
transform 1 0 12880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1231_
timestamp 18001
transform 1 0 16836 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o2111ai_1  _1232_
timestamp 18001
transform -1 0 16744 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1233_
timestamp 18001
transform 1 0 15088 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _1234_
timestamp 18001
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1235_
timestamp 18001
transform -1 0 11316 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_1  _1236_
timestamp 18001
transform 1 0 14076 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1237_
timestamp 18001
transform 1 0 15732 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1238_
timestamp 18001
transform -1 0 11684 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1239_
timestamp 18001
transform 1 0 13800 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _1240_
timestamp 18001
transform 1 0 11960 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1241_
timestamp 18001
transform 1 0 11776 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1242_
timestamp 18001
transform 1 0 15456 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1243_
timestamp 18001
transform 1 0 11592 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1244_
timestamp 18001
transform 1 0 12880 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1245_
timestamp 18001
transform -1 0 21068 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _1246_
timestamp 18001
transform 1 0 17204 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1247_
timestamp 18001
transform 1 0 17756 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o32ai_1  _1248_
timestamp 18001
transform 1 0 17296 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1249_
timestamp 18001
transform -1 0 15180 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _1250_
timestamp 18001
transform 1 0 14720 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1251_
timestamp 18001
transform -1 0 17388 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1252_
timestamp 18001
transform 1 0 16100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1253_
timestamp 18001
transform 1 0 16836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1254_
timestamp 18001
transform -1 0 25944 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1255_
timestamp 18001
transform -1 0 26864 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1256_
timestamp 18001
transform 1 0 26956 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1257_
timestamp 18001
transform -1 0 26128 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1258_
timestamp 18001
transform 1 0 26128 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1259_
timestamp 18001
transform 1 0 25944 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1260_
timestamp 18001
transform 1 0 26864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1261_
timestamp 18001
transform -1 0 19136 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1262_
timestamp 18001
transform 1 0 25576 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1263_
timestamp 18001
transform 1 0 26404 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1264_
timestamp 18001
transform 1 0 26496 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1265_
timestamp 18001
transform -1 0 20424 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1266_
timestamp 18001
transform -1 0 18492 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1267_
timestamp 18001
transform 1 0 24656 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1268_
timestamp 18001
transform 1 0 25668 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1269_
timestamp 18001
transform 1 0 19504 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _1270_
timestamp 18001
transform -1 0 19320 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1271_
timestamp 18001
transform 1 0 17756 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1272_
timestamp 18001
transform -1 0 21712 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1273_
timestamp 18001
transform -1 0 20332 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1274_
timestamp 18001
transform 1 0 17756 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1275_
timestamp 18001
transform 1 0 20884 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1276_
timestamp 18001
transform -1 0 22908 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1277_
timestamp 18001
transform 1 0 24196 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1278_
timestamp 18001
transform -1 0 24288 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1279_
timestamp 18001
transform -1 0 19964 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1280_
timestamp 18001
transform -1 0 18308 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _1281_
timestamp 18001
transform 1 0 24380 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1282_
timestamp 18001
transform -1 0 26128 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _1283_
timestamp 18001
transform -1 0 21252 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _1284_
timestamp 18001
transform 1 0 22356 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1285_
timestamp 18001
transform 1 0 25208 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1286_
timestamp 18001
transform 1 0 26220 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1287_
timestamp 18001
transform -1 0 19504 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1288_
timestamp 18001
transform -1 0 20608 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1289_
timestamp 18001
transform 1 0 23092 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _1290_
timestamp 18001
transform -1 0 22908 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _1291_
timestamp 18001
transform 1 0 22908 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1292_
timestamp 18001
transform 1 0 25668 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1293_
timestamp 18001
transform -1 0 21252 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1294_
timestamp 18001
transform 1 0 21804 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1295_
timestamp 18001
transform 1 0 17204 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1296_
timestamp 18001
transform 1 0 24932 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1297_
timestamp 18001
transform -1 0 20884 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1298_
timestamp 18001
transform -1 0 18216 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1299_
timestamp 18001
transform 1 0 21528 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1300_
timestamp 18001
transform -1 0 26312 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1301_
timestamp 18001
transform 1 0 17480 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1302_
timestamp 18001
transform 1 0 26312 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1303_
timestamp 18001
transform 1 0 24748 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1304_
timestamp 18001
transform 1 0 25944 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1305_
timestamp 18001
transform -1 0 26220 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1306_
timestamp 18001
transform -1 0 20608 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1307_
timestamp 18001
transform 1 0 19504 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1308_
timestamp 18001
transform 1 0 25208 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1309_
timestamp 18001
transform 1 0 26956 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1310_
timestamp 18001
transform -1 0 27416 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1311_
timestamp 18001
transform 1 0 26588 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  _1312_
timestamp 18001
transform 1 0 23276 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1313_
timestamp 18001
transform 1 0 24380 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1314_
timestamp 18001
transform 1 0 24380 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1315_
timestamp 18001
transform 1 0 22448 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1316_
timestamp 18001
transform 1 0 14076 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1317_
timestamp 18001
transform 1 0 10212 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1318_
timestamp 18001
transform 1 0 10212 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1319_
timestamp 18001
transform 1 0 11040 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1320_
timestamp 18001
transform 1 0 11500 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1321_
timestamp 18001
transform 1 0 14076 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1322_
timestamp 18001
transform 1 0 16100 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1323_
timestamp 18001
transform 1 0 16192 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1324_
timestamp 18001
transform 1 0 17388 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1325_
timestamp 18001
transform 1 0 19780 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1326_
timestamp 18001
transform 1 0 20148 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1327_
timestamp 18001
transform 1 0 19504 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1328_
timestamp 18001
transform 1 0 23552 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1329_
timestamp 18001
transform 1 0 23368 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1330_
timestamp 18001
transform 1 0 22448 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1331_
timestamp 18001
transform 1 0 17020 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1332_
timestamp 18001
transform 1 0 21804 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1333_
timestamp 18001
transform 1 0 18952 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1334_
timestamp 18001
transform -1 0 21160 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1335_
timestamp 18001
transform 1 0 15640 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1336_
timestamp 18001
transform 1 0 13248 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1337_
timestamp 18001
transform 1 0 10304 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1338_
timestamp 18001
transform 1 0 14076 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1339_
timestamp 18001
transform 1 0 11684 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1340_
timestamp 18001
transform 1 0 22448 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1341_
timestamp 18001
transform 1 0 25024 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1342_
timestamp 18001
transform 1 0 24656 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1343_
timestamp 18001
transform -1 0 23644 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1344_
timestamp 18001
transform -1 0 21712 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1345_
timestamp 18001
transform 1 0 21528 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1346_
timestamp 18001
transform 1 0 23736 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1347_
timestamp 18001
transform 1 0 26036 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 18001
transform -1 0 20056 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 18001
transform -1 0 18492 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 18001
transform 1 0 19780 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 18001
transform 1 0 17112 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 18001
transform 1 0 20056 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkload0
timestamp 18001
transform 1 0 16652 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_2  clkload1
timestamp 18001
transform -1 0 19780 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  clkload2
timestamp 18001
transform 1 0 16744 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout53
timestamp 18001
transform 1 0 22540 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout54
timestamp 18001
transform -1 0 19596 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout55
timestamp 18001
transform 1 0 18032 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout56
timestamp 18001
transform 1 0 20240 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout57
timestamp 18001
transform 1 0 19412 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout58
timestamp 18001
transform -1 0 16284 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout59
timestamp 18001
transform -1 0 13064 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout60
timestamp 18001
transform 1 0 15456 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout61
timestamp 18001
transform -1 0 15824 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout62
timestamp 18001
transform -1 0 17756 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout63
timestamp 18001
transform -1 0 20332 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout64
timestamp 18001
transform 1 0 21896 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout65
timestamp 18001
transform 1 0 23000 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout66
timestamp 18001
transform 1 0 21896 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout67
timestamp 18001
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout68
timestamp 18001
transform -1 0 22540 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout69
timestamp 18001
transform -1 0 21988 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout70
timestamp 18001
transform -1 0 23736 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout71
timestamp 18001
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout72
timestamp 18001
transform -1 0 25852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout73
timestamp 18001
transform -1 0 27324 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout74
timestamp 18001
transform -1 0 27692 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  fanout75
timestamp 18001
transform 1 0 21620 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout76
timestamp 18001
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout77
timestamp 18001
transform -1 0 22080 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout78
timestamp 18001
transform 1 0 7452 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout79
timestamp 18001
transform -1 0 3496 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout80
timestamp 18001
transform -1 0 3680 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout81
timestamp 18001
transform 1 0 12788 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout82
timestamp 18001
transform -1 0 2760 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout83
timestamp 18001
transform -1 0 25024 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout84
timestamp 18001
transform 1 0 25208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout85
timestamp 18001
transform 1 0 24564 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout86
timestamp 18001
transform -1 0 25300 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout87
timestamp 18001
transform -1 0 2484 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout88
timestamp 18001
transform -1 0 23460 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout89
timestamp 18001
transform 1 0 22540 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout90
timestamp 18001
transform 1 0 25392 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout91
timestamp 18001
transform -1 0 22724 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636986456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636986456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 18001
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636986456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_41
timestamp 18001
transform 1 0 4876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_49
timestamp 18001
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 18001
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636986456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_69
timestamp 18001
transform 1 0 7452 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_77
timestamp 18001
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1636986456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1636986456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 18001
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1636986456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1636986456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 18001
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1636986456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1636986456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 18001
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1636986456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1636986456
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 18001
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1636986456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1636986456
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 18001
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1636986456
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1636986456
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 18001
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1636986456
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1636986456
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 18001
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_281
timestamp 18001
transform 1 0 26956 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_289
timestamp 18001
transform 1 0 27692 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636986456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636986456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636986456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1636986456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 18001
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 18001
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1636986456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1636986456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1636986456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1636986456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 18001
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 18001
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1636986456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1636986456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1636986456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1636986456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 18001
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 18001
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1636986456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1636986456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1636986456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1636986456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 18001
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 18001
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1636986456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1636986456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1636986456
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1636986456
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 18001
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 18001
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_281
timestamp 18001
transform 1 0 26956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_289
timestamp 18001
transform 1 0 27692 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636986456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636986456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 18001
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1636986456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1636986456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1636986456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1636986456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 18001
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 18001
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1636986456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1636986456
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1636986456
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1636986456
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 18001
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 18001
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1636986456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1636986456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1636986456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1636986456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 18001
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 18001
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1636986456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1636986456
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1636986456
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1636986456
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 18001
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 18001
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1636986456
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1636986456
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1636986456
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_289
timestamp 18001
transform 1 0 27692 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636986456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636986456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1636986456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1636986456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 18001
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 18001
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1636986456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1636986456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1636986456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1636986456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 18001
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 18001
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1636986456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1636986456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1636986456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1636986456
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 18001
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 18001
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1636986456
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1636986456
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1636986456
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1636986456
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 18001
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 18001
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1636986456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1636986456
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1636986456
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1636986456
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 18001
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 18001
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_281
timestamp 18001
transform 1 0 26956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_289
timestamp 18001
transform 1 0 27692 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1636986456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1636986456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 18001
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1636986456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1636986456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1636986456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1636986456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 18001
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 18001
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1636986456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1636986456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1636986456
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1636986456
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 18001
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 18001
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1636986456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1636986456
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1636986456
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1636986456
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 18001
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 18001
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1636986456
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1636986456
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1636986456
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1636986456
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 18001
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 18001
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1636986456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1636986456
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1636986456
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_289
timestamp 18001
transform 1 0 27692 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1636986456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1636986456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1636986456
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1636986456
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 18001
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 18001
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1636986456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1636986456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1636986456
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1636986456
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 18001
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 18001
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_133
timestamp 1636986456
transform 1 0 13340 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_145
timestamp 1636986456
transform 1 0 14444 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_157
timestamp 18001
transform 1 0 15548 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_165
timestamp 18001
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1636986456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1636986456
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1636986456
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1636986456
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 18001
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 18001
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1636986456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1636986456
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1636986456
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1636986456
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 18001
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 18001
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_281
timestamp 18001
transform 1 0 26956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_289
timestamp 18001
transform 1 0 27692 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1636986456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1636986456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 18001
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1636986456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1636986456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1636986456
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1636986456
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 18001
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 18001
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1636986456
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_97
timestamp 18001
transform 1 0 10028 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_119
timestamp 1636986456
transform 1 0 12052 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_131
timestamp 18001
transform 1 0 13156 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 18001
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_162
timestamp 18001
transform 1 0 16008 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_185
timestamp 18001
transform 1 0 18124 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_193
timestamp 18001
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1636986456
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1636986456
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1636986456
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1636986456
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 18001
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 18001
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1636986456
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1636986456
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_277
timestamp 18001
transform 1 0 26588 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_285
timestamp 18001
transform 1 0 27324 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1636986456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1636986456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1636986456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_39
timestamp 18001
transform 1 0 4692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_47
timestamp 18001
transform 1 0 5428 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_57
timestamp 18001
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_64
timestamp 18001
transform 1 0 6992 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_72
timestamp 1636986456
transform 1 0 7728 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_84
timestamp 1636986456
transform 1 0 8832 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_96
timestamp 1636986456
transform 1 0 9936 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_108
timestamp 18001
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_113
timestamp 18001
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_129
timestamp 18001
transform 1 0 12972 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_135
timestamp 18001
transform 1 0 13524 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_143
timestamp 18001
transform 1 0 14260 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_156
timestamp 1636986456
transform 1 0 15456 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_169
timestamp 18001
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_197
timestamp 1636986456
transform 1 0 19228 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_209
timestamp 18001
transform 1 0 20332 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_218
timestamp 18001
transform 1 0 21160 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1636986456
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_240
timestamp 1636986456
transform 1 0 23184 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_252
timestamp 1636986456
transform 1 0 24288 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_264
timestamp 1636986456
transform 1 0 25392 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_276
timestamp 18001
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_281
timestamp 18001
transform 1 0 26956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_287
timestamp 18001
transform 1 0 27508 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1636986456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1636986456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 18001
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1636986456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_41
timestamp 18001
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_75
timestamp 18001
transform 1 0 8004 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 18001
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_93
timestamp 18001
transform 1 0 9660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_137
timestamp 18001
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_141
timestamp 18001
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_163
timestamp 18001
transform 1 0 16100 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_167
timestamp 18001
transform 1 0 16468 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_194
timestamp 18001
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_197
timestamp 18001
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_228
timestamp 18001
transform 1 0 22080 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1636986456
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1636986456
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1636986456
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_289
timestamp 18001
transform 1 0 27692 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1636986456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1636986456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_27
timestamp 18001
transform 1 0 3588 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_36
timestamp 1636986456
transform 1 0 4416 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_48
timestamp 18001
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_64
timestamp 1636986456
transform 1 0 6992 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_76
timestamp 18001
transform 1 0 8096 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_95
timestamp 18001
transform 1 0 9844 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_103
timestamp 18001
transform 1 0 10580 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 18001
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_119
timestamp 18001
transform 1 0 12052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_125
timestamp 18001
transform 1 0 12604 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_130
timestamp 1636986456
transform 1 0 13064 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_142
timestamp 18001
transform 1 0 14168 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_155
timestamp 18001
transform 1 0 15364 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 18001
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_169
timestamp 18001
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_254
timestamp 1636986456
transform 1 0 24472 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_266
timestamp 1636986456
transform 1 0 25576 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_278
timestamp 18001
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_281
timestamp 18001
transform 1 0 26956 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_289
timestamp 18001
transform 1 0 27692 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1636986456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1636986456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 18001
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_43
timestamp 1636986456
transform 1 0 5060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_55
timestamp 18001
transform 1 0 6164 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_61
timestamp 18001
transform 1 0 6716 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_69
timestamp 18001
transform 1 0 7452 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_77
timestamp 18001
transform 1 0 8188 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 18001
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_90
timestamp 1636986456
transform 1 0 9384 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_102
timestamp 18001
transform 1 0 10488 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_110
timestamp 18001
transform 1 0 11224 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_119
timestamp 18001
transform 1 0 12052 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_125
timestamp 18001
transform 1 0 12604 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 18001
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 18001
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1636986456
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_153
timestamp 18001
transform 1 0 15180 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_161
timestamp 18001
transform 1 0 15916 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_169
timestamp 18001
transform 1 0 16652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_176
timestamp 18001
transform 1 0 17296 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_194
timestamp 18001
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_205
timestamp 18001
transform 1 0 19964 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_229
timestamp 18001
transform 1 0 22172 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 18001
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_273
timestamp 1636986456
transform 1 0 26220 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_285
timestamp 18001
transform 1 0 27324 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1636986456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_15
timestamp 18001
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_32
timestamp 1636986456
transform 1 0 4048 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_44
timestamp 18001
transform 1 0 5152 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_49
timestamp 18001
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 18001
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_57
timestamp 18001
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_76
timestamp 18001
transform 1 0 8096 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_84
timestamp 18001
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_90
timestamp 18001
transform 1 0 9384 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_96
timestamp 18001
transform 1 0 9936 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_108
timestamp 18001
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_113
timestamp 18001
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_119
timestamp 1636986456
transform 1 0 12052 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_131
timestamp 1636986456
transform 1 0 13156 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_143
timestamp 1636986456
transform 1 0 14260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_155
timestamp 1636986456
transform 1 0 15364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 18001
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_178
timestamp 18001
transform 1 0 17480 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_187
timestamp 1636986456
transform 1 0 18308 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_199
timestamp 1636986456
transform 1 0 19412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_211
timestamp 1636986456
transform 1 0 20516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 18001
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1636986456
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_237
timestamp 18001
transform 1 0 22908 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_245
timestamp 18001
transform 1 0 23644 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_266
timestamp 1636986456
transform 1 0 25576 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_278
timestamp 18001
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_281
timestamp 18001
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_289
timestamp 18001
transform 1 0 27692 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1636986456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_15
timestamp 18001
transform 1 0 2484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp 18001
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_37
timestamp 18001
transform 1 0 4508 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_50
timestamp 1636986456
transform 1 0 5704 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_62
timestamp 1636986456
transform 1 0 6808 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 18001
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 18001
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1636986456
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_97
timestamp 18001
transform 1 0 10028 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_119
timestamp 18001
transform 1 0 12052 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_130
timestamp 18001
transform 1 0 13064 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 18001
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1636986456
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1636986456
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1636986456
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_177
timestamp 18001
transform 1 0 17388 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_185
timestamp 18001
transform 1 0 18124 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_190
timestamp 18001
transform 1 0 18584 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_202
timestamp 18001
transform 1 0 19688 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_210
timestamp 18001
transform 1 0 20424 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_217
timestamp 1636986456
transform 1 0 21068 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_229
timestamp 1636986456
transform 1 0 22172 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_241
timestamp 18001
transform 1 0 23276 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_249
timestamp 18001
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1636986456
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1636986456
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1636986456
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_289
timestamp 18001
transform 1 0 27692 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1636986456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1636986456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_27
timestamp 18001
transform 1 0 3588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_40
timestamp 18001
transform 1 0 4784 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_49
timestamp 18001
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 18001
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_57
timestamp 18001
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_65
timestamp 18001
transform 1 0 7084 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_71
timestamp 18001
transform 1 0 7636 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_84
timestamp 1636986456
transform 1 0 8832 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_96
timestamp 1636986456
transform 1 0 9936 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_108
timestamp 18001
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_113
timestamp 18001
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_121
timestamp 18001
transform 1 0 12236 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_133
timestamp 1636986456
transform 1 0 13340 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_145
timestamp 18001
transform 1 0 14444 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_149
timestamp 18001
transform 1 0 14812 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_160
timestamp 18001
transform 1 0 15824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 18001
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1636986456
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_181
timestamp 18001
transform 1 0 17756 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_189
timestamp 18001
transform 1 0 18492 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_196
timestamp 1636986456
transform 1 0 19136 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_208
timestamp 18001
transform 1 0 20240 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 18001
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1636986456
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1636986456
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_249
timestamp 18001
transform 1 0 24012 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_254
timestamp 1636986456
transform 1 0 24472 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_266
timestamp 1636986456
transform 1 0 25576 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_278
timestamp 18001
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_281
timestamp 18001
transform 1 0 26956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_289
timestamp 18001
transform 1 0 27692 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_3
timestamp 18001
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_9
timestamp 18001
transform 1 0 1932 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_17
timestamp 18001
transform 1 0 2668 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_25
timestamp 18001
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1636986456
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1636986456
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1636986456
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_65
timestamp 18001
transform 1 0 7084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_69
timestamp 18001
transform 1 0 7452 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_76
timestamp 18001
transform 1 0 8096 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_100
timestamp 18001
transform 1 0 10304 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_106
timestamp 18001
transform 1 0 10856 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_110
timestamp 1636986456
transform 1 0 11224 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_122
timestamp 18001
transform 1 0 12328 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_127
timestamp 18001
transform 1 0 12788 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_131
timestamp 18001
transform 1 0 13156 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_148
timestamp 18001
transform 1 0 14720 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_157
timestamp 18001
transform 1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_165
timestamp 18001
transform 1 0 16284 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_181
timestamp 18001
transform 1 0 17756 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_191
timestamp 18001
transform 1 0 18676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 18001
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_197
timestamp 18001
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_205
timestamp 18001
transform 1 0 19964 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_227
timestamp 1636986456
transform 1 0 21988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_239
timestamp 18001
transform 1 0 23092 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_250
timestamp 18001
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_273
timestamp 1636986456
transform 1 0 26220 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_285
timestamp 18001
transform 1 0 27324 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_3
timestamp 18001
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_16
timestamp 18001
transform 1 0 2576 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_29
timestamp 1636986456
transform 1 0 3772 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_41
timestamp 18001
transform 1 0 4876 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 18001
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_69
timestamp 18001
transform 1 0 7452 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_90
timestamp 1636986456
transform 1 0 9384 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_102
timestamp 18001
transform 1 0 10488 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_108
timestamp 18001
transform 1 0 11040 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_113
timestamp 18001
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_124
timestamp 18001
transform 1 0 12512 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_131
timestamp 18001
transform 1 0 13156 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_139
timestamp 18001
transform 1 0 13892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_196
timestamp 18001
transform 1 0 19136 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_202
timestamp 18001
transform 1 0 19688 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_222
timestamp 18001
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_225
timestamp 18001
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_233
timestamp 18001
transform 1 0 22540 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_264
timestamp 1636986456
transform 1 0 25392 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_276
timestamp 18001
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_281
timestamp 18001
transform 1 0 26956 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_289
timestamp 18001
transform 1 0 27692 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_3
timestamp 18001
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_18
timestamp 18001
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_26
timestamp 18001
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1636986456
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1636986456
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_53
timestamp 18001
transform 1 0 5980 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_68
timestamp 1636986456
transform 1 0 7360 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_80
timestamp 18001
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_85
timestamp 18001
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_93
timestamp 18001
transform 1 0 9660 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_127
timestamp 18001
transform 1 0 12788 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_131
timestamp 18001
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 18001
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_141
timestamp 18001
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_188
timestamp 18001
transform 1 0 18400 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_197
timestamp 18001
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_219
timestamp 1636986456
transform 1 0 21252 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_231
timestamp 18001
transform 1 0 22356 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_250
timestamp 18001
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_253
timestamp 18001
transform 1 0 24380 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_260
timestamp 1636986456
transform 1 0 25024 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_272
timestamp 1636986456
transform 1 0 26128 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_284
timestamp 18001
transform 1 0 27232 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_290
timestamp 18001
transform 1 0 27784 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_9
timestamp 18001
transform 1 0 1932 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_17
timestamp 18001
transform 1 0 2668 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_29
timestamp 18001
transform 1 0 3772 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_35
timestamp 18001
transform 1 0 4324 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_46
timestamp 18001
transform 1 0 5336 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 18001
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1636986456
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_69
timestamp 18001
transform 1 0 7452 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_73
timestamp 1636986456
transform 1 0 7820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_85
timestamp 1636986456
transform 1 0 8924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_97
timestamp 18001
transform 1 0 10028 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_105
timestamp 18001
transform 1 0 10764 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_126
timestamp 1636986456
transform 1 0 12696 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_138
timestamp 1636986456
transform 1 0 13800 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_150
timestamp 18001
transform 1 0 14904 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_180
timestamp 18001
transform 1 0 17664 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_188
timestamp 18001
transform 1 0 18400 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 18001
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1636986456
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_237
timestamp 18001
transform 1 0 22908 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_246
timestamp 1636986456
transform 1 0 23736 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_258
timestamp 1636986456
transform 1 0 24840 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_270
timestamp 18001
transform 1 0 25944 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_278
timestamp 18001
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_281
timestamp 18001
transform 1 0 26956 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_289
timestamp 18001
transform 1 0 27692 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1636986456
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_15
timestamp 18001
transform 1 0 2484 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_32
timestamp 18001
transform 1 0 4048 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_44
timestamp 18001
transform 1 0 5152 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_50
timestamp 18001
transform 1 0 5704 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_80
timestamp 18001
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1636986456
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1636986456
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_115
timestamp 18001
transform 1 0 11684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_131
timestamp 18001
transform 1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 18001
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1636986456
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_153
timestamp 18001
transform 1 0 15180 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_161
timestamp 18001
transform 1 0 15916 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_176
timestamp 18001
transform 1 0 17296 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_184
timestamp 18001
transform 1 0 18032 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_188
timestamp 18001
transform 1 0 18400 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_215
timestamp 18001
transform 1 0 20884 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_224
timestamp 1636986456
transform 1 0 21712 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_236
timestamp 1636986456
transform 1 0 22816 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_248
timestamp 18001
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1636986456
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1636986456
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1636986456
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_289
timestamp 18001
transform 1 0 27692 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_3
timestamp 18001
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_14
timestamp 1636986456
transform 1 0 2392 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_26
timestamp 1636986456
transform 1 0 3496 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_38
timestamp 18001
transform 1 0 4600 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_42
timestamp 18001
transform 1 0 4968 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_57
timestamp 18001
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_61
timestamp 1636986456
transform 1 0 6716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_73
timestamp 18001
transform 1 0 7820 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_94
timestamp 1636986456
transform 1 0 9752 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_106
timestamp 18001
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_113
timestamp 18001
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1636986456
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1636986456
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_149
timestamp 18001
transform 1 0 14812 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_162
timestamp 18001
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1636986456
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_185
timestamp 18001
transform 1 0 18124 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_189
timestamp 18001
transform 1 0 18492 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_220
timestamp 18001
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_230
timestamp 18001
transform 1 0 22264 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_238
timestamp 18001
transform 1 0 23000 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_247
timestamp 1636986456
transform 1 0 23828 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_259
timestamp 1636986456
transform 1 0 24932 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_271
timestamp 18001
transform 1 0 26036 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 18001
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_281
timestamp 18001
transform 1 0 26956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_289
timestamp 18001
transform 1 0 27692 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_3
timestamp 18001
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_16
timestamp 1636986456
transform 1 0 2576 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1636986456
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1636986456
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_53
timestamp 18001
transform 1 0 5980 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_61
timestamp 18001
transform 1 0 6716 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_74
timestamp 18001
transform 1 0 7912 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_98
timestamp 1636986456
transform 1 0 10120 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_110
timestamp 18001
transform 1 0 11224 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_118
timestamp 18001
transform 1 0 11960 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_130
timestamp 18001
transform 1 0 13064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 18001
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_167
timestamp 18001
transform 1 0 16468 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_175
timestamp 18001
transform 1 0 17204 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_183
timestamp 1636986456
transform 1 0 17940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 18001
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_197
timestamp 18001
transform 1 0 19228 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_212
timestamp 1636986456
transform 1 0 20608 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_224
timestamp 18001
transform 1 0 21712 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_231
timestamp 18001
transform 1 0 22356 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_247
timestamp 18001
transform 1 0 23828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 18001
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_260
timestamp 1636986456
transform 1 0 25024 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_272
timestamp 1636986456
transform 1 0 26128 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_284
timestamp 18001
transform 1 0 27232 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_290
timestamp 18001
transform 1 0 27784 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_14
timestamp 18001
transform 1 0 2392 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_25
timestamp 18001
transform 1 0 3404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_45
timestamp 18001
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_53
timestamp 18001
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_64
timestamp 1636986456
transform 1 0 6992 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_76
timestamp 18001
transform 1 0 8096 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_86
timestamp 1636986456
transform 1 0 9016 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_98
timestamp 18001
transform 1 0 10120 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_102
timestamp 18001
transform 1 0 10488 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_106
timestamp 18001
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_116
timestamp 18001
transform 1 0 11776 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_127
timestamp 1636986456
transform 1 0 12788 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_139
timestamp 18001
transform 1 0 13892 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_143
timestamp 18001
transform 1 0 14260 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_153
timestamp 18001
transform 1 0 15180 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 18001
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 18001
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1636986456
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_181
timestamp 18001
transform 1 0 17756 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_191
timestamp 1636986456
transform 1 0 18676 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_203
timestamp 1636986456
transform 1 0 19780 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_215
timestamp 18001
transform 1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 18001
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_270
timestamp 18001
transform 1 0 25944 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_278
timestamp 18001
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_281
timestamp 18001
transform 1 0 26956 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_3
timestamp 18001
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_9
timestamp 18001
transform 1 0 1932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_17
timestamp 18001
transform 1 0 2668 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_25
timestamp 18001
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_36
timestamp 18001
transform 1 0 4416 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_44
timestamp 18001
transform 1 0 5152 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_51
timestamp 18001
transform 1 0 5796 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_67
timestamp 1636986456
transform 1 0 7268 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_79
timestamp 18001
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 18001
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1636986456
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_97
timestamp 18001
transform 1 0 10028 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_105
timestamp 18001
transform 1 0 10764 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_135
timestamp 18001
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 18001
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_141
timestamp 18001
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_147
timestamp 18001
transform 1 0 14628 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_154
timestamp 1636986456
transform 1 0 15272 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_166
timestamp 18001
transform 1 0 16376 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_170
timestamp 18001
transform 1 0 16744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_181
timestamp 18001
transform 1 0 17756 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_191
timestamp 18001
transform 1 0 18676 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 18001
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_204
timestamp 18001
transform 1 0 19872 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_219
timestamp 18001
transform 1 0 21252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_225
timestamp 18001
transform 1 0 21804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_239
timestamp 18001
transform 1 0 23092 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 18001
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_259
timestamp 1636986456
transform 1 0 24932 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_271
timestamp 1636986456
transform 1 0 26036 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_283
timestamp 18001
transform 1 0 27140 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1636986456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_18
timestamp 18001
transform 1 0 2760 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_36
timestamp 18001
transform 1 0 4416 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 18001
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_72
timestamp 18001
transform 1 0 7728 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_76
timestamp 18001
transform 1 0 8096 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_109
timestamp 18001
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_113
timestamp 18001
transform 1 0 11500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_130
timestamp 18001
transform 1 0 13064 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_138
timestamp 18001
transform 1 0 13800 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_148
timestamp 1636986456
transform 1 0 14720 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_160
timestamp 18001
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_169
timestamp 18001
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1636986456
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_237
timestamp 18001
transform 1 0 22908 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_244
timestamp 18001
transform 1 0 23552 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_250
timestamp 1636986456
transform 1 0 24104 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_262
timestamp 1636986456
transform 1 0 25208 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_274
timestamp 18001
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_281
timestamp 18001
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_289
timestamp 18001
transform 1 0 27692 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1636986456
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1636986456
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 18001
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_29
timestamp 18001
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_40
timestamp 1636986456
transform 1 0 4784 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_52
timestamp 18001
transform 1 0 5888 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_60
timestamp 18001
transform 1 0 6624 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_85
timestamp 18001
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_109
timestamp 18001
transform 1 0 11132 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_113
timestamp 18001
transform 1 0 11500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1636986456
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 18001
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 18001
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1636986456
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_153
timestamp 18001
transform 1 0 15180 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_161
timestamp 18001
transform 1 0 15916 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_169
timestamp 18001
transform 1 0 16652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_197
timestamp 18001
transform 1 0 19228 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_209
timestamp 18001
transform 1 0 20332 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_218
timestamp 1636986456
transform 1 0 21160 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_230
timestamp 18001
transform 1 0 22264 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_238
timestamp 18001
transform 1 0 23000 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_249
timestamp 18001
transform 1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_258
timestamp 1636986456
transform 1 0 24840 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_270
timestamp 1636986456
transform 1 0 25944 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_282
timestamp 18001
transform 1 0 27048 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_290
timestamp 18001
transform 1 0 27784 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_9
timestamp 18001
transform 1 0 1932 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_17
timestamp 18001
transform 1 0 2668 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_25
timestamp 18001
transform 1 0 3404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_47
timestamp 18001
transform 1 0 5428 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_52
timestamp 18001
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_57
timestamp 18001
transform 1 0 6348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_102
timestamp 18001
transform 1 0 10488 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_110
timestamp 18001
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_113
timestamp 18001
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_117
timestamp 18001
transform 1 0 11868 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_126
timestamp 1636986456
transform 1 0 12696 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_156
timestamp 1636986456
transform 1 0 15456 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_178
timestamp 18001
transform 1 0 17480 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_186
timestamp 18001
transform 1 0 18216 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_190
timestamp 18001
transform 1 0 18584 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_194
timestamp 18001
transform 1 0 18952 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_206
timestamp 1636986456
transform 1 0 20056 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_218
timestamp 18001
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1636986456
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_237
timestamp 18001
transform 1 0 22908 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_262
timestamp 1636986456
transform 1 0 25208 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_274
timestamp 18001
transform 1 0 26312 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_281
timestamp 18001
transform 1 0 26956 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_289
timestamp 18001
transform 1 0 27692 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_3
timestamp 18001
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_11
timestamp 18001
transform 1 0 2116 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 18001
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_29
timestamp 18001
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_35
timestamp 18001
transform 1 0 4324 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_80
timestamp 18001
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_107
timestamp 1636986456
transform 1 0 10948 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_134
timestamp 18001
transform 1 0 13432 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_164
timestamp 1636986456
transform 1 0 16192 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_176
timestamp 1636986456
transform 1 0 17296 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_188
timestamp 18001
transform 1 0 18400 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_197
timestamp 18001
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_203
timestamp 18001
transform 1 0 19780 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 18001
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_253
timestamp 18001
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_261
timestamp 1636986456
transform 1 0 25116 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_273
timestamp 1636986456
transform 1 0 26220 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_285
timestamp 18001
transform 1 0 27324 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_3
timestamp 18001
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_16
timestamp 18001
transform 1 0 2576 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_24
timestamp 18001
transform 1 0 3312 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_41
timestamp 1636986456
transform 1 0 4876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_53
timestamp 18001
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1636986456
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_69
timestamp 18001
transform 1 0 7452 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_74
timestamp 18001
transform 1 0 7912 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_82
timestamp 18001
transform 1 0 8648 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_113
timestamp 18001
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_139
timestamp 18001
transform 1 0 13892 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_147
timestamp 18001
transform 1 0 14628 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_155
timestamp 18001
transform 1 0 15364 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_164
timestamp 18001
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_169
timestamp 18001
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_174
timestamp 1636986456
transform 1 0 17112 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_186
timestamp 18001
transform 1 0 18216 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_194
timestamp 18001
transform 1 0 18952 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_211
timestamp 18001
transform 1 0 20516 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_217
timestamp 18001
transform 1 0 21068 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_221
timestamp 18001
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_225
timestamp 18001
transform 1 0 21804 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_236
timestamp 18001
transform 1 0 22816 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_246
timestamp 18001
transform 1 0 23736 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_254
timestamp 18001
transform 1 0 24472 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_263
timestamp 1636986456
transform 1 0 25300 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_275
timestamp 18001
transform 1 0 26404 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 18001
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_281
timestamp 18001
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_289
timestamp 18001
transform 1 0 27692 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_26
timestamp 18001
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1636986456
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1636986456
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_53
timestamp 18001
transform 1 0 5980 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_81
timestamp 18001
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_85
timestamp 18001
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_104
timestamp 1636986456
transform 1 0 10672 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_116
timestamp 18001
transform 1 0 11776 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_123
timestamp 1636986456
transform 1 0 12420 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_135
timestamp 18001
transform 1 0 13524 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 18001
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_141
timestamp 18001
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_155
timestamp 18001
transform 1 0 15364 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_163
timestamp 18001
transform 1 0 16100 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1636986456
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_209
timestamp 18001
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1636986456
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1636986456
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 1636986456
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_289
timestamp 18001
transform 1 0 27692 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_15
timestamp 18001
transform 1 0 2484 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_26
timestamp 1636986456
transform 1 0 3496 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_38
timestamp 18001
transform 1 0 4600 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_44
timestamp 1636986456
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_60
timestamp 18001
transform 1 0 6624 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_70
timestamp 1636986456
transform 1 0 7544 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_82
timestamp 18001
transform 1 0 8648 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_101
timestamp 18001
transform 1 0 10396 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_109
timestamp 18001
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_113
timestamp 18001
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_117
timestamp 18001
transform 1 0 11868 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_129
timestamp 18001
transform 1 0 12972 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_137
timestamp 18001
transform 1 0 13708 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_143
timestamp 18001
transform 1 0 14260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_154
timestamp 18001
transform 1 0 15272 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_160
timestamp 18001
transform 1 0 15824 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_166
timestamp 18001
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_169
timestamp 18001
transform 1 0 16652 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_214
timestamp 18001
transform 1 0 20792 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_222
timestamp 18001
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_232
timestamp 18001
transform 1 0 22448 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_239
timestamp 1636986456
transform 1 0 23092 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_251
timestamp 1636986456
transform 1 0 24196 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_263
timestamp 1636986456
transform 1 0 25300 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_275
timestamp 18001
transform 1 0 26404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 18001
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_281
timestamp 18001
transform 1 0 26956 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_289
timestamp 18001
transform 1 0 27692 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1636986456
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1636986456
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 18001
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_29
timestamp 18001
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_37
timestamp 18001
transform 1 0 4508 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_73
timestamp 18001
transform 1 0 7820 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_95
timestamp 1636986456
transform 1 0 9844 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_107
timestamp 1636986456
transform 1 0 10948 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_119
timestamp 18001
transform 1 0 12052 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_132
timestamp 18001
transform 1 0 13248 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_136
timestamp 18001
transform 1 0 13616 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_149
timestamp 1636986456
transform 1 0 14812 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_161
timestamp 1636986456
transform 1 0 15916 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_173
timestamp 18001
transform 1 0 17020 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 18001
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_197
timestamp 18001
transform 1 0 19228 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_205
timestamp 18001
transform 1 0 19964 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_226
timestamp 18001
transform 1 0 21896 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1636986456
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1636986456
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1636986456
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_289
timestamp 18001
transform 1 0 27692 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1636986456
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_15
timestamp 18001
transform 1 0 2484 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_34
timestamp 18001
transform 1 0 4232 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_60
timestamp 1636986456
transform 1 0 6624 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_72
timestamp 18001
transform 1 0 7728 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_100
timestamp 1636986456
transform 1 0 10304 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_113
timestamp 18001
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_121
timestamp 18001
transform 1 0 12236 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_131
timestamp 1636986456
transform 1 0 13156 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_143
timestamp 1636986456
transform 1 0 14260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_155
timestamp 1636986456
transform 1 0 15364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 18001
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1636986456
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_181
timestamp 18001
transform 1 0 17756 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_187
timestamp 18001
transform 1 0 18308 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_215
timestamp 18001
transform 1 0 20884 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 18001
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_234
timestamp 1636986456
transform 1 0 22632 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_246
timestamp 1636986456
transform 1 0 23736 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_258
timestamp 1636986456
transform 1 0 24840 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_270
timestamp 18001
transform 1 0 25944 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_278
timestamp 18001
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_281
timestamp 18001
transform 1 0 26956 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_289
timestamp 18001
transform 1 0 27692 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_19
timestamp 18001
transform 1 0 2852 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_29
timestamp 18001
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_49
timestamp 1636986456
transform 1 0 5612 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_61
timestamp 18001
transform 1 0 6716 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_76
timestamp 18001
transform 1 0 8096 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1636986456
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_97
timestamp 18001
transform 1 0 10028 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_128
timestamp 18001
transform 1 0 12880 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 18001
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_148
timestamp 1636986456
transform 1 0 14720 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_160
timestamp 1636986456
transform 1 0 15824 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_172
timestamp 1636986456
transform 1 0 16928 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_184
timestamp 1636986456
transform 1 0 18032 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_197
timestamp 18001
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_205
timestamp 18001
transform 1 0 19964 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_213
timestamp 18001
transform 1 0 20700 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_220
timestamp 18001
transform 1 0 21344 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_235
timestamp 1636986456
transform 1 0 22724 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_247
timestamp 18001
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 18001
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1636986456
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_265
timestamp 18001
transform 1 0 25484 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_3
timestamp 18001
transform 1 0 1380 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_9
timestamp 18001
transform 1 0 1932 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_29
timestamp 1636986456
transform 1 0 3772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_41
timestamp 1636986456
transform 1 0 4876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 18001
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_57
timestamp 18001
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_64
timestamp 18001
transform 1 0 6992 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1636986456
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 1636986456
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_126
timestamp 18001
transform 1 0 12696 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_148
timestamp 18001
transform 1 0 14720 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_160
timestamp 18001
transform 1 0 15824 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_185
timestamp 18001
transform 1 0 18124 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_191
timestamp 18001
transform 1 0 18676 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_205
timestamp 18001
transform 1 0 19964 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_245
timestamp 1636986456
transform 1 0 23644 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_257
timestamp 18001
transform 1 0 24748 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_269
timestamp 18001
transform 1 0 25852 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_277
timestamp 18001
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_281
timestamp 18001
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_289
timestamp 18001
transform 1 0 27692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_3
timestamp 18001
transform 1 0 1380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_19
timestamp 18001
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 18001
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1636986456
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_41
timestamp 18001
transform 1 0 4876 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_82
timestamp 18001
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1636986456
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_97
timestamp 18001
transform 1 0 10028 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_105
timestamp 18001
transform 1 0 10764 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_123
timestamp 18001
transform 1 0 12420 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_131
timestamp 18001
transform 1 0 13156 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_137
timestamp 18001
transform 1 0 13708 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_212
timestamp 18001
transform 1 0 20608 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_220
timestamp 18001
transform 1 0 21344 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_235
timestamp 1636986456
transform 1 0 22724 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_247
timestamp 18001
transform 1 0 23828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 18001
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_253
timestamp 18001
transform 1 0 24380 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_276
timestamp 1636986456
transform 1 0 26496 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_288
timestamp 18001
transform 1 0 27600 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_20
timestamp 18001
transform 1 0 2944 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_39
timestamp 18001
transform 1 0 4692 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_44
timestamp 18001
transform 1 0 5152 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_54
timestamp 18001
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_57
timestamp 18001
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_65
timestamp 18001
transform 1 0 7084 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_89
timestamp 1636986456
transform 1 0 9292 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_101
timestamp 18001
transform 1 0 10396 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_109
timestamp 18001
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1636986456
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 1636986456
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_137
timestamp 18001
transform 1 0 13708 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_160
timestamp 18001
transform 1 0 15824 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_175
timestamp 18001
transform 1 0 17204 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 1636986456
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_217
timestamp 18001
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 18001
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1636986456
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 1636986456
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_249
timestamp 18001
transform 1 0 24012 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_285
timestamp 18001
transform 1 0 27324 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_25
timestamp 18001
transform 1 0 3404 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_29
timestamp 18001
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_34
timestamp 18001
transform 1 0 4232 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_60
timestamp 1636986456
transform 1 0 6624 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_72
timestamp 1636986456
transform 1 0 7728 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_85
timestamp 18001
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_89
timestamp 18001
transform 1 0 9292 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_106
timestamp 18001
transform 1 0 10856 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_130
timestamp 18001
transform 1 0 13064 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_138
timestamp 18001
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_141
timestamp 18001
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 1636986456
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_165
timestamp 18001
transform 1 0 16284 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_171
timestamp 18001
transform 1 0 16836 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_177
timestamp 1636986456
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_189
timestamp 18001
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 18001
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 1636986456
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_209
timestamp 18001
transform 1 0 20332 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 1636986456
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_233
timestamp 1636986456
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_245
timestamp 18001
transform 1 0 23644 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_253
timestamp 18001
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_261
timestamp 18001
transform 1 0 25116 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_276
timestamp 18001
transform 1 0 26496 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_284
timestamp 18001
transform 1 0 27232 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_36
timestamp 1636986456
transform 1 0 4416 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_48
timestamp 18001
transform 1 0 5520 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_57
timestamp 18001
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_64
timestamp 18001
transform 1 0 6992 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_68
timestamp 18001
transform 1 0 7360 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_72
timestamp 18001
transform 1 0 7728 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_77
timestamp 18001
transform 1 0 8188 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_83
timestamp 18001
transform 1 0 8740 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_89
timestamp 18001
transform 1 0 9292 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_98
timestamp 1636986456
transform 1 0 10120 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_110
timestamp 18001
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_113
timestamp 18001
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_121
timestamp 18001
transform 1 0 12236 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_130
timestamp 1636986456
transform 1 0 13064 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_142
timestamp 1636986456
transform 1 0 14168 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_154
timestamp 1636986456
transform 1 0 15272 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_166
timestamp 18001
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 1636986456
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_181
timestamp 18001
transform 1 0 17756 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_203
timestamp 18001
transform 1 0 19780 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_210
timestamp 1636986456
transform 1 0 20424 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_222
timestamp 18001
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_225
timestamp 18001
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_233
timestamp 1636986456
transform 1 0 22540 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_245
timestamp 1636986456
transform 1 0 23644 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_268
timestamp 18001
transform 1 0 25760 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_275
timestamp 18001
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 18001
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_286
timestamp 18001
transform 1 0 27416 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_7
timestamp 18001
transform 1 0 1748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_11
timestamp 18001
transform 1 0 2116 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_24
timestamp 18001
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1636986456
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_85
timestamp 18001
transform 1 0 8924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_91
timestamp 18001
transform 1 0 9476 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_95
timestamp 18001
transform 1 0 9844 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_113
timestamp 18001
transform 1 0 11500 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_119
timestamp 18001
transform 1 0 12052 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_130
timestamp 18001
transform 1 0 13064 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_138
timestamp 18001
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_148
timestamp 1636986456
transform 1 0 14720 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_160
timestamp 18001
transform 1 0 15824 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_168
timestamp 18001
transform 1 0 16560 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_174
timestamp 1636986456
transform 1 0 17112 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_186
timestamp 18001
transform 1 0 18216 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_194
timestamp 18001
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_203
timestamp 1636986456
transform 1 0 19780 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_215
timestamp 18001
transform 1 0 20884 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_223
timestamp 18001
transform 1 0 21620 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_240
timestamp 18001
transform 1 0 23184 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 18001
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_261
timestamp 18001
transform 1 0 25116 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_267
timestamp 18001
transform 1 0 25668 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_275
timestamp 18001
transform 1 0 26404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_289
timestamp 18001
transform 1 0 27692 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_3
timestamp 18001
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_19
timestamp 1636986456
transform 1 0 2852 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_31
timestamp 18001
transform 1 0 3956 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_45
timestamp 18001
transform 1 0 5244 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_57
timestamp 18001
transform 1 0 6348 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_72
timestamp 1636986456
transform 1 0 7728 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_84
timestamp 18001
transform 1 0 8832 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_95
timestamp 18001
transform 1 0 9844 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_102
timestamp 18001
transform 1 0 10488 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_110
timestamp 18001
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_113
timestamp 18001
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_152
timestamp 18001
transform 1 0 15088 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_160
timestamp 18001
transform 1 0 15824 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_164
timestamp 18001
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_169
timestamp 18001
transform 1 0 16652 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_173
timestamp 18001
transform 1 0 17020 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_198
timestamp 18001
transform 1 0 19320 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_245
timestamp 18001
transform 1 0 23644 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_274
timestamp 18001
transform 1 0 26312 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_281
timestamp 18001
transform 1 0 26956 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_29
timestamp 18001
transform 1 0 3772 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1636986456
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_65
timestamp 18001
transform 1 0 7084 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_74
timestamp 18001
transform 1 0 7912 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_82
timestamp 18001
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_85
timestamp 18001
transform 1 0 8924 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_106
timestamp 18001
transform 1 0 10856 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_130
timestamp 18001
transform 1 0 13064 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_138
timestamp 18001
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_144
timestamp 18001
transform 1 0 14352 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_157
timestamp 18001
transform 1 0 15548 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_186
timestamp 18001
transform 1 0 18216 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_194
timestamp 18001
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_218
timestamp 18001
transform 1 0 21160 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_248
timestamp 18001
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_253
timestamp 18001
transform 1 0 24380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_262
timestamp 18001
transform 1 0 25208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_266
timestamp 18001
transform 1 0 25576 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_283
timestamp 18001
transform 1 0 27140 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_6
timestamp 18001
transform 1 0 1656 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_14
timestamp 18001
transform 1 0 2392 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_34
timestamp 18001
transform 1 0 4232 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_39
timestamp 18001
transform 1 0 4692 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_49
timestamp 18001
transform 1 0 5612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 18001
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1636986456
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_69
timestamp 18001
transform 1 0 7452 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_91
timestamp 18001
transform 1 0 9476 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_97
timestamp 18001
transform 1 0 10028 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 18001
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_113
timestamp 18001
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_121
timestamp 1636986456
transform 1 0 12236 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_133
timestamp 1636986456
transform 1 0 13340 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_145
timestamp 18001
transform 1 0 14444 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 18001
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_182
timestamp 1636986456
transform 1 0 17848 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_194
timestamp 1636986456
transform 1 0 18952 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_206
timestamp 1636986456
transform 1 0 20056 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_218
timestamp 18001
transform 1 0 21160 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_241
timestamp 1636986456
transform 1 0 23276 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_253
timestamp 1636986456
transform 1 0 24380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_265
timestamp 18001
transform 1 0 25484 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_278
timestamp 18001
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_286
timestamp 18001
transform 1 0 27416 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1636986456
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1636986456
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 18001
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1636986456
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1636986456
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1636986456
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1636986456
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 18001
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 18001
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_85
timestamp 18001
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_96
timestamp 18001
transform 1 0 9936 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_107
timestamp 1636986456
transform 1 0 10948 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_119
timestamp 18001
transform 1 0 12052 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_131
timestamp 18001
transform 1 0 13156 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 18001
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1636986456
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_153
timestamp 18001
transform 1 0 15180 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_162
timestamp 18001
transform 1 0 16008 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_175
timestamp 1636986456
transform 1 0 17204 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_187
timestamp 18001
transform 1 0 18308 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 18001
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 1636986456
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_209
timestamp 1636986456
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_221
timestamp 18001
transform 1 0 21436 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_225
timestamp 18001
transform 1 0 21804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_230
timestamp 1636986456
transform 1 0 22264 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_242
timestamp 18001
transform 1 0 23368 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_250
timestamp 18001
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1636986456
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_265
timestamp 18001
transform 1 0 25484 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_277
timestamp 18001
transform 1 0 26588 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_285
timestamp 18001
transform 1 0 27324 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_3
timestamp 18001
transform 1 0 1380 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_11
timestamp 18001
transform 1 0 2116 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1636986456
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1636986456
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 18001
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 18001
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_57
timestamp 18001
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_72
timestamp 18001
transform 1 0 7728 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_85
timestamp 1636986456
transform 1 0 8924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_97
timestamp 1636986456
transform 1 0 10028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_109
timestamp 18001
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_113
timestamp 18001
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_129
timestamp 1636986456
transform 1 0 12972 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_141
timestamp 1636986456
transform 1 0 14076 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_153
timestamp 1636986456
transform 1 0 15180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_165
timestamp 18001
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1636986456
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 1636986456
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_193
timestamp 1636986456
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_205
timestamp 18001
transform 1 0 19964 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_209
timestamp 18001
transform 1 0 20332 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_213
timestamp 18001
transform 1 0 20700 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_221
timestamp 18001
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_225
timestamp 18001
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_233
timestamp 18001
transform 1 0 22540 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_239
timestamp 1636986456
transform 1 0 23092 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_251
timestamp 18001
transform 1 0 24196 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_259
timestamp 18001
transform 1 0 24932 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_269
timestamp 18001
transform 1 0 25852 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_278
timestamp 18001
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_281
timestamp 18001
transform 1 0 26956 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_289
timestamp 18001
transform 1 0 27692 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_3
timestamp 18001
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_26
timestamp 18001
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_29
timestamp 18001
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_37
timestamp 18001
transform 1 0 4508 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_41
timestamp 18001
transform 1 0 4876 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_49
timestamp 18001
transform 1 0 5612 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1636986456
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 18001
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 18001
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_85
timestamp 18001
transform 1 0 8924 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_96
timestamp 18001
transform 1 0 9936 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_102
timestamp 18001
transform 1 0 10488 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_107
timestamp 18001
transform 1 0 10948 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_115
timestamp 18001
transform 1 0 11684 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_134
timestamp 18001
transform 1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1636986456
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1636986456
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 1636986456
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 1636986456
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 18001
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 18001
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_197
timestamp 18001
transform 1 0 19228 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_201
timestamp 18001
transform 1 0 19596 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_214
timestamp 1636986456
transform 1 0 20792 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_226
timestamp 18001
transform 1 0 21896 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_233
timestamp 18001
transform 1 0 22540 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 18001
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 18001
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_253
timestamp 18001
transform 1 0 24380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_265
timestamp 18001
transform 1 0 25484 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_283
timestamp 18001
transform 1 0 27140 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_3
timestamp 18001
transform 1 0 1380 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_11
timestamp 18001
transform 1 0 2116 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_19
timestamp 18001
transform 1 0 2852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_54
timestamp 18001
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_61
timestamp 18001
transform 1 0 6716 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_78
timestamp 1636986456
transform 1 0 8280 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_90
timestamp 18001
transform 1 0 9384 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_96
timestamp 18001
transform 1 0 9936 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 18001
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_130
timestamp 1636986456
transform 1 0 13064 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_142
timestamp 1636986456
transform 1 0 14168 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_154
timestamp 1636986456
transform 1 0 15272 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_166
timestamp 18001
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1636986456
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_184
timestamp 18001
transform 1 0 18032 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_189
timestamp 18001
transform 1 0 18492 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_198
timestamp 18001
transform 1 0 19320 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_210
timestamp 18001
transform 1 0 20424 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_225
timestamp 18001
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_246
timestamp 18001
transform 1 0 23736 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_250
timestamp 18001
transform 1 0 24104 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_262
timestamp 18001
transform 1 0 25208 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_266
timestamp 18001
transform 1 0 25576 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_276
timestamp 18001
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_281
timestamp 18001
transform 1 0 26956 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1636986456
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1636986456
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 18001
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_32
timestamp 18001
transform 1 0 4048 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_52
timestamp 18001
transform 1 0 5888 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_57
timestamp 18001
transform 1 0 6348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_76
timestamp 18001
transform 1 0 8096 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_85
timestamp 18001
transform 1 0 8924 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_95
timestamp 18001
transform 1 0 9844 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_129
timestamp 18001
transform 1 0 12972 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_137
timestamp 18001
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1636986456
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 1636986456
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_165
timestamp 18001
transform 1 0 16284 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_173
timestamp 18001
transform 1 0 17020 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_187
timestamp 18001
transform 1 0 18308 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_229
timestamp 18001
transform 1 0 22172 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_244
timestamp 18001
transform 1 0 23552 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_248
timestamp 18001
transform 1 0 23920 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_277
timestamp 18001
transform 1 0 26588 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1636986456
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1636986456
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1636986456
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1636986456
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 18001
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 18001
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_57
timestamp 18001
transform 1 0 6348 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_61
timestamp 18001
transform 1 0 6716 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_65
timestamp 1636986456
transform 1 0 7084 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_77
timestamp 1636986456
transform 1 0 8188 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_89
timestamp 1636986456
transform 1 0 9292 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_101
timestamp 18001
transform 1 0 10396 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 18001
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_118
timestamp 1636986456
transform 1 0 11960 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_130
timestamp 1636986456
transform 1 0 13064 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_142
timestamp 1636986456
transform 1 0 14168 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_154
timestamp 1636986456
transform 1 0 15272 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_166
timestamp 18001
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1636986456
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_181
timestamp 18001
transform 1 0 17756 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_186
timestamp 18001
transform 1 0 18216 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_194
timestamp 18001
transform 1 0 18952 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_212
timestamp 18001
transform 1 0 20608 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_219
timestamp 18001
transform 1 0 21252 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 18001
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_232
timestamp 1636986456
transform 1 0 22448 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_244
timestamp 1636986456
transform 1 0 23552 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_264
timestamp 18001
transform 1 0 25392 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_268
timestamp 18001
transform 1 0 25760 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_272
timestamp 18001
transform 1 0 26128 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_281
timestamp 18001
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_289
timestamp 18001
transform 1 0 27692 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1636986456
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1636986456
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 18001
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1636986456
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1636986456
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_53
timestamp 18001
transform 1 0 5980 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_57
timestamp 1636986456
transform 1 0 6348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_69
timestamp 1636986456
transform 1 0 7452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_81
timestamp 18001
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1636986456
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 1636986456
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_109
timestamp 18001
transform 1 0 11132 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_113
timestamp 1636986456
transform 1 0 11500 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_125
timestamp 18001
transform 1 0 12604 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_141
timestamp 18001
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_149
timestamp 18001
transform 1 0 14812 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_156
timestamp 18001
transform 1 0 15456 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_163
timestamp 18001
transform 1 0 16100 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_167
timestamp 18001
transform 1 0 16468 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_193
timestamp 18001
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_221
timestamp 18001
transform 1 0 21436 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_249
timestamp 18001
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_277
timestamp 18001
transform 1 0 26588 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_287
timestamp 18001
transform 1 0 27508 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 18001
transform 1 0 27600 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 18001
transform -1 0 27876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 18001
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 18001
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 18001
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 18001
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 18001
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 18001
transform 1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input9
timestamp 18001
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input10
timestamp 18001
transform 1 0 1380 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input11
timestamp 18001
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input12
timestamp 18001
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input13
timestamp 18001
transform 1 0 1380 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input14
timestamp 18001
transform 1 0 2852 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input15
timestamp 18001
transform 1 0 2392 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 18001
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 18001
transform -1 0 27876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 18001
transform -1 0 27876 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 18001
transform 1 0 27508 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 18001
transform 1 0 23460 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 18001
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 18001
transform -1 0 13432 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 18001
transform -1 0 14812 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 18001
transform 1 0 24380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 18001
transform -1 0 17204 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 18001
transform 1 0 27508 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 18001
transform 1 0 22908 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 18001
transform 1 0 17204 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 18001
transform 1 0 25484 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 18001
transform 1 0 27508 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 18001
transform 1 0 20884 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 18001
transform 1 0 18308 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output33
timestamp 18001
transform 1 0 22356 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output34
timestamp 18001
transform 1 0 27324 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 18001
transform -1 0 15456 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 18001
transform -1 0 26588 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 18001
transform 1 0 27508 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output38
timestamp 18001
transform 1 0 26956 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 18001
transform 1 0 20332 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 18001
transform -1 0 20332 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 18001
transform 1 0 19228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 18001
transform 1 0 27508 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 18001
transform 1 0 27508 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 18001
transform 1 0 27508 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 18001
transform 1 0 27508 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output46
timestamp 18001
transform 1 0 26772 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output47
timestamp 18001
transform -1 0 16100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output48
timestamp 18001
transform -1 0 13984 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output49
timestamp 18001
transform 1 0 21804 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output50
timestamp 18001
transform 1 0 24932 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output51
timestamp 18001
transform -1 0 18308 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output52
timestamp 18001
transform 1 0 27140 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_49
timestamp 18001
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 18001
transform -1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_50
timestamp 18001
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 18001
transform -1 0 28152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_51
timestamp 18001
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 18001
transform -1 0 28152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_52
timestamp 18001
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 18001
transform -1 0 28152 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_53
timestamp 18001
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 18001
transform -1 0 28152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_54
timestamp 18001
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 18001
transform -1 0 28152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_55
timestamp 18001
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 18001
transform -1 0 28152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_56
timestamp 18001
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 18001
transform -1 0 28152 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_57
timestamp 18001
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 18001
transform -1 0 28152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_58
timestamp 18001
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 18001
transform -1 0 28152 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_59
timestamp 18001
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 18001
transform -1 0 28152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_60
timestamp 18001
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 18001
transform -1 0 28152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_61
timestamp 18001
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 18001
transform -1 0 28152 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_62
timestamp 18001
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 18001
transform -1 0 28152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_63
timestamp 18001
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 18001
transform -1 0 28152 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_64
timestamp 18001
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 18001
transform -1 0 28152 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_65
timestamp 18001
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 18001
transform -1 0 28152 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_66
timestamp 18001
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 18001
transform -1 0 28152 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_67
timestamp 18001
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 18001
transform -1 0 28152 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_68
timestamp 18001
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 18001
transform -1 0 28152 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_69
timestamp 18001
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 18001
transform -1 0 28152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_70
timestamp 18001
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 18001
transform -1 0 28152 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_71
timestamp 18001
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 18001
transform -1 0 28152 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_72
timestamp 18001
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 18001
transform -1 0 28152 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_73
timestamp 18001
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 18001
transform -1 0 28152 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_74
timestamp 18001
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 18001
transform -1 0 28152 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_75
timestamp 18001
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 18001
transform -1 0 28152 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_76
timestamp 18001
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 18001
transform -1 0 28152 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_77
timestamp 18001
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 18001
transform -1 0 28152 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_78
timestamp 18001
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 18001
transform -1 0 28152 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_79
timestamp 18001
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 18001
transform -1 0 28152 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_80
timestamp 18001
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 18001
transform -1 0 28152 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_81
timestamp 18001
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 18001
transform -1 0 28152 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_82
timestamp 18001
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 18001
transform -1 0 28152 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_83
timestamp 18001
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 18001
transform -1 0 28152 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_84
timestamp 18001
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 18001
transform -1 0 28152 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_85
timestamp 18001
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 18001
transform -1 0 28152 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_86
timestamp 18001
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 18001
transform -1 0 28152 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_87
timestamp 18001
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 18001
transform -1 0 28152 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_88
timestamp 18001
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 18001
transform -1 0 28152 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_89
timestamp 18001
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 18001
transform -1 0 28152 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_90
timestamp 18001
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 18001
transform -1 0 28152 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_91
timestamp 18001
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 18001
transform -1 0 28152 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_92
timestamp 18001
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 18001
transform -1 0 28152 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_93
timestamp 18001
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 18001
transform -1 0 28152 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_94
timestamp 18001
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 18001
transform -1 0 28152 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_95
timestamp 18001
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 18001
transform -1 0 28152 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_96
timestamp 18001
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 18001
transform -1 0 28152 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_97
timestamp 18001
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 18001
transform -1 0 28152 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_98
timestamp 18001
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_99
timestamp 18001
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_100
timestamp 18001
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_101
timestamp 18001
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_102
timestamp 18001
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_103
timestamp 18001
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_104
timestamp 18001
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_105
timestamp 18001
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_106
timestamp 18001
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_107
timestamp 18001
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_108
timestamp 18001
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_109
timestamp 18001
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_110
timestamp 18001
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_111
timestamp 18001
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_112
timestamp 18001
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_113
timestamp 18001
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_114
timestamp 18001
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_115
timestamp 18001
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_116
timestamp 18001
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_117
timestamp 18001
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_118
timestamp 18001
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_119
timestamp 18001
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_120
timestamp 18001
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_121
timestamp 18001
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_122
timestamp 18001
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_123
timestamp 18001
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_124
timestamp 18001
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_125
timestamp 18001
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_126
timestamp 18001
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_127
timestamp 18001
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_128
timestamp 18001
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_129
timestamp 18001
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_130
timestamp 18001
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_131
timestamp 18001
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_132
timestamp 18001
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_133
timestamp 18001
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_134
timestamp 18001
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_135
timestamp 18001
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_136
timestamp 18001
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_137
timestamp 18001
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_138
timestamp 18001
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_139
timestamp 18001
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_140
timestamp 18001
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_141
timestamp 18001
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_142
timestamp 18001
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_143
timestamp 18001
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_144
timestamp 18001
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_145
timestamp 18001
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_146
timestamp 18001
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_147
timestamp 18001
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_148
timestamp 18001
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_149
timestamp 18001
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_150
timestamp 18001
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_151
timestamp 18001
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_152
timestamp 18001
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_153
timestamp 18001
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_154
timestamp 18001
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_155
timestamp 18001
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_156
timestamp 18001
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_157
timestamp 18001
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_158
timestamp 18001
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_159
timestamp 18001
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_160
timestamp 18001
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_161
timestamp 18001
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_162
timestamp 18001
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_163
timestamp 18001
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_164
timestamp 18001
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_165
timestamp 18001
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_166
timestamp 18001
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_167
timestamp 18001
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_168
timestamp 18001
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_169
timestamp 18001
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_170
timestamp 18001
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_171
timestamp 18001
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_172
timestamp 18001
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_173
timestamp 18001
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_174
timestamp 18001
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_175
timestamp 18001
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_176
timestamp 18001
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_177
timestamp 18001
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_178
timestamp 18001
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_179
timestamp 18001
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_180
timestamp 18001
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_181
timestamp 18001
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_182
timestamp 18001
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_183
timestamp 18001
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_184
timestamp 18001
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_185
timestamp 18001
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_186
timestamp 18001
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_187
timestamp 18001
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_188
timestamp 18001
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_189
timestamp 18001
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_190
timestamp 18001
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_191
timestamp 18001
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_192
timestamp 18001
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_193
timestamp 18001
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_194
timestamp 18001
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_195
timestamp 18001
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_196
timestamp 18001
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_197
timestamp 18001
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_198
timestamp 18001
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_199
timestamp 18001
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_200
timestamp 18001
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_201
timestamp 18001
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_202
timestamp 18001
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_203
timestamp 18001
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_204
timestamp 18001
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_205
timestamp 18001
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_206
timestamp 18001
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_207
timestamp 18001
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_208
timestamp 18001
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_209
timestamp 18001
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_210
timestamp 18001
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_211
timestamp 18001
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_212
timestamp 18001
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_213
timestamp 18001
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_214
timestamp 18001
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_215
timestamp 18001
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_216
timestamp 18001
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_217
timestamp 18001
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_218
timestamp 18001
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_219
timestamp 18001
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_220
timestamp 18001
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_221
timestamp 18001
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_222
timestamp 18001
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_223
timestamp 18001
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_224
timestamp 18001
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_225
timestamp 18001
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_226
timestamp 18001
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_227
timestamp 18001
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_228
timestamp 18001
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_229
timestamp 18001
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_230
timestamp 18001
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_231
timestamp 18001
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_232
timestamp 18001
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_233
timestamp 18001
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_234
timestamp 18001
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_235
timestamp 18001
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_236
timestamp 18001
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_237
timestamp 18001
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_238
timestamp 18001
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_239
timestamp 18001
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_240
timestamp 18001
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_241
timestamp 18001
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_242
timestamp 18001
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_243
timestamp 18001
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_244
timestamp 18001
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_245
timestamp 18001
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_246
timestamp 18001
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_247
timestamp 18001
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_248
timestamp 18001
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_249
timestamp 18001
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_250
timestamp 18001
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_251
timestamp 18001
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_252
timestamp 18001
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_253
timestamp 18001
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_254
timestamp 18001
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_255
timestamp 18001
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_256
timestamp 18001
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_257
timestamp 18001
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_258
timestamp 18001
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_259
timestamp 18001
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_260
timestamp 18001
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_261
timestamp 18001
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_262
timestamp 18001
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_263
timestamp 18001
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_264
timestamp 18001
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_265
timestamp 18001
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_266
timestamp 18001
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_267
timestamp 18001
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_268
timestamp 18001
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_269
timestamp 18001
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_270
timestamp 18001
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_271
timestamp 18001
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_272
timestamp 18001
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_273
timestamp 18001
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_274
timestamp 18001
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_275
timestamp 18001
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_276
timestamp 18001
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_277
timestamp 18001
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_278
timestamp 18001
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_279
timestamp 18001
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_280
timestamp 18001
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_281
timestamp 18001
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_282
timestamp 18001
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_283
timestamp 18001
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_284
timestamp 18001
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_285
timestamp 18001
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_286
timestamp 18001
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_287
timestamp 18001
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_288
timestamp 18001
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_289
timestamp 18001
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_290
timestamp 18001
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_291
timestamp 18001
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_292
timestamp 18001
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_293
timestamp 18001
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_294
timestamp 18001
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_295
timestamp 18001
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_296
timestamp 18001
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_297
timestamp 18001
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_298
timestamp 18001
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_299
timestamp 18001
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_300
timestamp 18001
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_301
timestamp 18001
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_302
timestamp 18001
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_303
timestamp 18001
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_304
timestamp 18001
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_305
timestamp 18001
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_306
timestamp 18001
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_307
timestamp 18001
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_308
timestamp 18001
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_309
timestamp 18001
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_310
timestamp 18001
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_311
timestamp 18001
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_312
timestamp 18001
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_313
timestamp 18001
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_314
timestamp 18001
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_315
timestamp 18001
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_316
timestamp 18001
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_317
timestamp 18001
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_318
timestamp 18001
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_319
timestamp 18001
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_320
timestamp 18001
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_321
timestamp 18001
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_322
timestamp 18001
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_323
timestamp 18001
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_324
timestamp 18001
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_325
timestamp 18001
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_326
timestamp 18001
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_327
timestamp 18001
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_328
timestamp 18001
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_329
timestamp 18001
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_330
timestamp 18001
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_331
timestamp 18001
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_332
timestamp 18001
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_333
timestamp 18001
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_334
timestamp 18001
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_335
timestamp 18001
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_336
timestamp 18001
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_337
timestamp 18001
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_338
timestamp 18001
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_339
timestamp 18001
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_340
timestamp 18001
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_341
timestamp 18001
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_342
timestamp 18001
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_343
timestamp 18001
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_344
timestamp 18001
transform 1 0 6256 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_345
timestamp 18001
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_346
timestamp 18001
transform 1 0 11408 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_347
timestamp 18001
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_348
timestamp 18001
transform 1 0 16560 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_349
timestamp 18001
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_350
timestamp 18001
transform 1 0 21712 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_351
timestamp 18001
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_352
timestamp 18001
transform 1 0 26864 0 1 28288
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 28880 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 28880 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 28532 4768 29332 4888 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 28532 21088 29332 21208 0 FreeSans 480 0 0 0 done
port 3 nsew signal output
flabel metal3 s 28532 6128 29332 6248 0 FreeSans 480 0 0 0 enable
port 4 nsew signal input
flabel metal3 s 28532 5448 29332 5568 0 FreeSans 480 0 0 0 nrst
port 5 nsew signal input
flabel metal3 s 28532 21768 29332 21888 0 FreeSans 480 0 0 0 out[0]
port 6 nsew signal output
flabel metal2 s 23202 30676 23258 31476 0 FreeSans 224 90 0 0 out[10]
port 7 nsew signal output
flabel metal2 s 28998 30676 29054 31476 0 FreeSans 224 90 0 0 out[11]
port 8 nsew signal output
flabel metal2 s 12898 30676 12954 31476 0 FreeSans 224 90 0 0 out[12]
port 9 nsew signal output
flabel metal2 s 14186 30676 14242 31476 0 FreeSans 224 90 0 0 out[13]
port 10 nsew signal output
flabel metal2 s 23846 30676 23902 31476 0 FreeSans 224 90 0 0 out[14]
port 11 nsew signal output
flabel metal2 s 16118 30676 16174 31476 0 FreeSans 224 90 0 0 out[15]
port 12 nsew signal output
flabel metal3 s 28532 23808 29332 23928 0 FreeSans 480 0 0 0 out[16]
port 13 nsew signal output
flabel metal2 s 22558 30676 22614 31476 0 FreeSans 224 90 0 0 out[17]
port 14 nsew signal output
flabel metal2 s 16762 30676 16818 31476 0 FreeSans 224 90 0 0 out[18]
port 15 nsew signal output
flabel metal2 s 25134 30676 25190 31476 0 FreeSans 224 90 0 0 out[19]
port 16 nsew signal output
flabel metal3 s 28532 25168 29332 25288 0 FreeSans 480 0 0 0 out[1]
port 17 nsew signal output
flabel metal2 s 20626 30676 20682 31476 0 FreeSans 224 90 0 0 out[20]
port 18 nsew signal output
flabel metal2 s 18050 30676 18106 31476 0 FreeSans 224 90 0 0 out[21]
port 19 nsew signal output
flabel metal2 s 21914 30676 21970 31476 0 FreeSans 224 90 0 0 out[22]
port 20 nsew signal output
flabel metal2 s 27710 30676 27766 31476 0 FreeSans 224 90 0 0 out[23]
port 21 nsew signal output
flabel metal2 s 14830 30676 14886 31476 0 FreeSans 224 90 0 0 out[24]
port 22 nsew signal output
flabel metal2 s 25778 30676 25834 31476 0 FreeSans 224 90 0 0 out[25]
port 23 nsew signal output
flabel metal3 s 28532 26528 29332 26648 0 FreeSans 480 0 0 0 out[26]
port 24 nsew signal output
flabel metal2 s 26422 30676 26478 31476 0 FreeSans 224 90 0 0 out[27]
port 25 nsew signal output
flabel metal2 s 19982 30676 20038 31476 0 FreeSans 224 90 0 0 out[28]
port 26 nsew signal output
flabel metal2 s 19338 30676 19394 31476 0 FreeSans 224 90 0 0 out[29]
port 27 nsew signal output
flabel metal2 s 18694 30676 18750 31476 0 FreeSans 224 90 0 0 out[2]
port 28 nsew signal output
flabel metal3 s 28532 25848 29332 25968 0 FreeSans 480 0 0 0 out[30]
port 29 nsew signal output
flabel metal3 s 28532 24488 29332 24608 0 FreeSans 480 0 0 0 out[31]
port 30 nsew signal output
flabel metal3 s 28532 22448 29332 22568 0 FreeSans 480 0 0 0 out[32]
port 31 nsew signal output
flabel metal3 s 28532 23128 29332 23248 0 FreeSans 480 0 0 0 out[33]
port 32 nsew signal output
flabel metal2 s 28354 30676 28410 31476 0 FreeSans 224 90 0 0 out[3]
port 33 nsew signal output
flabel metal2 s 15474 30676 15530 31476 0 FreeSans 224 90 0 0 out[4]
port 34 nsew signal output
flabel metal2 s 13542 30676 13598 31476 0 FreeSans 224 90 0 0 out[5]
port 35 nsew signal output
flabel metal2 s 21270 30676 21326 31476 0 FreeSans 224 90 0 0 out[6]
port 36 nsew signal output
flabel metal2 s 24490 30676 24546 31476 0 FreeSans 224 90 0 0 out[7]
port 37 nsew signal output
flabel metal2 s 17406 30676 17462 31476 0 FreeSans 224 90 0 0 out[8]
port 38 nsew signal output
flabel metal2 s 27066 30676 27122 31476 0 FreeSans 224 90 0 0 out[9]
port 39 nsew signal output
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 prescaler[0]
port 40 nsew signal input
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 prescaler[10]
port 41 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 prescaler[11]
port 42 nsew signal input
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 prescaler[12]
port 43 nsew signal input
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 prescaler[13]
port 44 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 prescaler[1]
port 45 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 prescaler[2]
port 46 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 prescaler[3]
port 47 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 prescaler[4]
port 48 nsew signal input
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 prescaler[5]
port 49 nsew signal input
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 prescaler[6]
port 50 nsew signal input
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 prescaler[7]
port 51 nsew signal input
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 prescaler[8]
port 52 nsew signal input
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 prescaler[9]
port 53 nsew signal input
flabel metal3 s 28532 13608 29332 13728 0 FreeSans 480 0 0 0 stop
port 54 nsew signal input
rlabel metal1 14628 28288 14628 28288 0 VGND
rlabel metal1 14628 28832 14628 28832 0 VPWR
rlabel metal2 20562 25534 20562 25534 0 _0000_
rlabel metal1 23552 10030 23552 10030 0 _0001_
rlabel metal1 12880 18190 12880 18190 0 _0002_
rlabel metal2 12558 26792 12558 26792 0 _0003_
rlabel metal1 6072 26554 6072 26554 0 _0004_
rlabel metal1 7958 25942 7958 25942 0 _0005_
rlabel metal1 4554 21862 4554 21862 0 _0006_
rlabel metal1 5014 19380 5014 19380 0 _0007_
rlabel metal1 6762 18054 6762 18054 0 _0008_
rlabel metal1 3818 16048 3818 16048 0 _0009_
rlabel metal1 11362 13838 11362 13838 0 _0010_
rlabel metal1 10396 10234 10396 10234 0 _0011_
rlabel metal2 5382 8942 5382 8942 0 _0012_
rlabel metal1 13018 7820 13018 7820 0 _0013_
rlabel metal1 13892 18802 13892 18802 0 _0014_
rlabel metal1 12236 21114 12236 21114 0 _0015_
rlabel metal1 15318 21386 15318 21386 0 _0016_
rlabel metal1 16790 17680 16790 17680 0 _0017_
rlabel metal2 19366 20604 19366 20604 0 _0018_
rlabel metal1 19366 19312 19366 19312 0 _0019_
rlabel metal1 21252 22066 21252 22066 0 _0020_
rlabel metal2 18078 15572 18078 15572 0 _0021_
rlabel metal1 20700 17170 20700 17170 0 _0022_
rlabel metal2 23230 16320 23230 16320 0 _0023_
rlabel metal2 21022 14688 21022 14688 0 _0024_
rlabel metal1 20378 13158 20378 13158 0 _0025_
rlabel metal1 21068 11118 21068 11118 0 _0026_
rlabel metal2 20930 7140 20930 7140 0 _0027_
rlabel metal2 18078 8160 18078 8160 0 _0028_
rlabel metal2 18078 6970 18078 6970 0 _0029_
rlabel metal1 17434 10642 17434 10642 0 _0030_
rlabel metal1 14858 12818 14858 12818 0 _0031_
rlabel metal2 12834 6970 12834 6970 0 _0032_
rlabel metal1 12420 13702 12420 13702 0 _0033_
rlabel metal1 10764 11798 10764 11798 0 _0034_
rlabel metal1 11914 6834 11914 6834 0 _0035_
rlabel metal1 15778 6800 15778 6800 0 _0036_
rlabel metal1 23920 9350 23920 9350 0 _0037_
rlabel metal2 22034 6596 22034 6596 0 _0038_
rlabel metal1 22770 25942 22770 25942 0 _0039_
rlabel metal2 22402 27302 22402 27302 0 _0040_
rlabel metal1 26358 22644 26358 22644 0 _0041_
rlabel metal1 25668 21930 25668 21930 0 _0042_
rlabel metal1 25484 22746 25484 22746 0 _0043_
rlabel metal1 25990 22066 25990 22066 0 _0044_
rlabel metal1 26174 22134 26174 22134 0 _0045_
rlabel metal1 24518 21454 24518 21454 0 _0046_
rlabel metal1 25208 22542 25208 22542 0 _0047_
rlabel metal2 24794 21692 24794 21692 0 _0048_
rlabel metal1 20194 27438 20194 27438 0 _0049_
rlabel metal1 21620 27642 21620 27642 0 _0050_
rlabel metal1 24472 23154 24472 23154 0 _0051_
rlabel metal1 24150 23052 24150 23052 0 _0052_
rlabel metal1 13064 26010 13064 26010 0 _0053_
rlabel metal1 5520 23154 5520 23154 0 _0054_
rlabel metal2 2530 23970 2530 23970 0 _0055_
rlabel metal1 3174 24752 3174 24752 0 _0056_
rlabel metal1 2852 26282 2852 26282 0 _0057_
rlabel metal1 2990 24820 2990 24820 0 _0058_
rlabel metal1 3634 24242 3634 24242 0 _0059_
rlabel metal1 4554 23732 4554 23732 0 _0060_
rlabel metal1 4646 24174 4646 24174 0 _0061_
rlabel metal2 5106 24514 5106 24514 0 _0062_
rlabel metal1 4462 26316 4462 26316 0 _0063_
rlabel metal1 3320 27030 3320 27030 0 _0064_
rlabel metal2 3910 26554 3910 26554 0 _0065_
rlabel metal1 3772 27098 3772 27098 0 _0066_
rlabel metal2 4094 27132 4094 27132 0 _0067_
rlabel metal2 5290 25840 5290 25840 0 _0068_
rlabel via1 5951 23698 5951 23698 0 _0069_
rlabel metal1 5612 23698 5612 23698 0 _0070_
rlabel metal2 6946 22848 6946 22848 0 _0071_
rlabel metal1 4922 27438 4922 27438 0 _0072_
rlabel metal1 5198 26996 5198 26996 0 _0073_
rlabel metal1 7406 26894 7406 26894 0 _0074_
rlabel metal1 5980 26894 5980 26894 0 _0075_
rlabel metal2 5290 27302 5290 27302 0 _0076_
rlabel metal1 5528 27302 5528 27302 0 _0077_
rlabel viali 5565 26962 5565 26962 0 _0078_
rlabel metal1 5934 26384 5934 26384 0 _0079_
rlabel metal1 7038 23052 7038 23052 0 _0080_
rlabel metal1 7452 22746 7452 22746 0 _0081_
rlabel metal1 7636 21522 7636 21522 0 _0082_
rlabel metal2 7866 22950 7866 22950 0 _0083_
rlabel metal1 6394 25874 6394 25874 0 _0084_
rlabel metal2 6486 26860 6486 26860 0 _0085_
rlabel metal2 6854 26010 6854 26010 0 _0086_
rlabel metal1 7958 24786 7958 24786 0 _0087_
rlabel metal1 7636 24174 7636 24174 0 _0088_
rlabel metal2 8418 24582 8418 24582 0 _0089_
rlabel metal2 8142 23120 8142 23120 0 _0090_
rlabel metal1 8602 22610 8602 22610 0 _0091_
rlabel metal1 10718 23154 10718 23154 0 _0092_
rlabel metal2 8878 22814 8878 22814 0 _0093_
rlabel metal1 10212 21998 10212 21998 0 _0094_
rlabel metal1 4646 11696 4646 11696 0 _0095_
rlabel metal1 2208 10438 2208 10438 0 _0096_
rlabel metal2 2346 11424 2346 11424 0 _0097_
rlabel metal1 8188 9894 8188 9894 0 _0098_
rlabel metal1 4370 13940 4370 13940 0 _0099_
rlabel metal2 2254 13056 2254 13056 0 _0100_
rlabel metal1 2346 14382 2346 14382 0 _0101_
rlabel metal2 2254 11900 2254 11900 0 _0102_
rlabel metal1 3128 11662 3128 11662 0 _0103_
rlabel metal1 3082 10608 3082 10608 0 _0104_
rlabel metal2 3542 11492 3542 11492 0 _0105_
rlabel metal1 3496 11866 3496 11866 0 _0106_
rlabel metal1 2714 13940 2714 13940 0 _0107_
rlabel metal1 4094 15470 4094 15470 0 _0108_
rlabel metal2 1978 17408 1978 17408 0 _0109_
rlabel metal2 2438 17510 2438 17510 0 _0110_
rlabel metal2 2714 16014 2714 16014 0 _0111_
rlabel metal2 2898 14620 2898 14620 0 _0112_
rlabel metal1 3174 14484 3174 14484 0 _0113_
rlabel metal1 3128 12274 3128 12274 0 _0114_
rlabel metal1 4094 12138 4094 12138 0 _0115_
rlabel metal1 4554 12138 4554 12138 0 _0116_
rlabel metal1 5474 12240 5474 12240 0 _0117_
rlabel metal1 3450 15028 3450 15028 0 _0118_
rlabel metal1 2944 16218 2944 16218 0 _0119_
rlabel metal1 4922 18394 4922 18394 0 _0120_
rlabel metal2 2070 20162 2070 20162 0 _0121_
rlabel metal1 2392 20366 2392 20366 0 _0122_
rlabel metal2 2622 17986 2622 17986 0 _0123_
rlabel metal1 3128 17850 3128 17850 0 _0124_
rlabel metal1 2944 17578 2944 17578 0 _0125_
rlabel metal2 3542 15810 3542 15810 0 _0126_
rlabel metal2 3910 14586 3910 14586 0 _0127_
rlabel metal1 4002 14348 4002 14348 0 _0128_
rlabel metal2 5566 13328 5566 13328 0 _0129_
rlabel metal1 7590 13226 7590 13226 0 _0130_
rlabel metal1 6348 12818 6348 12818 0 _0131_
rlabel metal2 7130 13124 7130 13124 0 _0132_
rlabel metal2 5290 14722 5290 14722 0 _0133_
rlabel metal1 3128 19414 3128 19414 0 _0134_
rlabel metal1 5474 20910 5474 20910 0 _0135_
rlabel metal1 2070 21930 2070 21930 0 _0136_
rlabel metal1 3082 23052 3082 23052 0 _0137_
rlabel metal1 3542 20468 3542 20468 0 _0138_
rlabel metal2 3174 20060 3174 20060 0 _0139_
rlabel metal2 3450 20128 3450 20128 0 _0140_
rlabel metal1 4002 17170 4002 17170 0 _0141_
rlabel metal1 3496 17170 3496 17170 0 _0142_
rlabel metal1 4968 16082 4968 16082 0 _0143_
rlabel metal2 4646 16558 4646 16558 0 _0144_
rlabel metal1 4922 14994 4922 14994 0 _0145_
rlabel metal1 6118 14416 6118 14416 0 _0146_
rlabel metal1 6900 14450 6900 14450 0 _0147_
rlabel metal2 6854 13498 6854 13498 0 _0148_
rlabel metal1 8234 13328 8234 13328 0 _0149_
rlabel metal2 5474 8772 5474 8772 0 _0150_
rlabel metal1 3956 8466 3956 8466 0 _0151_
rlabel metal1 3726 8500 3726 8500 0 _0152_
rlabel metal2 2990 9146 2990 9146 0 _0153_
rlabel metal1 3818 8602 3818 8602 0 _0154_
rlabel metal2 4370 7684 4370 7684 0 _0155_
rlabel metal1 4508 8942 4508 8942 0 _0156_
rlabel metal1 4738 9588 4738 9588 0 _0157_
rlabel metal2 4002 9996 4002 9996 0 _0158_
rlabel metal1 5106 9520 5106 9520 0 _0159_
rlabel metal1 4830 9418 4830 9418 0 _0160_
rlabel metal2 5658 10166 5658 10166 0 _0161_
rlabel metal2 5566 11084 5566 11084 0 _0162_
rlabel metal1 6670 10778 6670 10778 0 _0163_
rlabel metal1 6946 10540 6946 10540 0 _0164_
rlabel metal1 7360 11730 7360 11730 0 _0165_
rlabel metal1 7360 12138 7360 12138 0 _0166_
rlabel metal1 8280 12818 8280 12818 0 _0167_
rlabel metal1 8234 12954 8234 12954 0 _0168_
rlabel metal1 8188 10574 8188 10574 0 _0169_
rlabel metal2 5474 7310 5474 7310 0 _0170_
rlabel metal1 5934 6800 5934 6800 0 _0171_
rlabel metal2 7498 9792 7498 9792 0 _0172_
rlabel metal1 7268 8466 7268 8466 0 _0173_
rlabel metal2 6946 7038 6946 7038 0 _0174_
rlabel metal1 6762 7446 6762 7446 0 _0175_
rlabel metal1 8418 6290 8418 6290 0 _0176_
rlabel metal2 6302 6528 6302 6528 0 _0177_
rlabel metal2 5934 6698 5934 6698 0 _0178_
rlabel metal1 6716 6290 6716 6290 0 _0179_
rlabel metal2 6486 6562 6486 6562 0 _0180_
rlabel metal1 7130 7854 7130 7854 0 _0181_
rlabel metal2 6946 8364 6946 8364 0 _0182_
rlabel metal2 8418 9622 8418 9622 0 _0183_
rlabel metal1 7912 7854 7912 7854 0 _0184_
rlabel metal1 8510 6800 8510 6800 0 _0185_
rlabel metal2 8418 6494 8418 6494 0 _0186_
rlabel metal1 7590 8500 7590 8500 0 _0187_
rlabel metal2 7958 9214 7958 9214 0 _0188_
rlabel metal1 8280 10234 8280 10234 0 _0189_
rlabel metal1 8188 9146 8188 9146 0 _0190_
rlabel metal2 9154 7072 9154 7072 0 _0191_
rlabel metal2 8602 7412 8602 7412 0 _0192_
rlabel via1 9162 9962 9162 9962 0 _0193_
rlabel metal2 8050 12767 8050 12767 0 _0194_
rlabel metal1 8878 12954 8878 12954 0 _0195_
rlabel metal1 8694 13770 8694 13770 0 _0196_
rlabel metal2 8694 14246 8694 14246 0 _0197_
rlabel metal1 10212 14994 10212 14994 0 _0198_
rlabel metal2 7314 14994 7314 14994 0 _0199_
rlabel metal2 4830 16252 4830 16252 0 _0200_
rlabel metal1 4462 19856 4462 19856 0 _0201_
rlabel metal2 4002 21692 4002 21692 0 _0202_
rlabel metal1 3220 23086 3220 23086 0 _0203_
rlabel metal2 3818 22814 3818 22814 0 _0204_
rlabel metal1 3910 22610 3910 22610 0 _0205_
rlabel metal2 4738 20638 4738 20638 0 _0206_
rlabel metal2 6026 19516 6026 19516 0 _0207_
rlabel metal1 5428 19346 5428 19346 0 _0208_
rlabel metal1 5704 16082 5704 16082 0 _0209_
rlabel metal1 6072 14994 6072 14994 0 _0210_
rlabel metal1 7544 16558 7544 16558 0 _0211_
rlabel metal2 8142 16048 8142 16048 0 _0212_
rlabel metal1 9108 15130 9108 15130 0 _0213_
rlabel metal2 9890 15198 9890 15198 0 _0214_
rlabel metal1 6164 19142 6164 19142 0 _0215_
rlabel metal1 4876 21522 4876 21522 0 _0216_
rlabel metal2 5290 21760 5290 21760 0 _0217_
rlabel metal1 5198 21454 5198 21454 0 _0218_
rlabel metal1 5980 21454 5980 21454 0 _0219_
rlabel metal2 6578 20094 6578 20094 0 _0220_
rlabel metal1 6624 18326 6624 18326 0 _0221_
rlabel metal1 7544 18190 7544 18190 0 _0222_
rlabel metal1 8050 17306 8050 17306 0 _0223_
rlabel metal2 7222 15470 7222 15470 0 _0224_
rlabel metal2 9338 15674 9338 15674 0 _0225_
rlabel metal2 10258 16796 10258 16796 0 _0226_
rlabel metal2 6946 20876 6946 20876 0 _0227_
rlabel metal1 6532 20434 6532 20434 0 _0228_
rlabel metal1 7038 20366 7038 20366 0 _0229_
rlabel metal1 8280 20434 8280 20434 0 _0230_
rlabel metal2 8786 19210 8786 19210 0 _0231_
rlabel metal2 8694 18598 8694 18598 0 _0232_
rlabel metal1 9614 18258 9614 18258 0 _0233_
rlabel metal2 9246 18428 9246 18428 0 _0234_
rlabel metal1 9890 18292 9890 18292 0 _0235_
rlabel metal1 8234 19482 8234 19482 0 _0236_
rlabel metal2 8602 20366 8602 20366 0 _0237_
rlabel metal1 9430 18292 9430 18292 0 _0238_
rlabel metal1 9476 17646 9476 17646 0 _0239_
rlabel metal1 7544 16218 7544 16218 0 _0240_
rlabel metal1 8878 17068 8878 17068 0 _0241_
rlabel metal2 9614 19924 9614 19924 0 _0242_
rlabel metal2 8234 19142 8234 19142 0 _0243_
rlabel metal1 8694 16694 8694 16694 0 _0244_
rlabel metal1 9384 21998 9384 21998 0 _0245_
rlabel metal1 9706 22066 9706 22066 0 _0246_
rlabel metal1 10258 24174 10258 24174 0 _0247_
rlabel metal1 7222 27506 7222 27506 0 _0248_
rlabel metal2 7406 27132 7406 27132 0 _0249_
rlabel metal1 8234 27030 8234 27030 0 _0250_
rlabel metal1 8050 26928 8050 26928 0 _0251_
rlabel metal2 8234 26350 8234 26350 0 _0252_
rlabel metal1 9062 26282 9062 26282 0 _0253_
rlabel metal1 8694 25840 8694 25840 0 _0254_
rlabel metal2 8694 25228 8694 25228 0 _0255_
rlabel metal2 9338 24140 9338 24140 0 _0256_
rlabel metal2 9430 24378 9430 24378 0 _0257_
rlabel metal1 11040 23086 11040 23086 0 _0258_
rlabel metal1 11638 27438 11638 27438 0 _0259_
rlabel metal1 11822 27404 11822 27404 0 _0260_
rlabel metal1 11914 27472 11914 27472 0 _0261_
rlabel metal2 12466 26418 12466 26418 0 _0262_
rlabel metal2 11270 26690 11270 26690 0 _0263_
rlabel metal1 11132 27098 11132 27098 0 _0264_
rlabel metal1 12742 23120 12742 23120 0 _0265_
rlabel metal1 10672 27642 10672 27642 0 _0266_
rlabel metal2 10258 27370 10258 27370 0 _0267_
rlabel metal1 10534 26962 10534 26962 0 _0268_
rlabel metal2 10902 25738 10902 25738 0 _0269_
rlabel metal2 10718 26010 10718 26010 0 _0270_
rlabel metal1 15134 24718 15134 24718 0 _0271_
rlabel metal2 9338 26826 9338 26826 0 _0272_
rlabel metal1 15594 24854 15594 24854 0 _0273_
rlabel metal1 9752 25262 9752 25262 0 _0274_
rlabel metal1 10028 24854 10028 24854 0 _0275_
rlabel metal1 10488 24582 10488 24582 0 _0276_
rlabel metal2 10534 23290 10534 23290 0 _0277_
rlabel metal2 12006 23732 12006 23732 0 _0278_
rlabel metal1 9660 24106 9660 24106 0 _0279_
rlabel metal1 10718 24276 10718 24276 0 _0280_
rlabel metal1 10764 24786 10764 24786 0 _0281_
rlabel metal1 11638 24582 11638 24582 0 _0282_
rlabel metal1 13386 26384 13386 26384 0 _0283_
rlabel metal1 13064 26282 13064 26282 0 _0284_
rlabel metal2 13110 26554 13110 26554 0 _0285_
rlabel metal2 12650 26146 12650 26146 0 _0286_
rlabel metal2 12098 24922 12098 24922 0 _0287_
rlabel metal1 12696 24310 12696 24310 0 _0288_
rlabel metal2 12650 22780 12650 22780 0 _0289_
rlabel metal1 12880 22950 12880 22950 0 _0290_
rlabel metal2 13846 16626 13846 16626 0 _0291_
rlabel metal1 14306 19890 14306 19890 0 _0292_
rlabel metal2 14122 17136 14122 17136 0 _0293_
rlabel metal2 13294 20230 13294 20230 0 _0294_
rlabel metal1 13524 20502 13524 20502 0 _0295_
rlabel metal1 13984 21386 13984 21386 0 _0296_
rlabel metal2 14030 20706 14030 20706 0 _0297_
rlabel metal1 12466 22032 12466 22032 0 _0298_
rlabel metal1 11960 16082 11960 16082 0 _0299_
rlabel metal1 14444 21930 14444 21930 0 _0300_
rlabel metal2 14306 21794 14306 21794 0 _0301_
rlabel metal2 13018 24378 13018 24378 0 _0302_
rlabel metal1 14858 14926 14858 14926 0 _0303_
rlabel via1 14682 21930 14682 21930 0 _0304_
rlabel metal1 15824 21454 15824 21454 0 _0305_
rlabel metal1 17158 21488 17158 21488 0 _0306_
rlabel metal1 17802 20332 17802 20332 0 _0307_
rlabel metal1 15134 24310 15134 24310 0 _0308_
rlabel metal1 16560 24650 16560 24650 0 _0309_
rlabel metal1 16698 24752 16698 24752 0 _0310_
rlabel metal1 16468 25466 16468 25466 0 _0311_
rlabel metal1 17342 24752 17342 24752 0 _0312_
rlabel metal1 15870 17272 15870 17272 0 _0313_
rlabel metal2 17894 24106 17894 24106 0 _0314_
rlabel metal2 17158 24412 17158 24412 0 _0315_
rlabel metal1 18170 23834 18170 23834 0 _0316_
rlabel metal1 15318 24140 15318 24140 0 _0317_
rlabel metal2 18446 16320 18446 16320 0 _0318_
rlabel metal2 17526 23902 17526 23902 0 _0319_
rlabel metal1 18216 21522 18216 21522 0 _0320_
rlabel metal1 18170 22644 18170 22644 0 _0321_
rlabel metal1 18354 22576 18354 22576 0 _0322_
rlabel metal2 18170 18802 18170 18802 0 _0323_
rlabel metal1 19412 22474 19412 22474 0 _0324_
rlabel metal2 19366 22678 19366 22678 0 _0325_
rlabel metal1 21666 20400 21666 20400 0 _0326_
rlabel metal1 20194 22576 20194 22576 0 _0327_
rlabel metal1 18676 23290 18676 23290 0 _0328_
rlabel metal2 17250 24140 17250 24140 0 _0329_
rlabel metal1 17112 20978 17112 20978 0 _0330_
rlabel metal2 17250 21250 17250 21250 0 _0331_
rlabel metal1 14444 21590 14444 21590 0 _0332_
rlabel metal1 14306 20400 14306 20400 0 _0333_
rlabel metal1 13892 20434 13892 20434 0 _0334_
rlabel metal1 18262 17646 18262 17646 0 _0335_
rlabel metal2 15502 20383 15502 20383 0 _0336_
rlabel metal1 20562 22610 20562 22610 0 _0337_
rlabel metal1 19826 22678 19826 22678 0 _0338_
rlabel metal1 18538 21522 18538 21522 0 _0339_
rlabel metal2 17986 21964 17986 21964 0 _0340_
rlabel metal2 10074 17952 10074 17952 0 _0341_
rlabel metal1 9660 18122 9660 18122 0 _0342_
rlabel metal2 17434 16558 17434 16558 0 _0343_
rlabel metal2 17250 15130 17250 15130 0 _0344_
rlabel metal1 20010 16490 20010 16490 0 _0345_
rlabel via1 20928 16626 20928 16626 0 _0346_
rlabel metal1 20378 16082 20378 16082 0 _0347_
rlabel metal2 20286 15708 20286 15708 0 _0348_
rlabel metal2 9706 15674 9706 15674 0 _0349_
rlabel metal1 16100 16558 16100 16558 0 _0350_
rlabel metal2 16054 16966 16054 16966 0 _0351_
rlabel metal1 21114 14824 21114 14824 0 _0352_
rlabel metal1 21206 14994 21206 14994 0 _0353_
rlabel metal2 20930 14110 20930 14110 0 _0354_
rlabel metal2 20654 14722 20654 14722 0 _0355_
rlabel metal1 19872 14450 19872 14450 0 _0356_
rlabel metal2 8970 13498 8970 13498 0 _0357_
rlabel metal1 18308 12818 18308 12818 0 _0358_
rlabel metal1 18078 12750 18078 12750 0 _0359_
rlabel metal2 19090 11900 19090 11900 0 _0360_
rlabel metal2 18722 11424 18722 11424 0 _0361_
rlabel metal1 18124 12206 18124 12206 0 _0362_
rlabel metal1 18078 13940 18078 13940 0 _0363_
rlabel metal1 20056 11322 20056 11322 0 _0364_
rlabel metal1 18446 14552 18446 14552 0 _0365_
rlabel metal1 9384 6970 9384 6970 0 _0366_
rlabel metal1 15134 7276 15134 7276 0 _0367_
rlabel metal1 16054 9622 16054 9622 0 _0368_
rlabel metal1 8924 7378 8924 7378 0 _0369_
rlabel metal2 16790 9911 16790 9911 0 _0370_
rlabel metal1 15778 11050 15778 11050 0 _0371_
rlabel metal1 8372 9554 8372 9554 0 _0372_
rlabel metal2 14490 9860 14490 9860 0 _0373_
rlabel metal1 14766 14348 14766 14348 0 _0374_
rlabel metal1 15962 10676 15962 10676 0 _0375_
rlabel metal1 8694 10676 8694 10676 0 _0376_
rlabel metal2 11362 10812 11362 10812 0 _0377_
rlabel metal1 14858 9894 14858 9894 0 _0378_
rlabel metal1 12190 8466 12190 8466 0 _0379_
rlabel metal1 13202 7922 13202 7922 0 _0380_
rlabel metal2 11914 9622 11914 9622 0 _0381_
rlabel metal1 12926 9894 12926 9894 0 _0382_
rlabel metal2 10810 11220 10810 11220 0 _0383_
rlabel metal1 11730 10778 11730 10778 0 _0384_
rlabel metal1 11914 10574 11914 10574 0 _0385_
rlabel metal1 11730 10574 11730 10574 0 _0386_
rlabel metal1 13478 10064 13478 10064 0 _0387_
rlabel metal2 13938 10370 13938 10370 0 _0388_
rlabel metal1 18170 10064 18170 10064 0 _0389_
rlabel metal2 9338 10438 9338 10438 0 _0390_
rlabel metal1 15824 7310 15824 7310 0 _0391_
rlabel metal2 20470 7616 20470 7616 0 _0392_
rlabel metal1 18952 9690 18952 9690 0 _0393_
rlabel metal1 18446 8976 18446 8976 0 _0394_
rlabel metal2 9338 8262 9338 8262 0 _0395_
rlabel metal1 16928 12682 16928 12682 0 _0396_
rlabel metal1 18308 8602 18308 8602 0 _0397_
rlabel metal1 18124 14450 18124 14450 0 _0398_
rlabel metal1 18584 10234 18584 10234 0 _0399_
rlabel metal1 18630 9146 18630 9146 0 _0400_
rlabel metal1 18722 10778 18722 10778 0 _0401_
rlabel metal1 19412 11866 19412 11866 0 _0402_
rlabel metal1 20562 16660 20562 16660 0 _0403_
rlabel metal2 20010 15946 20010 15946 0 _0404_
rlabel metal2 20838 15300 20838 15300 0 _0405_
rlabel metal2 19826 14858 19826 14858 0 _0406_
rlabel metal1 18998 21556 18998 21556 0 _0407_
rlabel metal2 18078 17476 18078 17476 0 _0408_
rlabel metal1 20286 20944 20286 20944 0 _0409_
rlabel metal2 21022 17714 21022 17714 0 _0410_
rlabel metal1 24012 11050 24012 11050 0 _0411_
rlabel metal2 13294 7905 13294 7905 0 _0412_
rlabel metal2 12742 8500 12742 8500 0 _0413_
rlabel metal1 14214 9146 14214 9146 0 _0414_
rlabel metal1 16146 9690 16146 9690 0 _0415_
rlabel metal1 17664 10234 17664 10234 0 _0416_
rlabel metal2 18630 17510 18630 17510 0 _0417_
rlabel metal1 19642 20910 19642 20910 0 _0418_
rlabel metal2 17802 14314 17802 14314 0 _0419_
rlabel metal1 9292 10030 9292 10030 0 _0420_
rlabel metal2 9982 10608 9982 10608 0 _0421_
rlabel metal1 18768 12886 18768 12886 0 _0422_
rlabel metal2 22126 12954 22126 12954 0 _0423_
rlabel metal1 23230 12716 23230 12716 0 _0424_
rlabel metal1 14214 13464 14214 13464 0 _0425_
rlabel metal2 22402 14518 22402 14518 0 _0426_
rlabel viali 23138 11118 23138 11118 0 _0427_
rlabel metal1 23368 10982 23368 10982 0 _0428_
rlabel via1 23154 10710 23154 10710 0 _0429_
rlabel metal2 23322 8670 23322 8670 0 _0430_
rlabel metal2 24242 7820 24242 7820 0 _0431_
rlabel metal1 24012 7310 24012 7310 0 _0432_
rlabel metal1 24518 8432 24518 8432 0 _0433_
rlabel metal1 23552 7854 23552 7854 0 _0434_
rlabel metal2 24058 6698 24058 6698 0 _0435_
rlabel metal1 22770 23222 22770 23222 0 _0436_
rlabel metal1 22356 23290 22356 23290 0 _0437_
rlabel metal2 21482 24412 21482 24412 0 _0438_
rlabel metal1 21758 24378 21758 24378 0 _0439_
rlabel metal1 22678 24786 22678 24786 0 _0440_
rlabel metal1 14858 6732 14858 6732 0 _0441_
rlabel metal1 14346 6290 14346 6290 0 _0442_
rlabel metal1 14950 6800 14950 6800 0 _0443_
rlabel metal2 14582 6562 14582 6562 0 _0444_
rlabel via1 10994 6630 10994 6630 0 _0445_
rlabel metal2 12558 6953 12558 6953 0 _0446_
rlabel metal1 12420 6154 12420 6154 0 _0447_
rlabel metal1 10810 6766 10810 6766 0 _0448_
rlabel metal2 10810 7174 10810 7174 0 _0449_
rlabel metal2 11546 11968 11546 11968 0 _0450_
rlabel metal1 12706 10778 12706 10778 0 _0451_
rlabel metal2 12282 12002 12282 12002 0 _0452_
rlabel metal1 11776 12206 11776 12206 0 _0453_
rlabel metal2 11362 12036 11362 12036 0 _0454_
rlabel metal1 11132 11186 11132 11186 0 _0455_
rlabel metal2 12282 14416 12282 14416 0 _0456_
rlabel metal1 12466 13260 12466 13260 0 _0457_
rlabel metal1 12558 12954 12558 12954 0 _0458_
rlabel metal1 12144 13498 12144 13498 0 _0459_
rlabel metal2 13018 14110 13018 14110 0 _0460_
rlabel metal1 11960 14042 11960 14042 0 _0461_
rlabel metal1 12420 6766 12420 6766 0 _0462_
rlabel metal1 15134 9520 15134 9520 0 _0463_
rlabel metal2 12926 9860 12926 9860 0 _0464_
rlabel metal2 12466 8092 12466 8092 0 _0465_
rlabel metal1 17036 8534 17036 8534 0 _0466_
rlabel metal1 14674 10710 14674 10710 0 _0467_
rlabel metal2 15134 11203 15134 11203 0 _0468_
rlabel metal2 14674 13396 14674 13396 0 _0469_
rlabel metal1 15364 13838 15364 13838 0 _0470_
rlabel metal1 16100 11594 16100 11594 0 _0471_
rlabel metal1 15502 10098 15502 10098 0 _0472_
rlabel metal2 14858 10472 14858 10472 0 _0473_
rlabel metal1 15824 10778 15824 10778 0 _0474_
rlabel metal1 16560 11730 16560 11730 0 _0475_
rlabel metal1 17388 6834 17388 6834 0 _0476_
rlabel metal2 17066 8092 17066 8092 0 _0477_
rlabel metal1 17342 7854 17342 7854 0 _0478_
rlabel metal2 17342 7242 17342 7242 0 _0479_
rlabel metal2 16698 6698 16698 6698 0 _0480_
rlabel metal2 18630 7548 18630 7548 0 _0481_
rlabel metal1 20470 7242 20470 7242 0 _0482_
rlabel metal2 20010 7514 20010 7514 0 _0483_
rlabel metal1 18722 7276 18722 7276 0 _0484_
rlabel metal1 20746 7344 20746 7344 0 _0485_
rlabel metal1 21528 7514 21528 7514 0 _0486_
rlabel metal2 20838 7004 20838 7004 0 _0487_
rlabel metal1 20562 7412 20562 7412 0 _0488_
rlabel metal1 20562 10710 20562 10710 0 _0489_
rlabel metal1 21022 9418 21022 9418 0 _0490_
rlabel metal2 21206 9248 21206 9248 0 _0491_
rlabel metal1 20792 9622 20792 9622 0 _0492_
rlabel metal1 20332 10642 20332 10642 0 _0493_
rlabel metal1 18400 13838 18400 13838 0 _0494_
rlabel metal2 22034 13124 22034 13124 0 _0495_
rlabel metal1 21528 12342 21528 12342 0 _0496_
rlabel metal1 20884 12954 20884 12954 0 _0497_
rlabel metal2 18078 13090 18078 13090 0 _0498_
rlabel metal1 18492 12614 18492 12614 0 _0499_
rlabel metal2 22954 14076 22954 14076 0 _0500_
rlabel metal1 24196 13430 24196 13430 0 _0501_
rlabel metal1 23046 13906 23046 13906 0 _0502_
rlabel metal1 23506 16592 23506 16592 0 _0503_
rlabel metal1 23966 15606 23966 15606 0 _0504_
rlabel metal1 23690 14858 23690 14858 0 _0505_
rlabel metal1 23782 15674 23782 15674 0 _0506_
rlabel metal1 23322 16524 23322 16524 0 _0507_
rlabel metal2 21022 17102 21022 17102 0 _0508_
rlabel metal2 21758 16898 21758 16898 0 _0509_
rlabel metal1 23184 17238 23184 17238 0 _0510_
rlabel metal2 20930 17476 20930 17476 0 _0511_
rlabel metal1 21528 17646 21528 17646 0 _0512_
rlabel metal1 17986 14960 17986 14960 0 _0513_
rlabel metal1 17204 15130 17204 15130 0 _0514_
rlabel metal1 16974 15538 16974 15538 0 _0515_
rlabel metal1 21298 20400 21298 20400 0 _0516_
rlabel metal2 20838 19550 20838 19550 0 _0517_
rlabel metal2 22310 19482 22310 19482 0 _0518_
rlabel metal2 21206 20230 21206 20230 0 _0519_
rlabel metal1 21298 19890 21298 19890 0 _0520_
rlabel metal2 21574 20638 21574 20638 0 _0521_
rlabel metal1 17101 21930 17101 21930 0 _0522_
rlabel metal1 19964 19482 19964 19482 0 _0523_
rlabel metal1 19274 19210 19274 19210 0 _0524_
rlabel metal1 18630 18700 18630 18700 0 _0525_
rlabel metal2 18722 18190 18722 18190 0 _0526_
rlabel metal1 18630 20570 18630 20570 0 _0527_
rlabel metal2 20010 21148 20010 21148 0 _0528_
rlabel metal1 18538 20944 18538 20944 0 _0529_
rlabel metal1 18262 20876 18262 20876 0 _0530_
rlabel metal1 18423 18666 18423 18666 0 _0531_
rlabel metal2 16974 21216 16974 21216 0 _0532_
rlabel metal1 17204 20502 17204 20502 0 _0533_
rlabel metal2 17526 18972 17526 18972 0 _0534_
rlabel metal1 16376 18190 16376 18190 0 _0535_
rlabel metal1 16054 17612 16054 17612 0 _0536_
rlabel metal1 14904 20570 14904 20570 0 _0537_
rlabel metal1 14628 20978 14628 20978 0 _0538_
rlabel metal2 14582 21386 14582 21386 0 _0539_
rlabel metal1 14858 21012 14858 21012 0 _0540_
rlabel metal1 15502 20978 15502 20978 0 _0541_
rlabel metal1 14582 20774 14582 20774 0 _0542_
rlabel metal1 11224 20570 11224 20570 0 _0543_
rlabel metal1 12466 18768 12466 18768 0 _0544_
rlabel metal2 12466 20230 12466 20230 0 _0545_
rlabel metal2 11546 20740 11546 20740 0 _0546_
rlabel metal1 15042 18326 15042 18326 0 _0547_
rlabel metal1 14628 17782 14628 17782 0 _0548_
rlabel metal1 14904 17714 14904 17714 0 _0549_
rlabel metal2 12282 17204 12282 17204 0 _0550_
rlabel metal2 12558 18768 12558 18768 0 _0551_
rlabel metal1 12650 18292 12650 18292 0 _0552_
rlabel metal1 12190 16626 12190 16626 0 _0553_
rlabel metal1 23000 8602 23000 8602 0 _0554_
rlabel metal1 21574 13872 21574 13872 0 _0555_
rlabel metal1 23092 13498 23092 13498 0 _0556_
rlabel metal1 22954 11866 22954 11866 0 _0557_
rlabel metal1 21390 13294 21390 13294 0 _0558_
rlabel metal1 15778 14042 15778 14042 0 _0559_
rlabel metal1 15329 7446 15329 7446 0 _0560_
rlabel metal1 15640 7514 15640 7514 0 _0561_
rlabel metal2 15226 8092 15226 8092 0 _0562_
rlabel via3 16675 15300 16675 15300 0 _0563_
rlabel metal1 19734 17170 19734 17170 0 _0564_
rlabel metal1 21436 16762 21436 16762 0 _0565_
rlabel metal2 19366 17340 19366 17340 0 _0566_
rlabel metal1 17342 16014 17342 16014 0 _0567_
rlabel metal1 14996 16082 14996 16082 0 _0568_
rlabel metal1 14536 15946 14536 15946 0 _0569_
rlabel metal2 15134 14824 15134 14824 0 _0570_
rlabel metal1 16054 16082 16054 16082 0 _0571_
rlabel metal2 17158 16694 17158 16694 0 _0572_
rlabel metal1 17388 12614 17388 12614 0 _0573_
rlabel metal1 13110 11322 13110 11322 0 _0574_
rlabel metal1 17158 12172 17158 12172 0 _0575_
rlabel metal1 16514 15470 16514 15470 0 _0576_
rlabel metal1 14444 14926 14444 14926 0 _0577_
rlabel via2 14306 15011 14306 15011 0 _0578_
rlabel metal2 14214 11220 14214 11220 0 _0579_
rlabel metal1 14260 15130 14260 15130 0 _0580_
rlabel metal1 14720 16014 14720 16014 0 _0581_
rlabel metal2 14122 13481 14122 13481 0 _0582_
rlabel metal1 14996 15674 14996 15674 0 _0583_
rlabel metal2 13202 16388 13202 16388 0 _0584_
rlabel metal2 12374 15946 12374 15946 0 _0585_
rlabel metal1 13110 16524 13110 16524 0 _0586_
rlabel metal2 12190 16082 12190 16082 0 _0587_
rlabel metal1 14812 15538 14812 15538 0 _0588_
rlabel metal3 17825 13804 17825 13804 0 _0589_
rlabel metal2 17066 14790 17066 14790 0 _0590_
rlabel metal2 17342 16694 17342 16694 0 _0591_
rlabel metal1 17342 14926 17342 14926 0 _0592_
rlabel metal3 15295 13804 15295 13804 0 _0593_
rlabel metal1 15226 14586 15226 14586 0 _0594_
rlabel metal1 16836 15130 16836 15130 0 _0595_
rlabel metal1 16744 15674 16744 15674 0 _0596_
rlabel metal2 26358 25058 26358 25058 0 _0597_
rlabel metal2 22954 26673 22954 26673 0 _0598_
rlabel metal1 26128 25194 26128 25194 0 _0599_
rlabel metal2 26358 25908 26358 25908 0 _0600_
rlabel metal2 26910 24378 26910 24378 0 _0601_
rlabel metal1 18446 27336 18446 27336 0 _0602_
rlabel metal2 26450 24854 26450 24854 0 _0603_
rlabel metal2 25622 26146 25622 26146 0 _0604_
rlabel metal1 18446 26894 18446 26894 0 _0605_
rlabel metal1 19964 27098 19964 27098 0 _0606_
rlabel metal1 25254 26962 25254 26962 0 _0607_
rlabel metal1 19734 27914 19734 27914 0 _0608_
rlabel metal1 18952 27030 18952 27030 0 _0609_
rlabel metal1 20516 26962 20516 26962 0 _0610_
rlabel metal1 17848 27438 17848 27438 0 _0611_
rlabel metal1 22954 26486 22954 26486 0 _0612_
rlabel metal1 24242 27472 24242 27472 0 _0613_
rlabel metal1 18400 27438 18400 27438 0 _0614_
rlabel metal1 26082 27982 26082 27982 0 _0615_
rlabel metal2 23322 26928 23322 26928 0 _0616_
rlabel metal2 25990 27132 25990 27132 0 _0617_
rlabel metal1 20838 27404 20838 27404 0 _0618_
rlabel metal1 20516 28050 20516 28050 0 _0619_
rlabel metal1 25814 26010 25814 26010 0 _0620_
rlabel metal3 20079 13804 20079 13804 0 clk
rlabel metal1 25162 8568 25162 8568 0 clk_divider.count_out\[0\]
rlabel metal1 17204 8602 17204 8602 0 clk_divider.count_out\[10\]
rlabel metal1 17526 7378 17526 7378 0 clk_divider.count_out\[11\]
rlabel metal1 18630 7854 18630 7854 0 clk_divider.count_out\[12\]
rlabel metal2 19458 9248 19458 9248 0 clk_divider.count_out\[13\]
rlabel metal2 21482 10846 21482 10846 0 clk_divider.count_out\[14\]
rlabel metal2 21298 13124 21298 13124 0 clk_divider.count_out\[15\]
rlabel metal2 24794 13668 24794 13668 0 clk_divider.count_out\[16\]
rlabel metal2 21666 15504 21666 15504 0 clk_divider.count_out\[17\]
rlabel metal1 21390 17136 21390 17136 0 clk_divider.count_out\[18\]
rlabel metal1 22264 19142 22264 19142 0 clk_divider.count_out\[19\]
rlabel metal2 24242 9724 24242 9724 0 clk_divider.count_out\[1\]
rlabel metal1 23138 20910 23138 20910 0 clk_divider.count_out\[20\]
rlabel metal1 20700 19346 20700 19346 0 clk_divider.count_out\[21\]
rlabel metal1 16790 21658 16790 21658 0 clk_divider.count_out\[22\]
rlabel metal2 17342 21760 17342 21760 0 clk_divider.count_out\[23\]
rlabel metal1 14996 21998 14996 21998 0 clk_divider.count_out\[24\]
rlabel metal2 12558 21454 12558 21454 0 clk_divider.count_out\[25\]
rlabel metal1 15364 17646 15364 17646 0 clk_divider.count_out\[26\]
rlabel metal1 13064 16966 13064 16966 0 clk_divider.count_out\[27\]
rlabel metal1 25016 8534 25016 8534 0 clk_divider.count_out\[2\]
rlabel metal2 24334 7854 24334 7854 0 clk_divider.count_out\[3\]
rlabel metal2 15870 6324 15870 6324 0 clk_divider.count_out\[4\]
rlabel metal2 12006 7650 12006 7650 0 clk_divider.count_out\[5\]
rlabel metal1 12052 9078 12052 9078 0 clk_divider.count_out\[6\]
rlabel metal1 12696 13906 12696 13906 0 clk_divider.count_out\[7\]
rlabel metal1 13156 7378 13156 7378 0 clk_divider.count_out\[8\]
rlabel metal2 15778 12988 15778 12988 0 clk_divider.count_out\[9\]
rlabel metal1 23552 11322 23552 11322 0 clk_divider.next_count\[0\]
rlabel metal1 16376 11866 16376 11866 0 clk_divider.next_count\[10\]
rlabel metal1 16284 7310 16284 7310 0 clk_divider.next_count\[11\]
rlabel metal1 17250 13294 17250 13294 0 clk_divider.next_count\[12\]
rlabel metal1 19412 6970 19412 6970 0 clk_divider.next_count\[13\]
rlabel metal1 20378 10098 20378 10098 0 clk_divider.next_count\[14\]
rlabel metal1 19596 12138 19596 12138 0 clk_divider.next_count\[15\]
rlabel metal1 23874 14008 23874 14008 0 clk_divider.next_count\[16\]
rlabel metal2 22310 16286 22310 16286 0 clk_divider.next_count\[17\]
rlabel metal1 18906 16966 18906 16966 0 clk_divider.next_count\[18\]
rlabel metal1 17112 15402 17112 15402 0 clk_divider.next_count\[19\]
rlabel metal2 24702 10268 24702 10268 0 clk_divider.next_count\[1\]
rlabel metal2 22126 20638 22126 20638 0 clk_divider.next_count\[20\]
rlabel metal2 19274 18394 19274 18394 0 clk_divider.next_count\[21\]
rlabel metal1 19734 23834 19734 23834 0 clk_divider.next_count\[22\]
rlabel metal2 15962 21250 15962 21250 0 clk_divider.next_count\[23\]
rlabel metal2 13570 23902 13570 23902 0 clk_divider.next_count\[24\]
rlabel metal1 10626 19720 10626 19720 0 clk_divider.next_count\[25\]
rlabel metal2 14398 16728 14398 16728 0 clk_divider.next_count\[26\]
rlabel metal1 13662 17136 13662 17136 0 clk_divider.next_count\[27\]
rlabel metal2 24702 8092 24702 8092 0 clk_divider.next_count\[2\]
rlabel metal1 23131 6970 23131 6970 0 clk_divider.next_count\[3\]
rlabel metal1 14444 7174 14444 7174 0 clk_divider.next_count\[4\]
rlabel metal1 10488 6970 10488 6970 0 clk_divider.next_count\[5\]
rlabel metal1 10810 9010 10810 9010 0 clk_divider.next_count\[6\]
rlabel metal2 11362 14552 11362 14552 0 clk_divider.next_count\[7\]
rlabel metal2 12190 5882 12190 5882 0 clk_divider.next_count\[8\]
rlabel metal2 14398 13464 14398 13464 0 clk_divider.next_count\[9\]
rlabel metal1 19458 17068 19458 17068 0 clk_divider.next_flag
rlabel metal1 26082 21862 26082 21862 0 clk_divider.rollover_flag
rlabel metal1 19228 14790 19228 14790 0 clknet_0_clk
rlabel metal1 15180 5746 15180 5746 0 clknet_2_0__leaf_clk
rlabel metal1 20332 11866 20332 11866 0 clknet_2_1__leaf_clk
rlabel metal1 16790 18292 16790 18292 0 clknet_2_2__leaf_clk
rlabel metal1 22954 18802 22954 18802 0 clknet_2_3__leaf_clk
rlabel metal1 27140 21658 27140 21658 0 counter_to_35.count_out\[0\]
rlabel metal1 26082 20502 26082 20502 0 counter_to_35.count_out\[1\]
rlabel metal2 21942 23290 21942 23290 0 counter_to_35.count_out\[2\]
rlabel metal2 19918 24208 19918 24208 0 counter_to_35.count_out\[3\]
rlabel metal2 23138 24582 23138 24582 0 counter_to_35.count_out\[4\]
rlabel metal1 27002 24242 27002 24242 0 counter_to_35.count_out\[5\]
rlabel metal1 25438 22202 25438 22202 0 counter_to_35.next_count\[0\]
rlabel metal1 25070 21658 25070 21658 0 counter_to_35.next_count\[1\]
rlabel metal1 23046 23290 23046 23290 0 counter_to_35.next_count\[2\]
rlabel metal2 21390 24174 21390 24174 0 counter_to_35.next_count\[3\]
rlabel metal2 22402 24412 22402 24412 0 counter_to_35.next_count\[4\]
rlabel metal1 24104 23290 24104 23290 0 counter_to_35.next_count\[5\]
rlabel metal2 25714 20808 25714 20808 0 counter_to_35.next_flag
rlabel metal2 27646 21233 27646 21233 0 done
rlabel metal2 27830 6239 27830 6239 0 enable
rlabel metal2 27646 6834 27646 6834 0 net1
rlabel metal1 1886 10676 1886 10676 0 net10
rlabel metal1 1702 17748 1702 17748 0 net11
rlabel metal2 1610 17850 1610 17850 0 net12
rlabel metal2 5152 15844 5152 15844 0 net13
rlabel metal1 2576 10642 2576 10642 0 net14
rlabel metal1 1978 23596 1978 23596 0 net15
rlabel metal2 2346 19006 2346 19006 0 net16
rlabel metal1 25990 21998 25990 21998 0 net17
rlabel metal2 27830 20774 27830 20774 0 net18
rlabel metal1 27462 22406 27462 22406 0 net19
rlabel metal1 26496 8466 26496 8466 0 net2
rlabel metal1 23092 27574 23092 27574 0 net20
rlabel metal2 26358 27574 26358 27574 0 net21
rlabel metal1 18814 28186 18814 28186 0 net22
rlabel via2 20010 27557 20010 27557 0 net23
rlabel metal1 24012 27642 24012 27642 0 net24
rlabel metal2 22034 27744 22034 27744 0 net25
rlabel metal1 27462 24174 27462 24174 0 net26
rlabel metal1 22724 28186 22724 28186 0 net27
rlabel metal2 17250 28152 17250 28152 0 net28
rlabel metal1 25346 27098 25346 27098 0 net29
rlabel metal1 14168 6766 14168 6766 0 net3
rlabel metal1 27232 24378 27232 24378 0 net30
rlabel metal1 20930 27642 20930 27642 0 net31
rlabel metal1 18262 28186 18262 28186 0 net32
rlabel metal1 22310 27642 22310 27642 0 net33
rlabel metal1 27232 27438 27232 27438 0 net34
rlabel metal1 17342 27574 17342 27574 0 net35
rlabel metal1 26404 27642 26404 27642 0 net36
rlabel metal1 26450 26010 26450 26010 0 net37
rlabel metal2 26082 27812 26082 27812 0 net38
rlabel metal1 20332 28186 20332 28186 0 net39
rlabel metal1 2208 19822 2208 19822 0 net4
rlabel metal2 20102 28322 20102 28322 0 net40
rlabel metal1 18860 27098 18860 27098 0 net41
rlabel metal1 26312 25806 26312 25806 0 net42
rlabel metal1 27462 24786 27462 24786 0 net43
rlabel metal1 27462 22610 27462 22610 0 net44
rlabel metal2 27002 23494 27002 23494 0 net45
rlabel metal1 25852 27098 25852 27098 0 net46
rlabel metal1 17388 27098 17388 27098 0 net47
rlabel metal2 17802 27982 17802 27982 0 net48
rlabel metal2 21482 28016 21482 28016 0 net49
rlabel metal1 2162 23086 2162 23086 0 net5
rlabel metal1 24656 27574 24656 27574 0 net50
rlabel metal1 18216 27642 18216 27642 0 net51
rlabel metal1 26634 28118 26634 28118 0 net52
rlabel via2 15594 11747 15594 11747 0 net53
rlabel metal2 15318 20230 15318 20230 0 net54
rlabel metal1 19964 7174 19964 7174 0 net55
rlabel metal2 15134 21063 15134 21063 0 net56
rlabel metal2 12466 16303 12466 16303 0 net57
rlabel metal2 20562 7769 20562 7769 0 net58
rlabel metal2 12834 13260 12834 13260 0 net59
rlabel metal2 2162 24344 2162 24344 0 net6
rlabel metal1 14352 20910 14352 20910 0 net60
rlabel metal1 15180 20434 15180 20434 0 net61
rlabel metal1 20654 7956 20654 7956 0 net62
rlabel metal1 18952 12818 18952 12818 0 net63
rlabel metal1 21896 20910 21896 20910 0 net64
rlabel metal1 20194 13328 20194 13328 0 net65
rlabel metal1 19044 27642 19044 27642 0 net66
rlabel metal2 20930 26996 20930 26996 0 net67
rlabel metal2 22034 22848 22034 22848 0 net68
rlabel metal1 20562 26316 20562 26316 0 net69
rlabel metal1 3496 21862 3496 21862 0 net7
rlabel metal1 19090 27404 19090 27404 0 net70
rlabel metal1 24334 21556 24334 21556 0 net71
rlabel metal1 22034 28016 22034 28016 0 net72
rlabel metal2 27094 24650 27094 24650 0 net73
rlabel metal1 26358 21998 26358 21998 0 net74
rlabel metal1 16146 13192 16146 13192 0 net75
rlabel metal1 21574 20910 21574 20910 0 net76
rlabel metal1 21804 6970 21804 6970 0 net77
rlabel metal2 10074 7956 10074 7956 0 net78
rlabel metal1 12926 25840 12926 25840 0 net79
rlabel metal1 6854 2618 6854 2618 0 net8
rlabel metal1 2438 24208 2438 24208 0 net80
rlabel metal2 13018 25908 13018 25908 0 net81
rlabel metal2 2346 22780 2346 22780 0 net82
rlabel metal1 19918 11764 19918 11764 0 net83
rlabel metal1 21850 9928 21850 9928 0 net84
rlabel metal1 24019 18666 24019 18666 0 net85
rlabel metal2 20378 16830 20378 16830 0 net86
rlabel metal2 1886 17748 1886 17748 0 net87
rlabel metal1 23000 6290 23000 6290 0 net88
rlabel metal1 21022 9554 21022 9554 0 net89
rlabel metal1 2070 10574 2070 10574 0 net9
rlabel via1 20654 15045 20654 15045 0 net90
rlabel metal3 22609 14212 22609 14212 0 net91
rlabel metal1 27692 5678 27692 5678 0 nrst
rlabel via2 27738 21845 27738 21845 0 out[0]
rlabel metal1 23460 28730 23460 28730 0 out[10]
rlabel metal1 27922 28050 27922 28050 0 out[11]
rlabel metal1 12972 28730 12972 28730 0 out[12]
rlabel metal2 14398 29767 14398 29767 0 out[13]
rlabel metal1 24242 28730 24242 28730 0 out[14]
rlabel metal1 16468 28730 16468 28730 0 out[15]
rlabel metal2 27738 23953 27738 23953 0 out[16]
rlabel metal1 22862 28730 22862 28730 0 out[17]
rlabel metal2 17526 28798 17526 28798 0 out[18]
rlabel metal1 25438 28730 25438 28730 0 out[19]
rlabel metal2 27738 25177 27738 25177 0 out[1]
rlabel metal1 20884 28730 20884 28730 0 out[20]
rlabel metal1 18308 28730 18308 28730 0 out[21]
rlabel metal2 21942 29760 21942 29760 0 out[22]
rlabel metal2 27738 29182 27738 29182 0 out[23]
rlabel metal1 14950 28730 14950 28730 0 out[24]
rlabel metal1 25990 28730 25990 28730 0 out[25]
rlabel metal2 27738 26673 27738 26673 0 out[26]
rlabel metal1 26818 28730 26818 28730 0 out[27]
rlabel metal1 20378 28662 20378 28662 0 out[28]
rlabel metal1 19642 28730 19642 28730 0 out[29]
rlabel metal1 19136 28662 19136 28662 0 out[2]
rlabel metal1 27646 26486 27646 26486 0 out[30]
rlabel via2 27738 24565 27738 24565 0 out[31]
rlabel via2 27738 22491 27738 22491 0 out[32]
rlabel metal1 27646 23494 27646 23494 0 out[33]
rlabel metal1 27830 27370 27830 27370 0 out[3]
rlabel metal2 15686 29767 15686 29767 0 out[4]
rlabel metal2 13570 29760 13570 29760 0 out[5]
rlabel metal2 21298 29726 21298 29726 0 out[6]
rlabel metal1 24886 28662 24886 28662 0 out[7]
rlabel metal1 17664 28730 17664 28730 0 out[8]
rlabel metal1 27232 28186 27232 28186 0 out[9]
rlabel metal2 8418 1588 8418 1588 0 prescaler[0]
rlabel metal3 751 23868 751 23868 0 prescaler[10]
rlabel metal3 751 23188 751 23188 0 prescaler[11]
rlabel metal3 751 24548 751 24548 0 prescaler[12]
rlabel metal3 1050 22508 1050 22508 0 prescaler[13]
rlabel metal2 5842 1588 5842 1588 0 prescaler[1]
rlabel metal3 751 11628 751 11628 0 prescaler[2]
rlabel metal3 1050 13668 1050 13668 0 prescaler[3]
rlabel metal3 751 15708 751 15708 0 prescaler[4]
rlabel metal3 1096 17748 1096 17748 0 prescaler[5]
rlabel metal3 1050 20468 1050 20468 0 prescaler[6]
rlabel metal2 2898 21913 2898 21913 0 prescaler[7]
rlabel metal3 1004 21148 1004 21148 0 prescaler[8]
rlabel metal3 751 19788 751 19788 0 prescaler[9]
rlabel metal1 27692 13906 27692 13906 0 stop
<< properties >>
string FIXED_BBOX 0 0 29332 31476
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1727274905
<< viali >>
rect 31033 41089 31067 41123
rect 31217 41021 31251 41055
rect 16313 40613 16347 40647
rect 15853 40545 15887 40579
rect 15761 40477 15795 40511
rect 16037 40477 16071 40511
rect 16589 40477 16623 40511
rect 16313 40409 16347 40443
rect 16221 40341 16255 40375
rect 16497 40341 16531 40375
rect 13546 40137 13580 40171
rect 13461 40069 13495 40103
rect 15301 40069 15335 40103
rect 11989 40001 12023 40035
rect 13369 40001 13403 40035
rect 13645 40001 13679 40035
rect 13921 40001 13955 40035
rect 14749 40001 14783 40035
rect 15025 40001 15059 40035
rect 15761 40001 15795 40035
rect 16221 40001 16255 40035
rect 16681 40001 16715 40035
rect 16865 40001 16899 40035
rect 12081 39933 12115 39967
rect 14013 39933 14047 39967
rect 14381 39933 14415 39967
rect 14657 39933 14691 39967
rect 15393 39933 15427 39967
rect 15853 39933 15887 39967
rect 16497 39933 16531 39967
rect 14289 39865 14323 39899
rect 15117 39865 15151 39899
rect 16037 39865 16071 39899
rect 12357 39797 12391 39831
rect 15209 39797 15243 39831
rect 16405 39797 16439 39831
rect 17049 39797 17083 39831
rect 11989 39593 12023 39627
rect 12357 39593 12391 39627
rect 16221 39593 16255 39627
rect 12541 39525 12575 39559
rect 16129 39525 16163 39559
rect 8309 39457 8343 39491
rect 11897 39457 11931 39491
rect 12725 39457 12759 39491
rect 14289 39457 14323 39491
rect 17049 39457 17083 39491
rect 17601 39457 17635 39491
rect 18061 39457 18095 39491
rect 8585 39389 8619 39423
rect 8769 39389 8803 39423
rect 11253 39389 11287 39423
rect 11437 39389 11471 39423
rect 11529 39389 11563 39423
rect 11713 39389 11747 39423
rect 12173 39389 12207 39423
rect 12449 39389 12483 39423
rect 12817 39389 12851 39423
rect 13001 39389 13035 39423
rect 14473 39389 14507 39423
rect 15577 39389 15611 39423
rect 15761 39389 15795 39423
rect 15853 39389 15887 39423
rect 16037 39389 16071 39423
rect 16313 39389 16347 39423
rect 17141 39389 17175 39423
rect 17969 39389 18003 39423
rect 8493 39253 8527 39287
rect 11345 39253 11379 39287
rect 11621 39253 11655 39287
rect 12449 39253 12483 39287
rect 12909 39253 12943 39287
rect 14657 39253 14691 39287
rect 15669 39253 15703 39287
rect 16589 39253 16623 39287
rect 17509 39253 17543 39287
rect 11989 39049 12023 39083
rect 12081 39049 12115 39083
rect 16865 39049 16899 39083
rect 25789 39049 25823 39083
rect 16681 38981 16715 39015
rect 18061 38981 18095 39015
rect 22937 38981 22971 39015
rect 24685 38981 24719 39015
rect 25697 38981 25731 39015
rect 10241 38913 10275 38947
rect 10425 38913 10459 38947
rect 10793 38913 10827 38947
rect 11069 38913 11103 38947
rect 11805 38913 11839 38947
rect 12265 38913 12299 38947
rect 16957 38913 16991 38947
rect 8309 38845 8343 38879
rect 8585 38845 8619 38879
rect 10885 38845 10919 38879
rect 11529 38845 11563 38879
rect 12449 38845 12483 38879
rect 19809 38845 19843 38879
rect 20085 38845 20119 38879
rect 22661 38845 22695 38879
rect 25513 38845 25547 38879
rect 10241 38777 10275 38811
rect 10977 38777 11011 38811
rect 11621 38777 11655 38811
rect 10057 38709 10091 38743
rect 10609 38709 10643 38743
rect 16681 38709 16715 38743
rect 26157 38709 26191 38743
rect 8033 38505 8067 38539
rect 8769 38505 8803 38539
rect 9413 38505 9447 38539
rect 9965 38505 9999 38539
rect 10517 38505 10551 38539
rect 11529 38505 11563 38539
rect 18521 38505 18555 38539
rect 23213 38505 23247 38539
rect 7941 38437 7975 38471
rect 21281 38437 21315 38471
rect 7757 38369 7791 38403
rect 13001 38369 13035 38403
rect 23857 38369 23891 38403
rect 26617 38369 26651 38403
rect 26709 38369 26743 38403
rect 28457 38369 28491 38403
rect 5457 38301 5491 38335
rect 5733 38301 5767 38335
rect 8033 38301 8067 38335
rect 8125 38301 8159 38335
rect 8309 38301 8343 38335
rect 8401 38301 8435 38335
rect 8493 38301 8527 38335
rect 8953 38301 8987 38335
rect 9045 38301 9079 38335
rect 9229 38301 9263 38335
rect 9781 38301 9815 38335
rect 9965 38301 9999 38335
rect 10241 38301 10275 38335
rect 10333 38301 10367 38335
rect 11345 38301 11379 38335
rect 11529 38301 11563 38335
rect 12633 38301 12667 38335
rect 12817 38301 12851 38335
rect 12909 38301 12943 38335
rect 13185 38301 13219 38335
rect 17785 38301 17819 38335
rect 17969 38301 18003 38335
rect 18061 38301 18095 38335
rect 18153 38301 18187 38335
rect 18337 38301 18371 38335
rect 20729 38301 20763 38335
rect 20913 38301 20947 38335
rect 21465 38301 21499 38335
rect 21557 38301 21591 38335
rect 21741 38301 21775 38335
rect 22937 38301 22971 38335
rect 24593 38301 24627 38335
rect 28733 38301 28767 38335
rect 5641 38233 5675 38267
rect 21097 38233 21131 38267
rect 23581 38233 23615 38267
rect 23673 38233 23707 38267
rect 24869 38233 24903 38267
rect 5273 38165 5307 38199
rect 13369 38165 13403 38199
rect 21649 38165 21683 38199
rect 23029 38165 23063 38199
rect 8677 37961 8711 37995
rect 18061 37961 18095 37995
rect 24961 37961 24995 37995
rect 25421 37961 25455 37995
rect 4445 37893 4479 37927
rect 6193 37893 6227 37927
rect 13277 37893 13311 37927
rect 15485 37893 15519 37927
rect 25329 37893 25363 37927
rect 8861 37825 8895 37859
rect 9137 37825 9171 37859
rect 9321 37825 9355 37859
rect 9413 37825 9447 37859
rect 9597 37825 9631 37859
rect 15117 37825 15151 37859
rect 15301 37825 15335 37859
rect 15577 37825 15611 37859
rect 15761 37825 15795 37859
rect 15853 37825 15887 37859
rect 15945 37825 15979 37859
rect 17601 37825 17635 37859
rect 17693 37825 17727 37859
rect 17877 37825 17911 37859
rect 18429 37825 18463 37859
rect 18981 37825 19015 37859
rect 19165 37825 19199 37859
rect 19349 37825 19383 37859
rect 19533 37825 19567 37859
rect 19809 37825 19843 37859
rect 22017 37825 22051 37859
rect 22109 37825 22143 37859
rect 4169 37757 4203 37791
rect 6377 37757 6411 37791
rect 6653 37757 6687 37791
rect 9045 37757 9079 37791
rect 9229 37757 9263 37791
rect 13001 37757 13035 37791
rect 15025 37757 15059 37791
rect 19257 37757 19291 37791
rect 19717 37757 19751 37791
rect 20085 37757 20119 37791
rect 21833 37757 21867 37791
rect 22385 37757 22419 37791
rect 22661 37757 22695 37791
rect 24409 37757 24443 37791
rect 25513 37757 25547 37791
rect 8125 37621 8159 37655
rect 9413 37621 9447 37655
rect 16221 37621 16255 37655
rect 18521 37621 18555 37655
rect 21557 37621 21591 37655
rect 21925 37621 21959 37655
rect 6469 37417 6503 37451
rect 7849 37417 7883 37451
rect 8953 37417 8987 37451
rect 12725 37417 12759 37451
rect 14933 37417 14967 37451
rect 17325 37417 17359 37451
rect 17601 37417 17635 37451
rect 20545 37417 20579 37451
rect 21373 37417 21407 37451
rect 23029 37417 23063 37451
rect 17417 37349 17451 37383
rect 21741 37349 21775 37383
rect 5181 37281 5215 37315
rect 6101 37281 6135 37315
rect 8125 37281 8159 37315
rect 12265 37281 12299 37315
rect 12449 37281 12483 37315
rect 15301 37281 15335 37315
rect 17233 37281 17267 37315
rect 18521 37281 18555 37315
rect 18613 37281 18647 37315
rect 20729 37281 20763 37315
rect 23489 37281 23523 37315
rect 23673 37281 23707 37315
rect 25973 37281 26007 37315
rect 5365 37213 5399 37247
rect 5549 37213 5583 37247
rect 5641 37213 5675 37247
rect 5733 37213 5767 37247
rect 5917 37213 5951 37247
rect 6009 37213 6043 37247
rect 6285 37213 6319 37247
rect 7757 37213 7791 37247
rect 7941 37213 7975 37247
rect 8401 37213 8435 37247
rect 8585 37213 8619 37247
rect 9137 37213 9171 37247
rect 9321 37213 9355 37247
rect 9413 37213 9447 37247
rect 12541 37213 12575 37247
rect 12633 37213 12667 37247
rect 12817 37213 12851 37247
rect 14473 37213 14507 37247
rect 14749 37213 14783 37247
rect 15025 37213 15059 37247
rect 17049 37213 17083 37247
rect 17509 37213 17543 37247
rect 17785 37213 17819 37247
rect 18061 37213 18095 37247
rect 18337 37213 18371 37247
rect 18429 37213 18463 37247
rect 19257 37213 19291 37247
rect 19717 37213 19751 37247
rect 20821 37213 20855 37247
rect 21281 37213 21315 37247
rect 21465 37213 21499 37247
rect 21557 37213 21591 37247
rect 21741 37213 21775 37247
rect 25881 37213 25915 37247
rect 25789 37145 25823 37179
rect 8309 37077 8343 37111
rect 12265 37077 12299 37111
rect 14565 37077 14599 37111
rect 17969 37077 18003 37111
rect 18797 37077 18831 37111
rect 19349 37077 19383 37111
rect 19441 37077 19475 37111
rect 23397 37077 23431 37111
rect 25421 37077 25455 37111
rect 6009 36873 6043 36907
rect 8493 36873 8527 36907
rect 11805 36873 11839 36907
rect 12541 36873 12575 36907
rect 15669 36873 15703 36907
rect 18245 36873 18279 36907
rect 18981 36873 19015 36907
rect 6469 36805 6503 36839
rect 8769 36805 8803 36839
rect 14473 36805 14507 36839
rect 15393 36805 15427 36839
rect 15577 36805 15611 36839
rect 25053 36805 25087 36839
rect 26801 36805 26835 36839
rect 5549 36737 5583 36771
rect 5825 36737 5859 36771
rect 6009 36737 6043 36771
rect 6377 36737 6411 36771
rect 6561 36737 6595 36771
rect 8493 36737 8527 36771
rect 8585 36737 8619 36771
rect 10701 36737 10735 36771
rect 10793 36737 10827 36771
rect 10977 36737 11011 36771
rect 11069 36737 11103 36771
rect 11713 36737 11747 36771
rect 12173 36737 12207 36771
rect 12909 36737 12943 36771
rect 13553 36737 13587 36771
rect 13829 36737 13863 36771
rect 14013 36737 14047 36771
rect 15209 36737 15243 36771
rect 15853 36737 15887 36771
rect 16129 36737 16163 36771
rect 16313 36737 16347 36771
rect 16865 36737 16899 36771
rect 17049 36737 17083 36771
rect 17141 36737 17175 36771
rect 18061 36737 18095 36771
rect 18705 36737 18739 36771
rect 23765 36737 23799 36771
rect 12265 36669 12299 36703
rect 13001 36669 13035 36703
rect 13369 36669 13403 36703
rect 14197 36669 14231 36703
rect 14381 36669 14415 36703
rect 17877 36669 17911 36703
rect 18981 36669 19015 36703
rect 23029 36669 23063 36703
rect 24777 36669 24811 36703
rect 17141 36601 17175 36635
rect 5687 36533 5721 36567
rect 10517 36533 10551 36567
rect 13185 36533 13219 36567
rect 14841 36533 14875 36567
rect 18797 36533 18831 36567
rect 6469 36329 6503 36363
rect 7849 36329 7883 36363
rect 7941 36329 7975 36363
rect 9229 36329 9263 36363
rect 9413 36329 9447 36363
rect 15761 36329 15795 36363
rect 5917 36261 5951 36295
rect 15301 36261 15335 36295
rect 21557 36261 21591 36295
rect 8309 36193 8343 36227
rect 10333 36193 10367 36227
rect 14565 36193 14599 36227
rect 14749 36193 14783 36227
rect 14933 36193 14967 36227
rect 15853 36193 15887 36227
rect 22017 36193 22051 36227
rect 22385 36193 22419 36227
rect 24133 36193 24167 36227
rect 25145 36193 25179 36227
rect 27169 36193 27203 36227
rect 3985 36125 4019 36159
rect 4261 36125 4295 36159
rect 6101 36125 6135 36159
rect 6193 36125 6227 36159
rect 7297 36125 7331 36159
rect 7665 36125 7699 36159
rect 8125 36125 8159 36159
rect 8401 36125 8435 36159
rect 9137 36125 9171 36159
rect 9229 36125 9263 36159
rect 9781 36125 9815 36159
rect 10057 36125 10091 36159
rect 10241 36125 10275 36159
rect 12357 36125 12391 36159
rect 12725 36125 12759 36159
rect 12817 36125 12851 36159
rect 15117 36125 15151 36159
rect 15577 36125 15611 36159
rect 15669 36125 15703 36159
rect 18153 36125 18187 36159
rect 18337 36125 18371 36159
rect 19625 36125 19659 36159
rect 21925 36125 21959 36159
rect 22293 36125 22327 36159
rect 22477 36125 22511 36159
rect 23305 36125 23339 36159
rect 3801 36057 3835 36091
rect 5917 36057 5951 36091
rect 6285 36057 6319 36091
rect 6485 36057 6519 36091
rect 6837 36057 6871 36091
rect 7021 36057 7055 36091
rect 7205 36057 7239 36091
rect 7481 36057 7515 36091
rect 7573 36057 7607 36091
rect 8953 36057 8987 36091
rect 10609 36057 10643 36091
rect 12449 36057 12483 36091
rect 13001 36057 13035 36091
rect 19901 36057 19935 36091
rect 23857 36057 23891 36091
rect 23949 36057 23983 36091
rect 25421 36057 25455 36091
rect 4169 35989 4203 36023
rect 6653 35989 6687 36023
rect 9597 35989 9631 36023
rect 12633 35989 12667 36023
rect 14105 35989 14139 36023
rect 14473 35989 14507 36023
rect 18245 35989 18279 36023
rect 21373 35989 21407 36023
rect 23489 35989 23523 36023
rect 6377 35785 6411 35819
rect 7573 35785 7607 35819
rect 8861 35785 8895 35819
rect 9045 35785 9079 35819
rect 10793 35785 10827 35819
rect 12081 35785 12115 35819
rect 19809 35785 19843 35819
rect 21189 35785 21223 35819
rect 25329 35785 25363 35819
rect 25789 35785 25823 35819
rect 2329 35717 2363 35751
rect 2513 35717 2547 35751
rect 4261 35717 4295 35751
rect 7113 35717 7147 35751
rect 11161 35717 11195 35751
rect 11621 35717 11655 35751
rect 17233 35717 17267 35751
rect 23305 35717 23339 35751
rect 25053 35717 25087 35751
rect 2145 35649 2179 35683
rect 2421 35649 2455 35683
rect 4537 35649 4571 35683
rect 6009 35649 6043 35683
rect 6561 35649 6595 35683
rect 6929 35649 6963 35683
rect 7481 35649 7515 35683
rect 7665 35649 7699 35683
rect 8493 35649 8527 35683
rect 8677 35649 8711 35683
rect 9229 35649 9263 35683
rect 9321 35649 9355 35683
rect 9505 35649 9539 35683
rect 10517 35649 10551 35683
rect 10876 35649 10910 35683
rect 10977 35649 11011 35683
rect 11713 35649 11747 35683
rect 11897 35649 11931 35683
rect 12081 35649 12115 35683
rect 13461 35649 13495 35683
rect 15669 35649 15703 35683
rect 15761 35649 15795 35683
rect 15853 35649 15887 35683
rect 15945 35649 15979 35683
rect 17141 35649 17175 35683
rect 17417 35649 17451 35683
rect 17601 35649 17635 35683
rect 18337 35649 18371 35683
rect 18521 35649 18555 35683
rect 19073 35649 19107 35683
rect 19257 35649 19291 35683
rect 19441 35649 19475 35683
rect 19625 35649 19659 35683
rect 21005 35649 21039 35683
rect 21189 35649 21223 35683
rect 21556 35649 21590 35683
rect 21649 35649 21683 35683
rect 21833 35649 21867 35683
rect 23029 35649 23063 35683
rect 25697 35649 25731 35683
rect 6837 35581 6871 35615
rect 10609 35581 10643 35615
rect 10793 35581 10827 35615
rect 13737 35581 13771 35615
rect 15485 35581 15519 35615
rect 16129 35581 16163 35615
rect 17877 35581 17911 35615
rect 17969 35581 18003 35615
rect 18061 35581 18095 35615
rect 18153 35581 18187 35615
rect 18429 35581 18463 35615
rect 19349 35581 19383 35615
rect 22569 35581 22603 35615
rect 25881 35581 25915 35615
rect 6101 35513 6135 35547
rect 11161 35513 11195 35547
rect 17693 35513 17727 35547
rect 1961 35445 1995 35479
rect 6745 35445 6779 35479
rect 7297 35445 7331 35479
rect 9321 35445 9355 35479
rect 21465 35445 21499 35479
rect 4169 35241 4203 35275
rect 7389 35241 7423 35275
rect 7757 35241 7791 35275
rect 8217 35241 8251 35275
rect 16221 35241 16255 35275
rect 16681 35241 16715 35275
rect 22293 35241 22327 35275
rect 7021 35173 7055 35207
rect 8953 35173 8987 35207
rect 17049 35173 17083 35207
rect 17233 35173 17267 35207
rect 19349 35173 19383 35207
rect 19717 35173 19751 35207
rect 3157 35105 3191 35139
rect 3433 35105 3467 35139
rect 5917 35105 5951 35139
rect 6009 35105 6043 35139
rect 6469 35105 6503 35139
rect 8309 35105 8343 35139
rect 8769 35105 8803 35139
rect 9229 35105 9263 35139
rect 9321 35105 9355 35139
rect 12541 35105 12575 35139
rect 16313 35105 16347 35139
rect 17601 35105 17635 35139
rect 21281 35105 21315 35139
rect 21557 35105 21591 35139
rect 6377 35037 6411 35071
rect 6929 35037 6963 35071
rect 7113 35037 7147 35071
rect 7205 35037 7239 35071
rect 7389 35037 7423 35071
rect 7573 35037 7607 35071
rect 8033 35037 8067 35071
rect 8217 35037 8251 35071
rect 8493 35037 8527 35071
rect 8677 35037 8711 35071
rect 9137 35037 9171 35071
rect 9413 35037 9447 35071
rect 12265 35037 12299 35071
rect 12449 35037 12483 35071
rect 12909 35037 12943 35071
rect 16497 35037 16531 35071
rect 17693 35037 17727 35071
rect 17877 35037 17911 35071
rect 18061 35037 18095 35071
rect 18337 35037 18371 35071
rect 19533 35037 19567 35071
rect 19901 35037 19935 35071
rect 20729 35037 20763 35071
rect 20913 35037 20947 35071
rect 21189 35037 21223 35071
rect 21925 35037 21959 35071
rect 22477 35037 22511 35071
rect 1409 34969 1443 35003
rect 5641 34969 5675 35003
rect 6745 34969 6779 35003
rect 16221 34969 16255 35003
rect 16773 34969 16807 35003
rect 17325 34969 17359 35003
rect 17785 34969 17819 35003
rect 22661 34969 22695 35003
rect 22937 34969 22971 35003
rect 6653 34901 6687 34935
rect 12081 34901 12115 34935
rect 12725 34901 12759 34935
rect 17417 34901 17451 34935
rect 18521 34901 18555 34935
rect 20913 34901 20947 34935
rect 22845 34901 22879 34935
rect 7021 34697 7055 34731
rect 8769 34697 8803 34731
rect 17417 34697 17451 34731
rect 18337 34697 18371 34731
rect 10977 34629 11011 34663
rect 17601 34629 17635 34663
rect 19533 34629 19567 34663
rect 19901 34629 19935 34663
rect 25605 34629 25639 34663
rect 4353 34561 4387 34595
rect 6377 34561 6411 34595
rect 6561 34561 6595 34595
rect 6653 34561 6687 34595
rect 6745 34561 6779 34595
rect 8677 34561 8711 34595
rect 8861 34561 8895 34595
rect 9229 34561 9263 34595
rect 9413 34561 9447 34595
rect 9965 34561 9999 34595
rect 10149 34561 10183 34595
rect 10609 34561 10643 34595
rect 10839 34561 10873 34595
rect 11069 34561 11103 34595
rect 11252 34561 11286 34595
rect 11345 34561 11379 34595
rect 11897 34561 11931 34595
rect 14381 34561 14415 34595
rect 17325 34561 17359 34595
rect 18245 34561 18279 34595
rect 18521 34561 18555 34595
rect 18705 34561 18739 34595
rect 18797 34561 18831 34595
rect 18981 34561 19015 34595
rect 19165 34561 19199 34595
rect 19349 34561 19383 34595
rect 22017 34561 22051 34595
rect 22109 34561 22143 34595
rect 22201 34561 22235 34595
rect 22339 34561 22373 34595
rect 22569 34561 22603 34595
rect 22937 34561 22971 34595
rect 23581 34561 23615 34595
rect 30389 34561 30423 34595
rect 2329 34493 2363 34527
rect 4077 34493 4111 34527
rect 10333 34493 10367 34527
rect 11989 34493 12023 34527
rect 12265 34493 12299 34527
rect 13737 34493 13771 34527
rect 14289 34493 14323 34527
rect 19073 34493 19107 34527
rect 19625 34493 19659 34527
rect 21649 34493 21683 34527
rect 22477 34493 22511 34527
rect 23857 34493 23891 34527
rect 28365 34493 28399 34527
rect 10517 34425 10551 34459
rect 9229 34357 9263 34391
rect 10149 34357 10183 34391
rect 10425 34357 10459 34391
rect 10701 34357 10735 34391
rect 11713 34357 11747 34391
rect 14657 34357 14691 34391
rect 17601 34357 17635 34391
rect 21833 34357 21867 34391
rect 29009 34357 29043 34391
rect 3065 34153 3099 34187
rect 8769 34153 8803 34187
rect 9229 34153 9263 34187
rect 9965 34153 9999 34187
rect 10793 34153 10827 34187
rect 10977 34153 11011 34187
rect 11989 34153 12023 34187
rect 12633 34153 12667 34187
rect 18429 34153 18463 34187
rect 18797 34153 18831 34187
rect 24409 34153 24443 34187
rect 27445 34153 27479 34187
rect 9597 34085 9631 34119
rect 18705 34085 18739 34119
rect 21649 34085 21683 34119
rect 9045 34017 9079 34051
rect 10057 34017 10091 34051
rect 10425 34017 10459 34051
rect 10885 34017 10919 34051
rect 12357 34017 12391 34051
rect 14473 34017 14507 34051
rect 14749 34017 14783 34051
rect 17049 34017 17083 34051
rect 17233 34017 17267 34051
rect 17601 34017 17635 34051
rect 17785 34017 17819 34051
rect 18889 34017 18923 34051
rect 20361 34017 20395 34051
rect 21925 34017 21959 34051
rect 25053 34017 25087 34051
rect 29193 34017 29227 34051
rect 29745 34017 29779 34051
rect 3249 33949 3283 33983
rect 3525 33949 3559 33983
rect 8493 33949 8527 33983
rect 8585 33949 8619 33983
rect 8953 33949 8987 33983
rect 9137 33949 9171 33983
rect 9413 33949 9447 33983
rect 9689 33949 9723 33983
rect 10149 33949 10183 33983
rect 10609 33949 10643 33983
rect 11161 33949 11195 33983
rect 11345 33949 11379 33983
rect 11805 33949 11839 33983
rect 11989 33949 12023 33983
rect 12265 33949 12299 33983
rect 12909 33949 12943 33983
rect 13093 33949 13127 33983
rect 17417 33949 17451 33983
rect 17509 33949 17543 33983
rect 17877 33949 17911 33983
rect 18153 33949 18187 33983
rect 18613 33949 18647 33983
rect 20453 33949 20487 33983
rect 22017 33949 22051 33983
rect 24869 33949 24903 33983
rect 30113 33949 30147 33983
rect 32137 33949 32171 33983
rect 3433 33881 3467 33915
rect 12725 33881 12759 33915
rect 28917 33881 28951 33915
rect 32413 33881 32447 33915
rect 9781 33813 9815 33847
rect 16221 33813 16255 33847
rect 17601 33813 17635 33847
rect 20085 33813 20119 33847
rect 24777 33813 24811 33847
rect 31539 33813 31573 33847
rect 33885 33813 33919 33847
rect 5641 33609 5675 33643
rect 6377 33609 6411 33643
rect 6745 33609 6779 33643
rect 8953 33609 8987 33643
rect 9873 33609 9907 33643
rect 10425 33609 10459 33643
rect 14197 33609 14231 33643
rect 15669 33609 15703 33643
rect 20177 33609 20211 33643
rect 30113 33609 30147 33643
rect 30205 33609 30239 33643
rect 32689 33609 32723 33643
rect 2329 33541 2363 33575
rect 6101 33541 6135 33575
rect 10149 33541 10183 33575
rect 15301 33541 15335 33575
rect 15485 33541 15519 33575
rect 29837 33541 29871 33575
rect 33057 33541 33091 33575
rect 33517 33541 33551 33575
rect 34437 33541 34471 33575
rect 2237 33473 2271 33507
rect 2513 33473 2547 33507
rect 3157 33473 3191 33507
rect 5549 33473 5583 33507
rect 6009 33473 6043 33507
rect 6193 33473 6227 33507
rect 7205 33473 7239 33507
rect 7389 33473 7423 33507
rect 7849 33473 7883 33507
rect 8033 33473 8067 33507
rect 8309 33473 8343 33507
rect 8493 33473 8527 33507
rect 9413 33473 9447 33507
rect 9597 33473 9631 33507
rect 9689 33473 9723 33507
rect 10057 33473 10091 33507
rect 10241 33473 10275 33507
rect 10333 33473 10367 33507
rect 10517 33473 10551 33507
rect 14565 33473 14599 33507
rect 19809 33473 19843 33507
rect 28733 33473 28767 33507
rect 29561 33473 29595 33507
rect 29745 33473 29779 33507
rect 29929 33473 29963 33507
rect 30481 33473 30515 33507
rect 30757 33473 30791 33507
rect 31401 33473 31435 33507
rect 31953 33473 31987 33507
rect 32873 33473 32907 33507
rect 33149 33473 33183 33507
rect 34069 33473 34103 33507
rect 34253 33473 34287 33507
rect 3249 33405 3283 33439
rect 3433 33405 3467 33439
rect 5825 33405 5859 33439
rect 6837 33405 6871 33439
rect 6929 33405 6963 33439
rect 8125 33405 8159 33439
rect 14657 33405 14691 33439
rect 14749 33405 14783 33439
rect 17693 33405 17727 33439
rect 17969 33405 18003 33439
rect 19717 33405 19751 33439
rect 28457 33405 28491 33439
rect 28825 33405 28859 33439
rect 30205 33405 30239 33439
rect 31677 33405 31711 33439
rect 2697 33337 2731 33371
rect 7297 33337 7331 33371
rect 9137 33337 9171 33371
rect 2789 33269 2823 33303
rect 5181 33269 5215 33303
rect 7665 33269 7699 33303
rect 19441 33269 19475 33303
rect 26985 33269 27019 33303
rect 29469 33269 29503 33303
rect 30389 33269 30423 33303
rect 34621 33269 34655 33303
rect 5641 33065 5675 33099
rect 8677 33065 8711 33099
rect 15577 33065 15611 33099
rect 16405 33065 16439 33099
rect 18337 33065 18371 33099
rect 28549 33065 28583 33099
rect 29653 33065 29687 33099
rect 33563 33065 33597 33099
rect 3249 32929 3283 32963
rect 4169 32929 4203 32963
rect 6653 32929 6687 32963
rect 6929 32929 6963 32963
rect 7205 32929 7239 32963
rect 29193 32929 29227 32963
rect 29929 32929 29963 32963
rect 31769 32929 31803 32963
rect 3525 32861 3559 32895
rect 3893 32861 3927 32895
rect 11621 32861 11655 32895
rect 11713 32861 11747 32895
rect 15577 32861 15611 32895
rect 15761 32861 15795 32895
rect 16313 32861 16347 32895
rect 16497 32861 16531 32895
rect 17601 32861 17635 32895
rect 17785 32861 17819 32895
rect 17877 32861 17911 32895
rect 17969 32861 18003 32895
rect 18153 32861 18187 32895
rect 23949 32861 23983 32895
rect 25697 32861 25731 32895
rect 25973 32861 26007 32895
rect 26127 32861 26161 32895
rect 28733 32861 28767 32895
rect 28825 32861 28859 32895
rect 29055 32861 29089 32895
rect 29561 32861 29595 32895
rect 29745 32861 29779 32895
rect 32137 32861 32171 32895
rect 33701 32861 33735 32895
rect 34713 32861 34747 32895
rect 36737 32861 36771 32895
rect 1501 32793 1535 32827
rect 6469 32793 6503 32827
rect 23673 32793 23707 32827
rect 28917 32793 28951 32827
rect 30205 32793 30239 32827
rect 34345 32793 34379 32827
rect 36461 32793 36495 32827
rect 6101 32725 6135 32759
rect 6561 32725 6595 32759
rect 11253 32725 11287 32759
rect 11897 32725 11931 32759
rect 16129 32725 16163 32759
rect 23771 32725 23805 32759
rect 23857 32725 23891 32759
rect 25513 32725 25547 32759
rect 26341 32725 26375 32759
rect 31677 32725 31711 32759
rect 34437 32725 34471 32759
rect 5365 32521 5399 32555
rect 6101 32521 6135 32555
rect 7389 32521 7423 32555
rect 7573 32521 7607 32555
rect 12909 32521 12943 32555
rect 24041 32521 24075 32555
rect 25506 32521 25540 32555
rect 29929 32521 29963 32555
rect 31861 32521 31895 32555
rect 34529 32521 34563 32555
rect 1869 32453 1903 32487
rect 3617 32453 3651 32487
rect 6529 32453 6563 32487
rect 6745 32453 6779 32487
rect 7757 32453 7791 32487
rect 8769 32453 8803 32487
rect 24685 32453 24719 32487
rect 26433 32453 26467 32487
rect 26617 32453 26651 32487
rect 28181 32453 28215 32487
rect 28365 32453 28399 32487
rect 30297 32453 30331 32487
rect 31125 32453 31159 32487
rect 32873 32453 32907 32487
rect 33701 32453 33735 32487
rect 34253 32453 34287 32487
rect 5181 32385 5215 32419
rect 5457 32385 5491 32419
rect 5733 32385 5767 32419
rect 7448 32385 7482 32419
rect 8585 32385 8619 32419
rect 12265 32385 12299 32419
rect 13093 32385 13127 32419
rect 14197 32385 14231 32419
rect 14841 32385 14875 32419
rect 20269 32385 20303 32419
rect 22017 32385 22051 32419
rect 22293 32385 22327 32419
rect 22477 32385 22511 32419
rect 22753 32385 22787 32419
rect 22845 32385 22879 32419
rect 22937 32385 22971 32419
rect 23121 32385 23155 32419
rect 23397 32385 23431 32419
rect 24225 32385 24259 32419
rect 24409 32385 24443 32419
rect 24869 32385 24903 32419
rect 24961 32385 24995 32419
rect 25058 32385 25092 32419
rect 25329 32385 25363 32419
rect 25421 32385 25455 32419
rect 25605 32385 25639 32419
rect 25789 32385 25823 32419
rect 25973 32385 26007 32419
rect 26065 32385 26099 32419
rect 26249 32385 26283 32419
rect 26341 32385 26375 32419
rect 28825 32385 28859 32419
rect 29009 32385 29043 32419
rect 29988 32385 30022 32419
rect 31217 32385 31251 32419
rect 31677 32385 31711 32419
rect 33977 32385 34011 32419
rect 34161 32385 34195 32419
rect 34345 32385 34379 32419
rect 36369 32385 36403 32419
rect 3893 32317 3927 32351
rect 5825 32317 5859 32351
rect 6929 32317 6963 32351
rect 7021 32317 7055 32351
rect 11529 32317 11563 32351
rect 12541 32317 12575 32351
rect 13277 32317 13311 32351
rect 14473 32317 14507 32351
rect 14749 32317 14783 32351
rect 20177 32317 20211 32351
rect 20361 32317 20395 32351
rect 20453 32317 20487 32351
rect 22109 32317 22143 32351
rect 23673 32317 23707 32351
rect 24317 32317 24351 32351
rect 24501 32317 24535 32351
rect 24777 32317 24811 32351
rect 28457 32317 28491 32351
rect 29469 32317 29503 32351
rect 31585 32317 31619 32351
rect 32689 32317 32723 32351
rect 36093 32317 36127 32351
rect 37473 32317 37507 32351
rect 37565 32317 37599 32351
rect 37657 32317 37691 32351
rect 37749 32317 37783 32351
rect 6377 32249 6411 32283
rect 11989 32249 12023 32283
rect 14657 32249 14691 32283
rect 22201 32249 22235 32283
rect 23213 32249 23247 32283
rect 26801 32249 26835 32283
rect 29561 32249 29595 32283
rect 30113 32249 30147 32283
rect 5181 32181 5215 32215
rect 6561 32181 6595 32215
rect 20637 32181 20671 32215
rect 21833 32181 21867 32215
rect 22569 32181 22603 32215
rect 23581 32181 23615 32215
rect 27997 32181 28031 32215
rect 31585 32181 31619 32215
rect 32137 32181 32171 32215
rect 34621 32181 34655 32215
rect 37289 32181 37323 32215
rect 4537 31977 4571 32011
rect 7849 31977 7883 32011
rect 8585 31977 8619 32011
rect 9045 31977 9079 32011
rect 10977 31977 11011 32011
rect 11069 31977 11103 32011
rect 14657 31977 14691 32011
rect 22569 31977 22603 32011
rect 26617 31977 26651 32011
rect 29837 31977 29871 32011
rect 30941 31977 30975 32011
rect 32137 31977 32171 32011
rect 32229 31977 32263 32011
rect 36093 31977 36127 32011
rect 37859 31977 37893 32011
rect 14105 31909 14139 31943
rect 25605 31909 25639 31943
rect 27445 31909 27479 31943
rect 27721 31909 27755 31943
rect 28733 31909 28767 31943
rect 35449 31909 35483 31943
rect 8033 31841 8067 31875
rect 10425 31841 10459 31875
rect 11621 31841 11655 31875
rect 12081 31841 12115 31875
rect 12909 31841 12943 31875
rect 14749 31841 14783 31875
rect 15209 31841 15243 31875
rect 16129 31841 16163 31875
rect 17233 31841 17267 31875
rect 17509 31841 17543 31875
rect 19349 31841 19383 31875
rect 21097 31841 21131 31875
rect 21741 31841 21775 31875
rect 22845 31841 22879 31875
rect 22937 31841 22971 31875
rect 25053 31841 25087 31875
rect 25513 31841 25547 31875
rect 25973 31841 26007 31875
rect 28457 31841 28491 31875
rect 31677 31841 31711 31875
rect 31861 31841 31895 31875
rect 31953 31841 31987 31875
rect 32597 31841 32631 31875
rect 34805 31841 34839 31875
rect 4813 31773 4847 31807
rect 5733 31773 5767 31807
rect 8125 31773 8159 31807
rect 9137 31773 9171 31807
rect 11529 31773 11563 31807
rect 12173 31773 12207 31807
rect 12540 31773 12574 31807
rect 13369 31773 13403 31807
rect 13737 31773 13771 31807
rect 13921 31773 13955 31807
rect 14230 31773 14264 31807
rect 15301 31773 15335 31807
rect 15945 31773 15979 31807
rect 16313 31773 16347 31807
rect 16405 31773 16439 31807
rect 22201 31773 22235 31807
rect 22745 31773 22779 31807
rect 23029 31773 23063 31807
rect 23397 31773 23431 31807
rect 23581 31773 23615 31807
rect 24961 31773 24995 31807
rect 25237 31773 25271 31807
rect 25421 31773 25455 31807
rect 25697 31773 25731 31807
rect 25881 31773 25915 31807
rect 26065 31773 26099 31807
rect 26436 31773 26470 31807
rect 27261 31773 27295 31807
rect 27629 31773 27663 31807
rect 27859 31773 27893 31807
rect 28089 31773 28123 31807
rect 28272 31773 28306 31807
rect 28365 31773 28399 31807
rect 28641 31773 28675 31807
rect 28825 31773 28859 31807
rect 28917 31773 28951 31807
rect 29561 31773 29595 31807
rect 29745 31773 29779 31807
rect 30481 31773 30515 31807
rect 31125 31773 31159 31807
rect 31217 31773 31251 31807
rect 31401 31773 31435 31807
rect 31493 31773 31527 31807
rect 31769 31773 31803 31807
rect 32413 31773 32447 31807
rect 32505 31773 32539 31807
rect 32689 31773 32723 31807
rect 32873 31773 32907 31807
rect 33057 31773 33091 31807
rect 33241 31773 33275 31807
rect 33333 31773 33367 31807
rect 35541 31773 35575 31807
rect 35817 31773 35851 31807
rect 35909 31773 35943 31807
rect 38117 31773 38151 31807
rect 38301 31773 38335 31807
rect 38485 31773 38519 31807
rect 38577 31773 38611 31807
rect 38669 31773 38703 31807
rect 8769 31705 8803 31739
rect 11437 31705 11471 31739
rect 19625 31705 19659 31739
rect 23765 31705 23799 31739
rect 23949 31705 23983 31739
rect 24133 31705 24167 31739
rect 27997 31705 28031 31739
rect 30665 31705 30699 31739
rect 35725 31705 35759 31739
rect 8401 31637 8435 31671
rect 8569 31637 8603 31671
rect 10517 31637 10551 31671
rect 10609 31637 10643 31671
rect 12633 31637 12667 31671
rect 14289 31637 14323 31671
rect 18981 31637 19015 31671
rect 21189 31637 21223 31671
rect 22385 31637 22419 31671
rect 23213 31637 23247 31671
rect 26433 31637 26467 31671
rect 27077 31637 27111 31671
rect 36369 31637 36403 31671
rect 38853 31637 38887 31671
rect 5733 31433 5767 31467
rect 7389 31433 7423 31467
rect 7665 31433 7699 31467
rect 8677 31433 8711 31467
rect 10977 31433 11011 31467
rect 11713 31433 11747 31467
rect 12725 31433 12759 31467
rect 13553 31433 13587 31467
rect 14105 31433 14139 31467
rect 16773 31433 16807 31467
rect 17969 31433 18003 31467
rect 19717 31433 19751 31467
rect 20085 31433 20119 31467
rect 21373 31433 21407 31467
rect 22569 31433 22603 31467
rect 24041 31433 24075 31467
rect 25881 31433 25915 31467
rect 26157 31433 26191 31467
rect 29653 31433 29687 31467
rect 34463 31433 34497 31467
rect 34713 31433 34747 31467
rect 37105 31433 37139 31467
rect 40233 31433 40267 31467
rect 5365 31365 5399 31399
rect 5581 31365 5615 31399
rect 6377 31365 6411 31399
rect 8953 31365 8987 31399
rect 9045 31365 9079 31399
rect 14289 31365 14323 31399
rect 21281 31365 21315 31399
rect 22201 31365 22235 31399
rect 27471 31365 27505 31399
rect 34253 31365 34287 31399
rect 36159 31365 36193 31399
rect 36277 31365 36311 31399
rect 36921 31365 36955 31399
rect 37565 31365 37599 31399
rect 38761 31365 38795 31399
rect 21971 31331 22005 31365
rect 8309 31297 8343 31331
rect 9321 31297 9355 31331
rect 9965 31297 9999 31331
rect 10425 31297 10459 31331
rect 10885 31297 10919 31331
rect 11710 31297 11744 31331
rect 12081 31297 12115 31331
rect 12173 31297 12207 31331
rect 12909 31297 12943 31331
rect 13001 31297 13035 31331
rect 13277 31297 13311 31331
rect 13369 31297 13403 31331
rect 13553 31297 13587 31331
rect 13737 31297 13771 31331
rect 13891 31297 13925 31331
rect 14197 31297 14231 31331
rect 14381 31297 14415 31331
rect 15577 31297 15611 31331
rect 15945 31297 15979 31331
rect 16681 31297 16715 31331
rect 17141 31297 17175 31331
rect 17509 31297 17543 31331
rect 18245 31297 18279 31331
rect 18521 31297 18555 31331
rect 20729 31297 20763 31331
rect 20821 31297 20855 31331
rect 20913 31297 20947 31331
rect 21097 31297 21131 31331
rect 22293 31297 22327 31331
rect 23121 31297 23155 31331
rect 23305 31297 23339 31331
rect 23673 31297 23707 31331
rect 24869 31297 24903 31331
rect 25237 31297 25271 31331
rect 25789 31297 25823 31331
rect 25973 31297 26007 31331
rect 26433 31297 26467 31331
rect 26525 31297 26559 31331
rect 26617 31297 26651 31331
rect 26801 31297 26835 31331
rect 27169 31297 27203 31331
rect 27261 31297 27295 31331
rect 27353 31297 27387 31331
rect 28273 31297 28307 31331
rect 28457 31297 28491 31331
rect 29561 31297 29595 31331
rect 29745 31297 29779 31331
rect 33425 31297 33459 31331
rect 33701 31297 33735 31331
rect 34897 31297 34931 31331
rect 36001 31297 36035 31331
rect 36369 31297 36403 31331
rect 36461 31297 36495 31331
rect 36645 31297 36679 31331
rect 36737 31297 36771 31331
rect 37289 31297 37323 31331
rect 37473 31297 37507 31331
rect 37657 31297 37691 31331
rect 38485 31297 38519 31331
rect 3249 31229 3283 31263
rect 4997 31229 5031 31263
rect 5273 31229 5307 31263
rect 7113 31229 7147 31263
rect 7548 31229 7582 31263
rect 7757 31229 7791 31263
rect 8033 31229 8067 31263
rect 8401 31229 8435 31263
rect 9413 31229 9447 31263
rect 10701 31229 10735 31263
rect 11161 31229 11195 31263
rect 11345 31229 11379 31263
rect 15117 31229 15151 31263
rect 15393 31229 15427 31263
rect 15853 31229 15887 31263
rect 17233 31229 17267 31263
rect 17417 31229 17451 31263
rect 18153 31229 18187 31263
rect 18613 31229 18647 31263
rect 18797 31229 18831 31263
rect 19349 31229 19383 31263
rect 20177 31229 20211 31263
rect 20361 31229 20395 31263
rect 22569 31229 22603 31263
rect 23857 31229 23891 31263
rect 24133 31229 24167 31263
rect 24961 31229 24995 31263
rect 25329 31229 25363 31263
rect 27629 31229 27663 31263
rect 33241 31229 33275 31263
rect 35081 31229 35115 31263
rect 9873 31161 9907 31195
rect 15209 31161 15243 31195
rect 26985 31161 27019 31195
rect 27813 31161 27847 31195
rect 27905 31161 27939 31195
rect 5549 31093 5583 31127
rect 9597 31093 9631 31127
rect 11529 31093 11563 31127
rect 13185 31093 13219 31127
rect 20545 31093 20579 31127
rect 21833 31093 21867 31127
rect 22017 31093 22051 31127
rect 22385 31093 22419 31127
rect 24317 31093 24351 31127
rect 28549 31093 28583 31127
rect 33609 31093 33643 31127
rect 34437 31093 34471 31127
rect 34621 31093 34655 31127
rect 37841 31093 37875 31127
rect 4169 30889 4203 30923
rect 7941 30889 7975 30923
rect 8585 30889 8619 30923
rect 10793 30889 10827 30923
rect 11345 30889 11379 30923
rect 15209 30889 15243 30923
rect 18429 30889 18463 30923
rect 18705 30889 18739 30923
rect 18889 30889 18923 30923
rect 22845 30889 22879 30923
rect 23121 30889 23155 30923
rect 23305 30889 23339 30923
rect 23673 30889 23707 30923
rect 24593 30889 24627 30923
rect 26617 30889 26651 30923
rect 33609 30889 33643 30923
rect 35173 30889 35207 30923
rect 35725 30889 35759 30923
rect 36921 30889 36955 30923
rect 38025 30889 38059 30923
rect 17969 30821 18003 30855
rect 27813 30821 27847 30855
rect 30389 30821 30423 30855
rect 34989 30821 35023 30855
rect 38209 30821 38243 30855
rect 4629 30753 4663 30787
rect 4813 30753 4847 30787
rect 7389 30753 7423 30787
rect 9689 30753 9723 30787
rect 19349 30753 19383 30787
rect 20821 30753 20855 30787
rect 21097 30753 21131 30787
rect 35357 30753 35391 30787
rect 36277 30753 36311 30787
rect 37749 30753 37783 30787
rect 3617 30685 3651 30719
rect 4537 30685 4571 30719
rect 6101 30685 6135 30719
rect 8033 30685 8067 30719
rect 8217 30685 8251 30719
rect 8401 30685 8435 30719
rect 8585 30685 8619 30719
rect 9873 30685 9907 30719
rect 10333 30685 10367 30719
rect 10701 30685 10735 30719
rect 10974 30685 11008 30719
rect 11437 30685 11471 30719
rect 13093 30685 13127 30719
rect 13277 30685 13311 30719
rect 15209 30685 15243 30719
rect 15301 30685 15335 30719
rect 15485 30685 15519 30719
rect 15577 30685 15611 30719
rect 15669 30685 15703 30719
rect 17785 30685 17819 30719
rect 17969 30685 18003 30719
rect 18061 30685 18095 30719
rect 21741 30685 21775 30719
rect 23213 30685 23247 30719
rect 23581 30685 23615 30719
rect 23857 30685 23891 30719
rect 23949 30685 23983 30719
rect 26893 30685 26927 30719
rect 27537 30685 27571 30719
rect 27721 30685 27755 30719
rect 28733 30685 28767 30719
rect 29009 30685 29043 30719
rect 29561 30685 29595 30719
rect 30849 30685 30883 30719
rect 31125 30685 31159 30719
rect 31217 30685 31251 30719
rect 31309 30685 31343 30719
rect 31493 30685 31527 30719
rect 31585 30685 31619 30719
rect 31769 30685 31803 30719
rect 33793 30685 33827 30719
rect 33885 30685 33919 30719
rect 34253 30685 34287 30719
rect 35173 30685 35207 30719
rect 35725 30685 35759 30719
rect 35909 30685 35943 30719
rect 36645 30685 36679 30719
rect 36829 30685 36863 30719
rect 36921 30685 36955 30719
rect 37105 30685 37139 30719
rect 37381 30685 37415 30719
rect 38485 30685 38519 30719
rect 1593 30617 1627 30651
rect 3341 30617 3375 30651
rect 7573 30617 7607 30651
rect 8125 30617 8159 30651
rect 18245 30617 18279 30651
rect 18521 30617 18555 30651
rect 18737 30617 18771 30651
rect 21925 30617 21959 30651
rect 24501 30617 24535 30651
rect 26617 30617 26651 30651
rect 26801 30617 26835 30651
rect 28365 30617 28399 30651
rect 28549 30617 28583 30651
rect 30665 30617 30699 30651
rect 31677 30617 31711 30651
rect 33977 30617 34011 30651
rect 34115 30617 34149 30651
rect 35633 30617 35667 30651
rect 37866 30617 37900 30651
rect 38393 30617 38427 30651
rect 38945 30617 38979 30651
rect 6193 30549 6227 30583
rect 7481 30549 7515 30583
rect 10977 30549 11011 30583
rect 13277 30549 13311 30583
rect 21649 30549 21683 30583
rect 23489 30549 23523 30583
rect 28825 30549 28859 30583
rect 30205 30549 30239 30583
rect 31401 30549 31435 30583
rect 36645 30549 36679 30583
rect 37657 30549 37691 30583
rect 3065 30345 3099 30379
rect 4537 30345 4571 30379
rect 10609 30345 10643 30379
rect 14473 30345 14507 30379
rect 18337 30345 18371 30379
rect 2697 30277 2731 30311
rect 12357 30277 12391 30311
rect 23213 30277 23247 30311
rect 25881 30277 25915 30311
rect 30665 30277 30699 30311
rect 31033 30277 31067 30311
rect 31661 30277 31695 30311
rect 31861 30277 31895 30311
rect 33793 30277 33827 30311
rect 38025 30277 38059 30311
rect 1501 30209 1535 30243
rect 2881 30209 2915 30243
rect 3157 30209 3191 30243
rect 7389 30209 7423 30243
rect 10885 30209 10919 30243
rect 12055 30209 12089 30243
rect 12449 30209 12483 30243
rect 12909 30209 12943 30243
rect 13461 30209 13495 30243
rect 13737 30209 13771 30243
rect 13921 30209 13955 30243
rect 14013 30209 14047 30243
rect 14289 30209 14323 30243
rect 14657 30209 14691 30243
rect 14933 30209 14967 30243
rect 15209 30209 15243 30243
rect 15393 30209 15427 30243
rect 15761 30209 15795 30243
rect 15945 30209 15979 30243
rect 16037 30209 16071 30243
rect 16221 30209 16255 30243
rect 16313 30209 16347 30243
rect 16425 30215 16459 30249
rect 16957 30209 16991 30243
rect 18705 30209 18739 30243
rect 23075 30209 23109 30243
rect 23305 30209 23339 30243
rect 23433 30209 23467 30243
rect 23581 30209 23615 30243
rect 26433 30209 26467 30243
rect 26525 30209 26559 30243
rect 30297 30209 30331 30243
rect 30455 30209 30489 30243
rect 30573 30209 30607 30243
rect 30757 30209 30791 30243
rect 31217 30209 31251 30243
rect 31401 30209 31435 30243
rect 32137 30209 32171 30243
rect 32413 30209 32447 30243
rect 32505 30209 32539 30243
rect 34437 30209 34471 30243
rect 36277 30209 36311 30243
rect 37289 30209 37323 30243
rect 37565 30209 37599 30243
rect 37933 30209 37967 30243
rect 38117 30209 38151 30243
rect 38209 30209 38243 30243
rect 4629 30141 4663 30175
rect 4813 30141 4847 30175
rect 11897 30141 11931 30175
rect 12725 30141 12759 30175
rect 13369 30141 13403 30175
rect 16681 30141 16715 30175
rect 18613 30141 18647 30175
rect 25513 30141 25547 30175
rect 26249 30141 26283 30175
rect 28457 30141 28491 30175
rect 29929 30141 29963 30175
rect 30205 30141 30239 30175
rect 32229 30141 32263 30175
rect 34253 30141 34287 30175
rect 36369 30141 36403 30175
rect 38485 30141 38519 30175
rect 40233 30141 40267 30175
rect 1777 30073 1811 30107
rect 15025 30073 15059 30107
rect 18245 30073 18279 30107
rect 26341 30073 26375 30107
rect 30941 30073 30975 30107
rect 31493 30073 31527 30107
rect 32137 30073 32171 30107
rect 33425 30073 33459 30107
rect 4169 30005 4203 30039
rect 7481 30005 7515 30039
rect 14197 30005 14231 30039
rect 16037 30005 16071 30039
rect 16773 30005 16807 30039
rect 17141 30005 17175 30039
rect 18613 30005 18647 30039
rect 22937 30005 22971 30039
rect 25881 30005 25915 30039
rect 26065 30005 26099 30039
rect 31677 30005 31711 30039
rect 32597 30005 32631 30039
rect 33793 30005 33827 30039
rect 33977 30005 34011 30039
rect 34621 30005 34655 30039
rect 36277 30005 36311 30039
rect 36645 30005 36679 30039
rect 37381 30005 37415 30039
rect 37841 30005 37875 30039
rect 5549 29801 5583 29835
rect 10517 29801 10551 29835
rect 18337 29801 18371 29835
rect 35817 29801 35851 29835
rect 36001 29801 36035 29835
rect 38393 29801 38427 29835
rect 12541 29733 12575 29767
rect 13553 29733 13587 29767
rect 14381 29733 14415 29767
rect 19625 29733 19659 29767
rect 27169 29733 27203 29767
rect 27261 29733 27295 29767
rect 34897 29733 34931 29767
rect 36369 29733 36403 29767
rect 38485 29733 38519 29767
rect 4077 29665 4111 29699
rect 6285 29665 6319 29699
rect 9873 29665 9907 29699
rect 10241 29665 10275 29699
rect 10333 29665 10367 29699
rect 12173 29665 12207 29699
rect 14197 29665 14231 29699
rect 15485 29665 15519 29699
rect 25237 29665 25271 29699
rect 30573 29665 30607 29699
rect 32505 29665 32539 29699
rect 33149 29665 33183 29699
rect 33241 29665 33275 29699
rect 35081 29665 35115 29699
rect 3801 29597 3835 29631
rect 6101 29597 6135 29631
rect 10609 29597 10643 29631
rect 11161 29597 11195 29631
rect 11437 29597 11471 29631
rect 11805 29597 11839 29631
rect 11970 29597 12004 29631
rect 12081 29597 12115 29631
rect 12357 29597 12391 29631
rect 12725 29597 12759 29631
rect 12909 29597 12943 29631
rect 13369 29597 13403 29631
rect 13461 29597 13495 29631
rect 13645 29597 13679 29631
rect 14105 29597 14139 29631
rect 14289 29597 14323 29631
rect 14381 29597 14415 29631
rect 14565 29597 14599 29631
rect 15117 29597 15151 29631
rect 15577 29597 15611 29631
rect 15945 29597 15979 29631
rect 16129 29597 16163 29631
rect 16497 29597 16531 29631
rect 16865 29597 16899 29631
rect 17141 29597 17175 29631
rect 17877 29597 17911 29631
rect 18521 29597 18555 29631
rect 18797 29597 18831 29631
rect 18889 29597 18923 29631
rect 19073 29597 19107 29631
rect 22293 29597 22327 29631
rect 22661 29597 22695 29631
rect 22845 29597 22879 29631
rect 23121 29597 23155 29631
rect 23213 29597 23247 29631
rect 23397 29597 23431 29631
rect 23489 29597 23523 29631
rect 23765 29597 23799 29631
rect 23949 29597 23983 29631
rect 24777 29597 24811 29631
rect 25145 29597 25179 29631
rect 25329 29597 25363 29631
rect 25789 29597 25823 29631
rect 25973 29597 26007 29631
rect 26249 29597 26283 29631
rect 26525 29597 26559 29631
rect 26617 29597 26651 29631
rect 27813 29597 27847 29631
rect 28181 29597 28215 29631
rect 28365 29597 28399 29631
rect 28825 29597 28859 29631
rect 30481 29597 30515 29631
rect 30665 29597 30699 29631
rect 32781 29597 32815 29631
rect 32873 29597 32907 29631
rect 34069 29597 34103 29631
rect 34161 29597 34195 29631
rect 34713 29597 34747 29631
rect 34897 29597 34931 29631
rect 35173 29597 35207 29631
rect 36277 29597 36311 29631
rect 36461 29597 36495 29631
rect 36553 29597 36587 29631
rect 38117 29597 38151 29631
rect 38669 29597 38703 29631
rect 39037 29597 39071 29631
rect 39129 29597 39163 29631
rect 39497 29597 39531 29631
rect 11713 29529 11747 29563
rect 12817 29529 12851 29563
rect 19257 29529 19291 29563
rect 19441 29529 19475 29563
rect 22385 29529 22419 29563
rect 24593 29529 24627 29563
rect 27077 29529 27111 29563
rect 32229 29529 32263 29563
rect 32597 29529 32631 29563
rect 33885 29529 33919 29563
rect 34437 29529 34471 29563
rect 35633 29529 35667 29563
rect 35849 29529 35883 29563
rect 36093 29529 36127 29563
rect 37565 29529 37599 29563
rect 37933 29529 37967 29563
rect 38393 29529 38427 29563
rect 38761 29529 38795 29563
rect 38853 29529 38887 29563
rect 39589 29529 39623 29563
rect 5641 29461 5675 29495
rect 6009 29461 6043 29495
rect 13185 29461 13219 29495
rect 15209 29461 15243 29495
rect 16313 29461 16347 29495
rect 18613 29461 18647 29495
rect 22937 29461 22971 29495
rect 23581 29461 23615 29495
rect 24501 29461 24535 29495
rect 24961 29461 24995 29495
rect 30757 29461 30791 29495
rect 32965 29461 32999 29495
rect 34253 29461 34287 29495
rect 38209 29461 38243 29495
rect 39313 29461 39347 29495
rect 11345 29257 11379 29291
rect 12081 29257 12115 29291
rect 16681 29257 16715 29291
rect 18705 29257 18739 29291
rect 19533 29257 19567 29291
rect 27261 29257 27295 29291
rect 27905 29257 27939 29291
rect 32229 29257 32263 29291
rect 35449 29257 35483 29291
rect 9781 29189 9815 29223
rect 11529 29189 11563 29223
rect 12541 29189 12575 29223
rect 19349 29189 19383 29223
rect 28575 29189 28609 29223
rect 31769 29189 31803 29223
rect 32505 29189 32539 29223
rect 32597 29189 32631 29223
rect 35541 29189 35575 29223
rect 35633 29189 35667 29223
rect 35909 29189 35943 29223
rect 36721 29189 36755 29223
rect 36921 29189 36955 29223
rect 38485 29189 38519 29223
rect 40233 29189 40267 29223
rect 4445 29121 4479 29155
rect 9413 29121 9447 29155
rect 9873 29121 9907 29155
rect 10149 29121 10183 29155
rect 10241 29121 10275 29155
rect 10977 29121 11011 29155
rect 11621 29121 11655 29155
rect 11897 29121 11931 29155
rect 12449 29121 12483 29155
rect 15117 29121 15151 29155
rect 15485 29121 15519 29155
rect 15853 29121 15887 29155
rect 15945 29121 15979 29155
rect 16865 29121 16899 29155
rect 17049 29121 17083 29155
rect 17141 29121 17175 29155
rect 17601 29121 17635 29155
rect 17877 29121 17911 29155
rect 19533 29121 19567 29155
rect 19717 29121 19751 29155
rect 20913 29121 20947 29155
rect 21097 29121 21131 29155
rect 21557 29121 21591 29155
rect 22109 29121 22143 29155
rect 23121 29121 23155 29155
rect 23305 29121 23339 29155
rect 23581 29121 23615 29155
rect 23857 29121 23891 29155
rect 24041 29121 24075 29155
rect 24133 29121 24167 29155
rect 24409 29121 24443 29155
rect 24593 29121 24627 29155
rect 24777 29121 24811 29155
rect 24869 29121 24903 29155
rect 25053 29121 25087 29155
rect 25421 29121 25455 29155
rect 25605 29121 25639 29155
rect 25697 29121 25731 29155
rect 25881 29121 25915 29155
rect 26433 29121 26467 29155
rect 26617 29121 26651 29155
rect 27169 29121 27203 29155
rect 27537 29121 27571 29155
rect 28273 29121 28307 29155
rect 28365 29121 28399 29155
rect 28457 29121 28491 29155
rect 29009 29121 29043 29155
rect 31953 29121 31987 29155
rect 32408 29121 32442 29155
rect 32725 29121 32759 29155
rect 32873 29121 32907 29155
rect 33608 29121 33642 29155
rect 33701 29121 33735 29155
rect 34069 29121 34103 29155
rect 34621 29121 34655 29155
rect 34989 29121 35023 29155
rect 36001 29121 36035 29155
rect 36185 29121 36219 29155
rect 36369 29121 36403 29155
rect 37289 29121 37323 29155
rect 37473 29121 37507 29155
rect 37565 29121 37599 29155
rect 37749 29121 37783 29155
rect 38209 29121 38243 29155
rect 6837 29053 6871 29087
rect 7113 29053 7147 29087
rect 9229 29053 9263 29087
rect 9597 29053 9631 29087
rect 10701 29053 10735 29087
rect 10885 29053 10919 29087
rect 12633 29053 12667 29087
rect 15025 29053 15059 29087
rect 15301 29053 15335 29087
rect 17325 29053 17359 29087
rect 18981 29053 19015 29087
rect 21281 29053 21315 29087
rect 22017 29053 22051 29087
rect 22477 29053 22511 29087
rect 23397 29053 23431 29087
rect 24225 29053 24259 29087
rect 24685 29053 24719 29087
rect 25145 29053 25179 29087
rect 25237 29053 25271 29087
rect 27445 29053 27479 29087
rect 28089 29053 28123 29087
rect 28733 29053 28767 29087
rect 33793 29053 33827 29087
rect 34437 29053 34471 29087
rect 37657 29053 37691 29087
rect 6193 28985 6227 29019
rect 8585 28985 8619 29019
rect 9965 28985 9999 29019
rect 16957 28985 16991 29019
rect 19073 28985 19107 29019
rect 20729 28985 20763 29019
rect 21833 28985 21867 29019
rect 23213 28985 23247 29019
rect 25697 28985 25731 29019
rect 26801 28985 26835 29019
rect 27629 28985 27663 29019
rect 28825 28985 28859 29019
rect 31585 28985 31619 29019
rect 33885 28985 33919 29019
rect 34897 28985 34931 29019
rect 35265 28985 35299 29019
rect 35817 28985 35851 29019
rect 36553 28985 36587 29019
rect 37289 28985 37323 29019
rect 4708 28917 4742 28951
rect 8677 28917 8711 28951
rect 9505 28917 9539 28951
rect 9597 28917 9631 28951
rect 10425 28917 10459 28951
rect 19184 28917 19218 28951
rect 22937 28917 22971 28951
rect 23673 28917 23707 28951
rect 33517 28917 33551 28951
rect 34253 28917 34287 28951
rect 36737 28917 36771 28951
rect 7573 28713 7607 28747
rect 11161 28713 11195 28747
rect 12081 28713 12115 28747
rect 21925 28713 21959 28747
rect 24041 28713 24075 28747
rect 24501 28713 24535 28747
rect 26249 28713 26283 28747
rect 26709 28713 26743 28747
rect 34253 28713 34287 28747
rect 35173 28713 35207 28747
rect 38209 28713 38243 28747
rect 10425 28645 10459 28679
rect 23857 28645 23891 28679
rect 5549 28577 5583 28611
rect 8217 28577 8251 28611
rect 10057 28577 10091 28611
rect 10609 28577 10643 28611
rect 17325 28577 17359 28611
rect 17877 28577 17911 28611
rect 23673 28577 23707 28611
rect 25237 28577 25271 28611
rect 25697 28577 25731 28611
rect 26249 28577 26283 28611
rect 26847 28577 26881 28611
rect 32873 28577 32907 28611
rect 38393 28577 38427 28611
rect 38853 28577 38887 28611
rect 8033 28509 8067 28543
rect 9781 28509 9815 28543
rect 10425 28509 10459 28543
rect 10885 28509 10919 28543
rect 11161 28509 11195 28543
rect 11805 28509 11839 28543
rect 11897 28509 11931 28543
rect 12173 28509 12207 28543
rect 14289 28509 14323 28543
rect 14657 28509 14691 28543
rect 17785 28509 17819 28543
rect 21189 28509 21223 28543
rect 22109 28509 22143 28543
rect 22201 28509 22235 28543
rect 22385 28509 22419 28543
rect 22477 28509 22511 28543
rect 23029 28509 23063 28543
rect 23305 28509 23339 28543
rect 23489 28509 23523 28543
rect 24777 28509 24811 28543
rect 24869 28509 24903 28543
rect 24961 28509 24995 28543
rect 25145 28509 25179 28543
rect 25421 28509 25455 28543
rect 25513 28509 25547 28543
rect 25789 28509 25823 28543
rect 26065 28509 26099 28543
rect 26341 28509 26375 28543
rect 26525 28509 26559 28543
rect 26985 28509 27019 28543
rect 27629 28509 27663 28543
rect 27997 28509 28031 28543
rect 28273 28509 28307 28543
rect 28641 28509 28675 28543
rect 29745 28509 29779 28543
rect 29929 28509 29963 28543
rect 30113 28509 30147 28543
rect 30205 28509 30239 28543
rect 32137 28509 32171 28543
rect 32597 28509 32631 28543
rect 33609 28509 33643 28543
rect 33885 28509 33919 28543
rect 35725 28509 35759 28543
rect 36001 28509 36035 28543
rect 38485 28509 38519 28543
rect 5825 28441 5859 28475
rect 9487 28441 9521 28475
rect 10793 28441 10827 28475
rect 11069 28441 11103 28475
rect 14381 28441 14415 28475
rect 14473 28441 14507 28475
rect 24225 28441 24259 28475
rect 29837 28441 29871 28475
rect 30481 28441 30515 28475
rect 34161 28441 34195 28475
rect 35173 28441 35207 28475
rect 35357 28441 35391 28475
rect 38761 28441 38795 28475
rect 7297 28373 7331 28407
rect 7941 28373 7975 28407
rect 9965 28373 9999 28407
rect 11621 28373 11655 28407
rect 14105 28373 14139 28407
rect 21005 28373 21039 28407
rect 23121 28373 23155 28407
rect 23397 28373 23431 28407
rect 24025 28373 24059 28407
rect 25881 28373 25915 28407
rect 26525 28373 26559 28407
rect 28549 28373 28583 28407
rect 29561 28373 29595 28407
rect 30573 28373 30607 28407
rect 33609 28373 33643 28407
rect 34989 28373 35023 28407
rect 35909 28373 35943 28407
rect 4261 28169 4295 28203
rect 6377 28169 6411 28203
rect 25421 28169 25455 28203
rect 25789 28169 25823 28203
rect 32505 28169 32539 28203
rect 4813 28101 4847 28135
rect 13921 28101 13955 28135
rect 14565 28101 14599 28135
rect 15669 28101 15703 28135
rect 15761 28101 15795 28135
rect 16957 28101 16991 28135
rect 17049 28101 17083 28135
rect 19257 28101 19291 28135
rect 21281 28101 21315 28135
rect 30849 28101 30883 28135
rect 31401 28101 31435 28135
rect 4721 28033 4755 28067
rect 6745 28033 6779 28067
rect 11713 28033 11747 28067
rect 11897 28033 11931 28067
rect 12081 28033 12115 28067
rect 12817 28033 12851 28067
rect 12910 28033 12944 28067
rect 13093 28033 13127 28067
rect 13185 28033 13219 28067
rect 13323 28033 13357 28067
rect 13553 28033 13587 28067
rect 13646 28033 13680 28067
rect 13829 28033 13863 28067
rect 14059 28033 14093 28067
rect 14468 28033 14502 28067
rect 14657 28033 14691 28067
rect 14795 28033 14829 28067
rect 14933 28033 14967 28067
rect 15393 28033 15427 28067
rect 15486 28033 15520 28067
rect 15877 28033 15911 28067
rect 16681 28033 16715 28067
rect 16774 28033 16808 28067
rect 17187 28033 17221 28067
rect 18429 28033 18463 28067
rect 18613 28033 18647 28067
rect 18889 28033 18923 28067
rect 19073 28033 19107 28067
rect 19533 28033 19567 28067
rect 19809 28033 19843 28067
rect 19993 28033 20027 28067
rect 20177 28033 20211 28067
rect 20637 28033 20671 28067
rect 21373 28033 21407 28067
rect 21833 28033 21867 28067
rect 22109 28033 22143 28067
rect 22385 28033 22419 28067
rect 22569 28033 22603 28067
rect 22845 28033 22879 28067
rect 23029 28033 23063 28067
rect 25145 28033 25179 28067
rect 28825 28033 28859 28067
rect 31309 28033 31343 28067
rect 32321 28033 32355 28067
rect 32689 28033 32723 28067
rect 2513 27965 2547 27999
rect 2789 27965 2823 27999
rect 4997 27965 5031 27999
rect 6837 27965 6871 27999
rect 7021 27965 7055 27999
rect 18245 27965 18279 27999
rect 19441 27965 19475 27999
rect 20085 27965 20119 27999
rect 20821 27965 20855 27999
rect 21557 27965 21591 27999
rect 22201 27965 22235 27999
rect 25513 27965 25547 27999
rect 25630 27965 25664 27999
rect 29193 27965 29227 27999
rect 4353 27897 4387 27931
rect 11713 27897 11747 27931
rect 14197 27897 14231 27931
rect 20913 27897 20947 27931
rect 13461 27829 13495 27863
rect 14289 27829 14323 27863
rect 16037 27829 16071 27863
rect 17325 27829 17359 27863
rect 18705 27829 18739 27863
rect 20453 27829 20487 27863
rect 23029 27829 23063 27863
rect 30619 27829 30653 27863
rect 31125 27829 31159 27863
rect 32781 27829 32815 27863
rect 7284 27625 7318 27659
rect 11345 27625 11379 27659
rect 17693 27625 17727 27659
rect 17877 27625 17911 27659
rect 36645 27625 36679 27659
rect 37289 27625 37323 27659
rect 5549 27557 5583 27591
rect 13001 27557 13035 27591
rect 18337 27557 18371 27591
rect 30941 27557 30975 27591
rect 33517 27557 33551 27591
rect 3801 27489 3835 27523
rect 7021 27489 7055 27523
rect 8769 27489 8803 27523
rect 9597 27489 9631 27523
rect 9689 27489 9723 27523
rect 12449 27489 12483 27523
rect 13185 27489 13219 27523
rect 13829 27489 13863 27523
rect 29745 27489 29779 27523
rect 31033 27489 31067 27523
rect 32137 27489 32171 27523
rect 33332 27489 33366 27523
rect 37105 27489 37139 27523
rect 39313 27489 39347 27523
rect 11069 27421 11103 27455
rect 12541 27421 12575 27455
rect 13277 27421 13311 27455
rect 13369 27421 13403 27455
rect 13461 27421 13495 27455
rect 13737 27421 13771 27455
rect 13921 27421 13955 27455
rect 14289 27421 14323 27455
rect 14381 27421 14415 27455
rect 14565 27421 14599 27455
rect 14657 27421 14691 27455
rect 14749 27421 14783 27455
rect 15209 27421 15243 27455
rect 15302 27421 15336 27455
rect 15485 27421 15519 27455
rect 15577 27421 15611 27455
rect 15715 27421 15749 27455
rect 17325 27421 17359 27455
rect 17509 27421 17543 27455
rect 18612 27399 18646 27433
rect 18705 27421 18739 27455
rect 18797 27421 18831 27455
rect 18981 27421 19015 27455
rect 19533 27421 19567 27455
rect 20453 27421 20487 27455
rect 20637 27421 20671 27455
rect 25421 27421 25455 27455
rect 25513 27421 25547 27455
rect 29929 27421 29963 27455
rect 30757 27421 30791 27455
rect 32295 27421 32329 27455
rect 32597 27421 32631 27455
rect 33057 27421 33091 27455
rect 33149 27421 33183 27455
rect 33241 27421 33275 27455
rect 36645 27421 36679 27455
rect 36829 27421 36863 27455
rect 37381 27421 37415 27455
rect 4077 27353 4111 27387
rect 17831 27353 17865 27387
rect 18245 27353 18279 27387
rect 19901 27353 19935 27387
rect 25697 27353 25731 27387
rect 31217 27353 31251 27387
rect 32413 27353 32447 27387
rect 32505 27353 32539 27387
rect 39589 27353 39623 27387
rect 9119 27285 9153 27319
rect 9597 27285 9631 27319
rect 14473 27285 14507 27319
rect 15853 27285 15887 27319
rect 17233 27285 17267 27319
rect 19349 27285 19383 27319
rect 19625 27285 19659 27319
rect 19717 27285 19751 27319
rect 20269 27285 20303 27319
rect 25421 27285 25455 27319
rect 32781 27285 32815 27319
rect 37013 27285 37047 27319
rect 37105 27285 37139 27319
rect 3985 27081 4019 27115
rect 4353 27081 4387 27115
rect 4445 27081 4479 27115
rect 8401 27081 8435 27115
rect 8769 27081 8803 27115
rect 9781 27081 9815 27115
rect 10241 27081 10275 27115
rect 11161 27081 11195 27115
rect 11713 27081 11747 27115
rect 13553 27081 13587 27115
rect 16681 27081 16715 27115
rect 19809 27081 19843 27115
rect 20177 27081 20211 27115
rect 20821 27081 20855 27115
rect 22569 27081 22603 27115
rect 29837 27081 29871 27115
rect 30205 27081 30239 27115
rect 31217 27081 31251 27115
rect 31401 27081 31435 27115
rect 38117 27081 38151 27115
rect 40049 27081 40083 27115
rect 6469 27013 6503 27047
rect 6653 27013 6687 27047
rect 10701 27013 10735 27047
rect 17509 27013 17543 27047
rect 18981 27013 19015 27047
rect 19625 27013 19659 27047
rect 23213 27013 23247 27047
rect 24869 27013 24903 27047
rect 32137 27013 32171 27047
rect 32321 27013 32355 27047
rect 36461 27013 36495 27047
rect 37565 27013 37599 27047
rect 39221 27013 39255 27047
rect 39405 27013 39439 27047
rect 5641 26945 5675 26979
rect 5825 26945 5859 26979
rect 5917 26945 5951 26979
rect 6009 26945 6043 26979
rect 6837 26945 6871 26979
rect 8861 26945 8895 26979
rect 9689 26945 9723 26979
rect 9873 26945 9907 26979
rect 10149 26945 10183 26979
rect 10333 26945 10367 26979
rect 10425 26945 10459 26979
rect 10517 26945 10551 26979
rect 10793 26945 10827 26979
rect 11529 26945 11563 26979
rect 13369 26945 13403 26979
rect 13645 26945 13679 26979
rect 14933 26945 14967 26979
rect 15301 26945 15335 26979
rect 15485 26945 15519 26979
rect 16819 26945 16853 26979
rect 16957 26945 16991 26979
rect 17049 26945 17083 26979
rect 17232 26945 17266 26979
rect 17325 26945 17359 26979
rect 17693 26945 17727 26979
rect 17877 26945 17911 26979
rect 18337 26945 18371 26979
rect 18429 26945 18463 26979
rect 18521 26945 18555 26979
rect 18613 26945 18647 26979
rect 19165 26945 19199 26979
rect 19809 26945 19843 26979
rect 19993 26945 20027 26979
rect 20085 26945 20119 26979
rect 20361 26945 20395 26979
rect 20545 26945 20579 26979
rect 21097 26945 21131 26979
rect 22017 26945 22051 26979
rect 22201 26945 22235 26979
rect 22477 26945 22511 26979
rect 22661 26945 22695 26979
rect 22937 26945 22971 26979
rect 23305 26945 23339 26979
rect 24501 26945 24535 26979
rect 24777 26945 24811 26979
rect 25605 26945 25639 26979
rect 25789 26945 25823 26979
rect 25881 26945 25915 26979
rect 30849 26945 30883 26979
rect 31677 26945 31711 26979
rect 31769 26945 31803 26979
rect 34437 26945 34471 26979
rect 34621 26945 34655 26979
rect 36185 26945 36219 26979
rect 36277 26945 36311 26979
rect 36553 26945 36587 26979
rect 36737 26945 36771 26979
rect 36829 26945 36863 26979
rect 36921 26945 36955 26979
rect 37473 26945 37507 26979
rect 37657 26945 37691 26979
rect 37775 26945 37809 26979
rect 37933 26945 37967 26979
rect 38393 26945 38427 26979
rect 38669 26945 38703 26979
rect 38945 26945 38979 26979
rect 39681 26945 39715 26979
rect 40233 26945 40267 26979
rect 4629 26877 4663 26911
rect 8953 26877 8987 26911
rect 10628 26877 10662 26911
rect 10885 26877 10919 26911
rect 11897 26877 11931 26911
rect 14841 26877 14875 26911
rect 15025 26877 15059 26911
rect 15117 26877 15151 26911
rect 18797 26877 18831 26911
rect 19257 26877 19291 26911
rect 20913 26877 20947 26911
rect 21373 26877 21407 26911
rect 23029 26877 23063 26911
rect 23397 26877 23431 26911
rect 24409 26877 24443 26911
rect 25421 26877 25455 26911
rect 30297 26877 30331 26911
rect 30389 26877 30423 26911
rect 38761 26877 38795 26911
rect 38853 26877 38887 26911
rect 13369 26809 13403 26843
rect 15393 26809 15427 26843
rect 21833 26809 21867 26843
rect 23673 26809 23707 26843
rect 31861 26809 31895 26843
rect 36461 26809 36495 26843
rect 37105 26809 37139 26843
rect 39129 26809 39163 26843
rect 6193 26741 6227 26775
rect 10793 26741 10827 26775
rect 12081 26741 12115 26775
rect 14657 26741 14691 26775
rect 20453 26741 20487 26775
rect 21281 26741 21315 26775
rect 22753 26741 22787 26775
rect 22937 26741 22971 26775
rect 23305 26741 23339 26775
rect 24225 26741 24259 26775
rect 31217 26741 31251 26775
rect 32321 26741 32355 26775
rect 32505 26741 32539 26775
rect 34621 26741 34655 26775
rect 37289 26741 37323 26775
rect 39405 26741 39439 26775
rect 6653 26537 6687 26571
rect 8677 26537 8711 26571
rect 10609 26537 10643 26571
rect 10977 26537 11011 26571
rect 11253 26537 11287 26571
rect 12081 26537 12115 26571
rect 12265 26537 12299 26571
rect 12633 26537 12667 26571
rect 16865 26537 16899 26571
rect 18613 26537 18647 26571
rect 20269 26537 20303 26571
rect 22477 26537 22511 26571
rect 23489 26537 23523 26571
rect 24409 26537 24443 26571
rect 24593 26537 24627 26571
rect 24961 26537 24995 26571
rect 25421 26537 25455 26571
rect 25697 26537 25731 26571
rect 26801 26537 26835 26571
rect 28457 26537 28491 26571
rect 29745 26537 29779 26571
rect 31493 26537 31527 26571
rect 34529 26537 34563 26571
rect 34989 26537 35023 26571
rect 40049 26537 40083 26571
rect 5917 26469 5951 26503
rect 8953 26469 8987 26503
rect 10149 26469 10183 26503
rect 11989 26469 12023 26503
rect 14105 26469 14139 26503
rect 20545 26469 20579 26503
rect 25513 26469 25547 26503
rect 29009 26469 29043 26503
rect 32413 26469 32447 26503
rect 34713 26469 34747 26503
rect 37749 26469 37783 26503
rect 3157 26401 3191 26435
rect 3341 26401 3375 26435
rect 6745 26401 6779 26435
rect 18797 26401 18831 26435
rect 20637 26401 20671 26435
rect 20729 26401 20763 26435
rect 21189 26401 21223 26435
rect 22293 26401 22327 26435
rect 22661 26401 22695 26435
rect 22753 26401 22787 26435
rect 26709 26401 26743 26435
rect 27629 26401 27663 26435
rect 28089 26401 28123 26435
rect 28733 26401 28767 26435
rect 38025 26401 38059 26435
rect 38117 26401 38151 26435
rect 4353 26333 4387 26367
rect 5365 26333 5399 26367
rect 5733 26333 5767 26367
rect 6009 26333 6043 26367
rect 6102 26333 6136 26367
rect 6515 26333 6549 26367
rect 6929 26333 6963 26367
rect 8033 26333 8067 26367
rect 8181 26333 8215 26367
rect 8401 26333 8435 26367
rect 8539 26333 8573 26367
rect 9321 26333 9355 26367
rect 9873 26333 9907 26367
rect 9965 26333 9999 26367
rect 10149 26333 10183 26367
rect 10609 26333 10643 26367
rect 10793 26333 10827 26367
rect 11253 26333 11287 26367
rect 11437 26333 11471 26367
rect 12081 26333 12115 26367
rect 12265 26333 12299 26367
rect 12449 26333 12483 26367
rect 14284 26333 14318 26367
rect 14473 26333 14507 26367
rect 14656 26333 14690 26367
rect 14749 26333 14783 26367
rect 15572 26333 15606 26367
rect 15889 26333 15923 26367
rect 16037 26333 16071 26367
rect 16129 26333 16163 26367
rect 16277 26333 16311 26367
rect 16405 26333 16439 26367
rect 16594 26333 16628 26367
rect 17253 26333 17287 26367
rect 17785 26333 17819 26367
rect 18153 26333 18187 26367
rect 18705 26333 18739 26367
rect 18981 26333 19015 26367
rect 20821 26333 20855 26367
rect 21005 26333 21039 26367
rect 21281 26333 21315 26367
rect 22201 26333 22235 26367
rect 22385 26333 22419 26367
rect 23121 26333 23155 26367
rect 23581 26333 23615 26367
rect 23673 26333 23707 26367
rect 24593 26333 24627 26367
rect 24685 26333 24719 26367
rect 25145 26333 25179 26367
rect 25237 26333 25271 26367
rect 26893 26333 26927 26367
rect 26985 26333 27019 26367
rect 27813 26333 27847 26367
rect 27905 26333 27939 26367
rect 27997 26333 28031 26367
rect 28273 26333 28307 26367
rect 28457 26333 28491 26367
rect 28825 26333 28859 26367
rect 29929 26333 29963 26367
rect 31125 26333 31159 26367
rect 31309 26333 31343 26367
rect 31401 26333 31435 26367
rect 31585 26333 31619 26367
rect 31677 26333 31711 26367
rect 31861 26333 31895 26367
rect 32321 26333 32355 26367
rect 32505 26333 32539 26367
rect 32597 26333 32631 26367
rect 34345 26333 34379 26367
rect 34529 26333 34563 26367
rect 34897 26333 34931 26367
rect 35265 26333 35299 26367
rect 35357 26333 35391 26367
rect 37933 26333 37967 26367
rect 40233 26333 40267 26367
rect 3065 26265 3099 26299
rect 3801 26265 3835 26299
rect 5549 26265 5583 26299
rect 5641 26265 5675 26299
rect 6285 26265 6319 26299
rect 6377 26265 6411 26299
rect 7113 26265 7147 26299
rect 8309 26265 8343 26299
rect 9137 26265 9171 26299
rect 11713 26265 11747 26299
rect 14381 26265 14415 26299
rect 15669 26265 15703 26299
rect 15761 26265 15795 26299
rect 16497 26265 16531 26299
rect 16865 26265 16899 26299
rect 17049 26265 17083 26299
rect 17141 26265 17175 26299
rect 17877 26265 17911 26299
rect 17969 26265 18003 26299
rect 19073 26265 19107 26299
rect 23029 26265 23063 26299
rect 24869 26265 24903 26299
rect 24961 26265 24995 26299
rect 25681 26265 25715 26299
rect 25881 26265 25915 26299
rect 31217 26265 31251 26299
rect 32781 26265 32815 26299
rect 35633 26265 35667 26299
rect 38393 26265 38427 26299
rect 2697 26197 2731 26231
rect 11805 26197 11839 26231
rect 15393 26197 15427 26231
rect 16773 26197 16807 26231
rect 17601 26197 17635 26231
rect 22845 26197 22879 26231
rect 23305 26197 23339 26231
rect 31861 26197 31895 26231
rect 35725 26197 35759 26231
rect 3341 25993 3375 26027
rect 5457 25993 5491 26027
rect 7757 25993 7791 26027
rect 10149 25993 10183 26027
rect 18429 25993 18463 26027
rect 26065 25993 26099 26027
rect 28365 25993 28399 26027
rect 29469 25993 29503 26027
rect 30573 25993 30607 26027
rect 38117 25993 38151 26027
rect 1869 25925 1903 25959
rect 6653 25925 6687 25959
rect 7389 25925 7423 25959
rect 10333 25925 10367 25959
rect 12633 25925 12667 25959
rect 19257 25925 19291 25959
rect 29193 25925 29227 25959
rect 30389 25925 30423 25959
rect 31217 25925 31251 25959
rect 34779 25925 34813 25959
rect 34989 25925 35023 25959
rect 3709 25857 3743 25891
rect 6101 25857 6135 25891
rect 6377 25857 6411 25891
rect 6525 25857 6559 25891
rect 6745 25857 6779 25891
rect 6883 25857 6917 25891
rect 7113 25857 7147 25891
rect 7206 25857 7240 25891
rect 7481 25857 7515 25891
rect 7619 25857 7653 25891
rect 10057 25857 10091 25891
rect 11529 25857 11563 25891
rect 11713 25857 11747 25891
rect 11897 25857 11931 25891
rect 12357 25857 12391 25891
rect 12449 25857 12483 25891
rect 13369 25857 13403 25891
rect 13553 25857 13587 25891
rect 13645 25857 13679 25891
rect 13829 25857 13863 25891
rect 13921 25857 13955 25891
rect 14013 25857 14047 25891
rect 14473 25857 14507 25891
rect 14565 25857 14599 25891
rect 14749 25857 14783 25891
rect 18153 25857 18187 25891
rect 18429 25857 18463 25891
rect 19073 25857 19107 25891
rect 25973 25857 26007 25891
rect 26157 25857 26191 25891
rect 28457 25857 28491 25891
rect 29009 25857 29043 25891
rect 29285 25857 29319 25891
rect 29377 25857 29411 25891
rect 29837 25857 29871 25891
rect 30205 25857 30239 25891
rect 30941 25857 30975 25891
rect 31677 25857 31711 25891
rect 32505 25857 32539 25891
rect 33885 25857 33919 25891
rect 34069 25857 34103 25891
rect 34161 25857 34195 25891
rect 34437 25857 34471 25891
rect 34621 25857 34655 25891
rect 34897 25857 34931 25891
rect 35081 25857 35115 25891
rect 38000 25857 38034 25891
rect 38485 25857 38519 25891
rect 1593 25789 1627 25823
rect 3985 25789 4019 25823
rect 14289 25789 14323 25823
rect 14381 25789 14415 25823
rect 15485 25789 15519 25823
rect 15945 25789 15979 25823
rect 31309 25789 31343 25823
rect 35449 25789 35483 25823
rect 38209 25789 38243 25823
rect 14197 25721 14231 25755
rect 15577 25721 15611 25755
rect 18337 25721 18371 25755
rect 34437 25721 34471 25755
rect 35725 25721 35759 25755
rect 5549 25653 5583 25687
rect 7021 25653 7055 25687
rect 10333 25653 10367 25687
rect 12633 25653 12667 25687
rect 13553 25653 13587 25687
rect 18981 25653 19015 25687
rect 29009 25653 29043 25687
rect 30757 25653 30791 25687
rect 32321 25653 32355 25687
rect 34069 25653 34103 25687
rect 35265 25653 35299 25687
rect 35909 25653 35943 25687
rect 37841 25653 37875 25687
rect 4537 25449 4571 25483
rect 6377 25449 6411 25483
rect 7297 25449 7331 25483
rect 11253 25449 11287 25483
rect 15485 25449 15519 25483
rect 16221 25449 16255 25483
rect 20361 25449 20395 25483
rect 23765 25449 23799 25483
rect 24869 25449 24903 25483
rect 30389 25449 30423 25483
rect 31861 25449 31895 25483
rect 32597 25449 32631 25483
rect 38025 25449 38059 25483
rect 25973 25381 26007 25415
rect 30573 25381 30607 25415
rect 1593 25313 1627 25347
rect 4997 25313 5031 25347
rect 5181 25313 5215 25347
rect 8493 25313 8527 25347
rect 18705 25313 18739 25347
rect 23305 25313 23339 25347
rect 23489 25313 23523 25347
rect 25237 25313 25271 25347
rect 25329 25313 25363 25347
rect 26525 25313 26559 25347
rect 30665 25313 30699 25347
rect 30941 25313 30975 25347
rect 32965 25313 32999 25347
rect 36001 25313 36035 25347
rect 38117 25313 38151 25347
rect 4445 25245 4479 25279
rect 4905 25245 4939 25279
rect 5733 25245 5767 25279
rect 6101 25245 6135 25279
rect 6561 25245 6595 25279
rect 6653 25245 6687 25279
rect 6929 25245 6963 25279
rect 7021 25245 7055 25279
rect 9505 25245 9539 25279
rect 16497 25245 16531 25279
rect 18521 25245 18555 25279
rect 20269 25245 20303 25279
rect 20453 25245 20487 25279
rect 23397 25245 23431 25279
rect 23581 25245 23615 25279
rect 25053 25245 25087 25279
rect 25605 25245 25639 25279
rect 25881 25245 25915 25279
rect 26157 25245 26191 25279
rect 26249 25245 26283 25279
rect 26341 25245 26375 25279
rect 26709 25245 26743 25279
rect 26801 25245 26835 25279
rect 31677 25245 31711 25279
rect 31861 25245 31895 25279
rect 31953 25245 31987 25279
rect 32137 25245 32171 25279
rect 33057 25245 33091 25279
rect 33149 25245 33183 25279
rect 33333 25245 33367 25279
rect 33425 25245 33459 25279
rect 33701 25245 33735 25279
rect 35541 25245 35575 25279
rect 35633 25245 35667 25279
rect 36093 25245 36127 25279
rect 36241 25245 36275 25279
rect 36369 25245 36403 25279
rect 36461 25245 36495 25279
rect 36599 25245 36633 25279
rect 38025 25245 38059 25279
rect 30435 25211 30469 25245
rect 1869 25177 1903 25211
rect 5917 25177 5951 25211
rect 6009 25177 6043 25211
rect 6745 25177 6779 25211
rect 7205 25177 7239 25211
rect 8953 25177 8987 25211
rect 11437 25177 11471 25211
rect 15669 25177 15703 25211
rect 16221 25177 16255 25211
rect 25421 25177 25455 25211
rect 26525 25177 26559 25211
rect 30205 25177 30239 25211
rect 35909 25177 35943 25211
rect 3341 25109 3375 25143
rect 3801 25109 3835 25143
rect 6285 25109 6319 25143
rect 7941 25109 7975 25143
rect 8309 25109 8343 25143
rect 8401 25109 8435 25143
rect 11069 25109 11103 25143
rect 11237 25109 11271 25143
rect 15301 25109 15335 25143
rect 15469 25109 15503 25143
rect 16405 25109 16439 25143
rect 18337 25109 18371 25143
rect 25789 25109 25823 25143
rect 32045 25109 32079 25143
rect 32413 25109 32447 25143
rect 32597 25109 32631 25143
rect 33609 25109 33643 25143
rect 33885 25109 33919 25143
rect 35357 25109 35391 25143
rect 35817 25109 35851 25143
rect 36737 25109 36771 25143
rect 38393 25109 38427 25143
rect 2605 24905 2639 24939
rect 2973 24905 3007 24939
rect 9045 24905 9079 24939
rect 11069 24905 11103 24939
rect 12173 24905 12207 24939
rect 20361 24905 20395 24939
rect 22017 24905 22051 24939
rect 24777 24905 24811 24939
rect 25145 24905 25179 24939
rect 25989 24905 26023 24939
rect 40049 24905 40083 24939
rect 3065 24837 3099 24871
rect 7573 24837 7607 24871
rect 9413 24837 9447 24871
rect 10793 24837 10827 24871
rect 11897 24837 11931 24871
rect 17693 24837 17727 24871
rect 19993 24837 20027 24871
rect 24409 24837 24443 24871
rect 25605 24837 25639 24871
rect 25789 24837 25823 24871
rect 26433 24837 26467 24871
rect 38853 24837 38887 24871
rect 5457 24769 5491 24803
rect 5641 24769 5675 24803
rect 5733 24769 5767 24803
rect 5825 24769 5859 24803
rect 9316 24769 9350 24803
rect 9505 24769 9539 24803
rect 9688 24769 9722 24803
rect 9781 24769 9815 24803
rect 10517 24769 10551 24803
rect 10701 24769 10735 24803
rect 10885 24769 10919 24803
rect 11529 24769 11563 24803
rect 11622 24769 11656 24803
rect 11805 24769 11839 24803
rect 11994 24769 12028 24803
rect 12265 24769 12299 24803
rect 12449 24769 12483 24803
rect 14473 24769 14507 24803
rect 14565 24769 14599 24803
rect 14749 24769 14783 24803
rect 14841 24769 14875 24803
rect 14933 24769 14967 24803
rect 15301 24769 15335 24803
rect 15485 24769 15519 24803
rect 16037 24769 16071 24803
rect 16221 24769 16255 24803
rect 16497 24769 16531 24803
rect 16956 24775 16990 24809
rect 39083 24803 39117 24837
rect 17049 24769 17083 24803
rect 17141 24769 17175 24803
rect 17325 24769 17359 24803
rect 17417 24769 17451 24803
rect 19073 24769 19107 24803
rect 19257 24769 19291 24803
rect 19809 24769 19843 24803
rect 20085 24769 20119 24803
rect 20177 24769 20211 24803
rect 20729 24769 20763 24803
rect 21097 24769 21131 24803
rect 21281 24769 21315 24803
rect 21557 24769 21591 24803
rect 21958 24769 21992 24803
rect 22477 24769 22511 24803
rect 24317 24769 24351 24803
rect 24501 24769 24535 24803
rect 24593 24769 24627 24803
rect 24777 24769 24811 24803
rect 24869 24769 24903 24803
rect 27261 24769 27295 24803
rect 27721 24769 27755 24803
rect 27905 24769 27939 24803
rect 28181 24769 28215 24803
rect 28365 24769 28399 24803
rect 28549 24769 28583 24803
rect 30481 24769 30515 24803
rect 31309 24769 31343 24803
rect 31493 24769 31527 24803
rect 31585 24769 31619 24803
rect 31677 24769 31711 24803
rect 35173 24769 35207 24803
rect 35265 24769 35299 24803
rect 35449 24769 35483 24803
rect 35633 24769 35667 24803
rect 37473 24769 37507 24803
rect 37749 24769 37783 24803
rect 38393 24769 38427 24803
rect 38577 24769 38611 24803
rect 40233 24769 40267 24803
rect 3249 24701 3283 24735
rect 3985 24701 4019 24735
rect 7297 24701 7331 24735
rect 15025 24701 15059 24735
rect 15669 24701 15703 24735
rect 16405 24701 16439 24735
rect 17509 24701 17543 24735
rect 18981 24701 19015 24735
rect 21373 24701 21407 24735
rect 25053 24701 25087 24735
rect 26985 24701 27019 24735
rect 27077 24701 27111 24735
rect 30297 24701 30331 24735
rect 37657 24701 37691 24735
rect 38761 24701 38795 24735
rect 16681 24633 16715 24667
rect 25605 24633 25639 24667
rect 26157 24633 26191 24667
rect 26249 24633 26283 24667
rect 26801 24633 26835 24667
rect 27445 24633 27479 24667
rect 30665 24633 30699 24667
rect 3433 24565 3467 24599
rect 6009 24565 6043 24599
rect 9137 24565 9171 24599
rect 12541 24565 12575 24599
rect 17417 24565 17451 24599
rect 21833 24565 21867 24599
rect 22385 24565 22419 24599
rect 25973 24565 26007 24599
rect 26433 24565 26467 24599
rect 27537 24565 27571 24599
rect 27997 24565 28031 24599
rect 28181 24565 28215 24599
rect 28733 24565 28767 24599
rect 31861 24565 31895 24599
rect 37289 24565 37323 24599
rect 37473 24565 37507 24599
rect 39037 24565 39071 24599
rect 39221 24565 39255 24599
rect 3157 24361 3191 24395
rect 6929 24361 6963 24395
rect 9597 24361 9631 24395
rect 14749 24361 14783 24395
rect 17785 24361 17819 24395
rect 19993 24361 20027 24395
rect 20361 24361 20395 24395
rect 23857 24361 23891 24395
rect 24133 24361 24167 24395
rect 26157 24361 26191 24395
rect 26617 24361 26651 24395
rect 27261 24361 27295 24395
rect 28825 24361 28859 24395
rect 37933 24361 37967 24395
rect 40049 24361 40083 24395
rect 15117 24293 15151 24327
rect 15301 24293 15335 24327
rect 15761 24293 15795 24327
rect 20453 24293 20487 24327
rect 23673 24293 23707 24327
rect 24961 24293 24995 24327
rect 29285 24293 29319 24327
rect 1409 24225 1443 24259
rect 3801 24225 3835 24259
rect 5549 24225 5583 24259
rect 6193 24225 6227 24259
rect 11345 24225 11379 24259
rect 15577 24225 15611 24259
rect 16589 24225 16623 24259
rect 18521 24225 18555 24259
rect 20269 24225 20303 24259
rect 24501 24225 24535 24259
rect 6377 24157 6411 24191
rect 6561 24157 6595 24191
rect 6653 24157 6687 24191
rect 6745 24157 6779 24191
rect 8033 24157 8067 24191
rect 8126 24157 8160 24191
rect 8309 24157 8343 24191
rect 8517 24157 8551 24191
rect 8941 24157 8975 24191
rect 9046 24157 9080 24191
rect 9229 24157 9263 24191
rect 9418 24157 9452 24191
rect 10977 24157 11011 24191
rect 11161 24157 11195 24191
rect 14105 24157 14139 24191
rect 14381 24157 14415 24191
rect 14472 24157 14506 24191
rect 14565 24157 14599 24191
rect 15761 24157 15795 24191
rect 16037 24157 16071 24191
rect 16405 24157 16439 24191
rect 17969 24157 18003 24191
rect 18153 24157 18187 24191
rect 18245 24157 18279 24191
rect 19625 24157 19659 24191
rect 20545 24157 20579 24191
rect 23029 24157 23063 24191
rect 23177 24157 23211 24191
rect 23494 24157 23528 24191
rect 23765 24157 23799 24191
rect 23949 24157 23983 24191
rect 25237 24157 25271 24191
rect 25697 24157 25731 24191
rect 25881 24157 25915 24191
rect 26157 24157 26191 24191
rect 27445 24157 27479 24191
rect 27537 24157 27571 24191
rect 27721 24157 27755 24191
rect 27813 24157 27847 24191
rect 28089 24157 28123 24191
rect 28182 24157 28216 24191
rect 28457 24157 28491 24191
rect 28554 24157 28588 24191
rect 29009 24157 29043 24191
rect 29101 24157 29135 24191
rect 38117 24157 38151 24191
rect 38301 24157 38335 24191
rect 38485 24157 38519 24191
rect 38577 24157 38611 24191
rect 39681 24157 39715 24191
rect 40233 24157 40267 24191
rect 1685 24089 1719 24123
rect 4077 24089 4111 24123
rect 8401 24089 8435 24123
rect 9321 24089 9355 24123
rect 14263 24089 14297 24123
rect 16221 24089 16255 24123
rect 18705 24089 18739 24123
rect 18889 24089 18923 24123
rect 23305 24089 23339 24123
rect 23397 24089 23431 24123
rect 25973 24089 26007 24123
rect 26249 24089 26283 24123
rect 26433 24089 26467 24123
rect 28365 24089 28399 24123
rect 28825 24089 28859 24123
rect 38209 24089 38243 24123
rect 5641 24021 5675 24055
rect 8677 24021 8711 24055
rect 19993 24021 20027 24055
rect 20177 24021 20211 24055
rect 28733 24021 28767 24055
rect 39497 24021 39531 24055
rect 2513 23817 2547 23851
rect 2881 23817 2915 23851
rect 4997 23817 5031 23851
rect 7849 23817 7883 23851
rect 18613 23817 18647 23851
rect 19165 23817 19199 23851
rect 20085 23817 20119 23851
rect 20453 23817 20487 23851
rect 23765 23817 23799 23851
rect 27905 23817 27939 23851
rect 29101 23817 29135 23851
rect 31125 23817 31159 23851
rect 33517 23817 33551 23851
rect 34621 23817 34655 23851
rect 3709 23749 3743 23783
rect 4537 23749 4571 23783
rect 5917 23749 5951 23783
rect 6653 23749 6687 23783
rect 8125 23749 8159 23783
rect 11345 23749 11379 23783
rect 19349 23749 19383 23783
rect 20621 23749 20655 23783
rect 20821 23749 20855 23783
rect 23213 23749 23247 23783
rect 23305 23749 23339 23783
rect 27169 23749 27203 23783
rect 29653 23749 29687 23783
rect 34713 23749 34747 23783
rect 36369 23749 36403 23783
rect 38485 23749 38519 23783
rect 2973 23681 3007 23715
rect 5825 23681 5859 23715
rect 6009 23681 6043 23715
rect 6193 23681 6227 23715
rect 6561 23681 6595 23715
rect 6745 23681 6779 23715
rect 6929 23681 6963 23715
rect 7987 23681 8021 23715
rect 8217 23681 8251 23715
rect 8400 23681 8434 23715
rect 8486 23681 8520 23715
rect 8769 23681 8803 23715
rect 8861 23681 8895 23715
rect 8953 23681 8987 23715
rect 9137 23681 9171 23715
rect 10977 23681 11011 23715
rect 15025 23681 15059 23715
rect 15209 23681 15243 23715
rect 15485 23681 15519 23715
rect 15761 23681 15795 23715
rect 15945 23681 15979 23715
rect 17325 23681 17359 23715
rect 18153 23681 18187 23715
rect 18797 23681 18831 23715
rect 19533 23681 19567 23715
rect 19901 23681 19935 23715
rect 20177 23681 20211 23715
rect 22569 23681 22603 23715
rect 22753 23681 22787 23715
rect 22937 23681 22971 23715
rect 23029 23681 23063 23715
rect 23397 23681 23431 23715
rect 23949 23681 23983 23715
rect 26985 23681 27019 23715
rect 28089 23681 28123 23715
rect 28254 23681 28288 23715
rect 28365 23681 28399 23715
rect 28457 23681 28491 23715
rect 28549 23681 28583 23715
rect 28825 23681 28859 23715
rect 28917 23681 28951 23715
rect 31033 23681 31067 23715
rect 31217 23681 31251 23715
rect 33057 23681 33091 23715
rect 33333 23681 33367 23715
rect 33977 23681 34011 23715
rect 34125 23681 34159 23715
rect 34253 23681 34287 23715
rect 34345 23681 34379 23715
rect 34442 23681 34476 23715
rect 34897 23681 34931 23715
rect 36553 23681 36587 23715
rect 3157 23613 3191 23647
rect 5089 23613 5123 23647
rect 5273 23613 5307 23647
rect 10865 23613 10899 23647
rect 11253 23613 11287 23647
rect 12173 23613 12207 23647
rect 12449 23613 12483 23647
rect 14565 23613 14599 23647
rect 17049 23613 17083 23647
rect 17601 23613 17635 23647
rect 18337 23613 18371 23647
rect 18981 23613 19015 23647
rect 19073 23613 19107 23647
rect 24133 23613 24167 23647
rect 24225 23613 24259 23647
rect 29193 23613 29227 23647
rect 33241 23613 33275 23647
rect 36737 23613 36771 23647
rect 38209 23613 38243 23647
rect 40233 23613 40267 23647
rect 4629 23545 4663 23579
rect 10701 23545 10735 23579
rect 15393 23545 15427 23579
rect 23581 23545 23615 23579
rect 27353 23545 27387 23579
rect 29285 23545 29319 23579
rect 5641 23477 5675 23511
rect 6377 23477 6411 23511
rect 8585 23477 8619 23511
rect 13921 23477 13955 23511
rect 14013 23477 14047 23511
rect 15577 23477 15611 23511
rect 15945 23477 15979 23511
rect 19901 23477 19935 23511
rect 20637 23477 20671 23511
rect 28641 23477 28675 23511
rect 33057 23477 33091 23511
rect 35081 23477 35115 23511
rect 4445 23273 4479 23307
rect 9045 23273 9079 23307
rect 9873 23273 9907 23307
rect 10333 23273 10367 23307
rect 11529 23273 11563 23307
rect 12173 23273 12207 23307
rect 12633 23273 12667 23307
rect 16589 23273 16623 23307
rect 16773 23273 16807 23307
rect 18061 23273 18095 23307
rect 18153 23273 18187 23307
rect 29101 23273 29135 23307
rect 38301 23273 38335 23307
rect 38669 23273 38703 23307
rect 39497 23273 39531 23307
rect 5273 23205 5307 23239
rect 5549 23205 5583 23239
rect 5641 23205 5675 23239
rect 5917 23205 5951 23239
rect 14749 23205 14783 23239
rect 31769 23205 31803 23239
rect 3617 23137 3651 23171
rect 10241 23137 10275 23171
rect 11621 23137 11655 23171
rect 13093 23137 13127 23171
rect 13277 23137 13311 23171
rect 17969 23137 18003 23171
rect 30481 23137 30515 23171
rect 33057 23137 33091 23171
rect 33149 23137 33183 23171
rect 33517 23137 33551 23171
rect 2421 23069 2455 23103
rect 4721 23069 4755 23103
rect 4997 23069 5031 23103
rect 5089 23069 5123 23103
rect 5457 23069 5491 23103
rect 5733 23069 5767 23103
rect 6101 23069 6135 23103
rect 6377 23069 6411 23103
rect 6745 23069 6779 23103
rect 7481 23069 7515 23103
rect 8953 23069 8987 23103
rect 9137 23069 9171 23103
rect 10517 23069 10551 23103
rect 10609 23069 10643 23103
rect 11158 23069 11192 23103
rect 11897 23069 11931 23103
rect 11989 23069 12023 23103
rect 12265 23069 12299 23103
rect 13001 23069 13035 23103
rect 14473 23069 14507 23103
rect 16865 23069 16899 23103
rect 17141 23069 17175 23103
rect 18061 23069 18095 23103
rect 18337 23069 18371 23103
rect 18429 23069 18463 23103
rect 18797 23069 18831 23103
rect 22293 23069 22327 23103
rect 22477 23069 22511 23103
rect 30113 23069 30147 23103
rect 30297 23069 30331 23103
rect 31217 23069 31251 23103
rect 31493 23069 31527 23103
rect 31585 23069 31619 23103
rect 36093 23069 36127 23103
rect 36186 23069 36220 23103
rect 36461 23069 36495 23103
rect 36558 23069 36592 23103
rect 38485 23069 38519 23103
rect 38577 23069 38611 23103
rect 39589 23069 39623 23103
rect 4537 23001 4571 23035
rect 4905 23001 4939 23035
rect 7205 23001 7239 23035
rect 9781 23001 9815 23035
rect 11713 23001 11747 23035
rect 13645 23001 13679 23035
rect 13829 23001 13863 23035
rect 14197 23001 14231 23035
rect 29285 23001 29319 23035
rect 31401 23001 31435 23035
rect 33425 23001 33459 23035
rect 36369 23001 36403 23035
rect 38761 23001 38795 23035
rect 2973 22933 3007 22967
rect 10793 22933 10827 22967
rect 10977 22933 11011 22967
rect 11161 22933 11195 22967
rect 14289 22933 14323 22967
rect 17693 22933 17727 22967
rect 18521 22933 18555 22967
rect 18705 22933 18739 22967
rect 22293 22933 22327 22967
rect 28917 22933 28951 22967
rect 29085 22933 29119 22967
rect 32873 22933 32907 22967
rect 33333 22933 33367 22967
rect 36737 22933 36771 22967
rect 2605 22729 2639 22763
rect 2697 22729 2731 22763
rect 6193 22729 6227 22763
rect 11897 22729 11931 22763
rect 21281 22729 21315 22763
rect 25421 22729 25455 22763
rect 25697 22729 25731 22763
rect 27537 22729 27571 22763
rect 29653 22729 29687 22763
rect 30665 22729 30699 22763
rect 32689 22729 32723 22763
rect 5825 22661 5859 22695
rect 14197 22661 14231 22695
rect 21465 22661 21499 22695
rect 28181 22661 28215 22695
rect 29285 22661 29319 22695
rect 31585 22661 31619 22695
rect 36093 22661 36127 22695
rect 3065 22593 3099 22627
rect 5641 22593 5675 22627
rect 5917 22593 5951 22627
rect 6009 22593 6043 22627
rect 8493 22593 8527 22627
rect 8677 22593 8711 22627
rect 8769 22593 8803 22627
rect 10793 22593 10827 22627
rect 10885 22593 10919 22627
rect 11161 22593 11195 22627
rect 11989 22593 12023 22627
rect 12449 22593 12483 22627
rect 14013 22593 14047 22627
rect 20361 22593 20395 22627
rect 20453 22593 20487 22627
rect 20637 22593 20671 22627
rect 20729 22593 20763 22627
rect 24041 22593 24075 22627
rect 24133 22593 24167 22627
rect 24317 22593 24351 22627
rect 24409 22593 24443 22627
rect 25580 22593 25614 22627
rect 26157 22593 26191 22627
rect 26617 22593 26651 22627
rect 26709 22593 26743 22627
rect 27721 22593 27755 22627
rect 28457 22593 28491 22627
rect 28912 22593 28946 22627
rect 29009 22593 29043 22627
rect 29101 22593 29135 22627
rect 29837 22593 29871 22627
rect 29929 22593 29963 22627
rect 30297 22593 30331 22627
rect 30389 22593 30423 22627
rect 30849 22593 30883 22627
rect 31401 22593 31435 22627
rect 31677 22593 31711 22627
rect 31769 22593 31803 22627
rect 32137 22593 32171 22627
rect 32321 22593 32355 22627
rect 32413 22593 32447 22627
rect 32505 22593 32539 22627
rect 32873 22593 32907 22627
rect 33057 22593 33091 22627
rect 35817 22593 35851 22627
rect 35910 22593 35944 22627
rect 36185 22593 36219 22627
rect 36323 22593 36357 22627
rect 38025 22593 38059 22627
rect 2789 22525 2823 22559
rect 3341 22525 3375 22559
rect 4813 22525 4847 22559
rect 5457 22525 5491 22559
rect 9505 22525 9539 22559
rect 11713 22525 11747 22559
rect 12541 22525 12575 22559
rect 25789 22525 25823 22559
rect 26065 22525 26099 22559
rect 26433 22525 26467 22559
rect 27905 22525 27939 22559
rect 28273 22525 28307 22559
rect 28733 22525 28767 22559
rect 29193 22525 29227 22559
rect 32965 22525 32999 22559
rect 33149 22525 33183 22559
rect 38117 22525 38151 22559
rect 4905 22457 4939 22491
rect 8585 22457 8619 22491
rect 10609 22457 10643 22491
rect 26341 22457 26375 22491
rect 28641 22457 28675 22491
rect 31953 22457 31987 22491
rect 33333 22457 33367 22491
rect 2237 22389 2271 22423
rect 8953 22389 8987 22423
rect 10057 22389 10091 22423
rect 11069 22389 11103 22423
rect 12357 22389 12391 22423
rect 13829 22389 13863 22423
rect 20913 22389 20947 22423
rect 21097 22389 21131 22423
rect 21281 22389 21315 22423
rect 24501 22389 24535 22423
rect 26525 22389 26559 22423
rect 28089 22389 28123 22423
rect 30113 22389 30147 22423
rect 36461 22389 36495 22423
rect 38025 22389 38059 22423
rect 38393 22389 38427 22423
rect 1764 22185 1798 22219
rect 3249 22185 3283 22219
rect 8677 22185 8711 22219
rect 19717 22185 19751 22219
rect 20085 22185 20119 22219
rect 20177 22185 20211 22219
rect 25329 22185 25363 22219
rect 26065 22185 26099 22219
rect 27353 22185 27387 22219
rect 31953 22185 31987 22219
rect 38209 22185 38243 22219
rect 38301 22185 38335 22219
rect 38669 22185 38703 22219
rect 7297 22117 7331 22151
rect 11529 22117 11563 22151
rect 14381 22117 14415 22151
rect 19993 22117 20027 22151
rect 22109 22117 22143 22151
rect 38393 22117 38427 22151
rect 38761 22117 38795 22151
rect 10701 22049 10735 22083
rect 12449 22049 12483 22083
rect 12909 22049 12943 22083
rect 13829 22049 13863 22083
rect 21005 22049 21039 22083
rect 21465 22049 21499 22083
rect 23765 22049 23799 22083
rect 24777 22049 24811 22083
rect 25053 22049 25087 22083
rect 25973 22049 26007 22083
rect 26617 22049 26651 22083
rect 30297 22049 30331 22083
rect 1501 21981 1535 22015
rect 4353 21981 4387 22015
rect 5917 21981 5951 22015
rect 6193 21981 6227 22015
rect 6285 21981 6319 22015
rect 6377 21981 6411 22015
rect 6469 21981 6503 22015
rect 7021 21981 7055 22015
rect 7205 21981 7239 22015
rect 7389 21981 7423 22015
rect 8125 21981 8159 22015
rect 8493 21981 8527 22015
rect 10793 21981 10827 22015
rect 10885 21981 10919 22015
rect 11069 21981 11103 22015
rect 11161 21981 11195 22015
rect 11345 21981 11379 22015
rect 11437 21981 11471 22015
rect 11621 21981 11655 22015
rect 12541 21981 12575 22015
rect 12633 21981 12667 22015
rect 12725 21981 12759 22015
rect 13001 21981 13035 22015
rect 13093 21981 13127 22015
rect 13461 21981 13495 22015
rect 13737 21981 13771 22015
rect 13921 21981 13955 22015
rect 14381 21981 14415 22015
rect 14749 21981 14783 22015
rect 15117 21981 15151 22015
rect 17049 21981 17083 22015
rect 17142 21981 17176 22015
rect 17325 21981 17359 22015
rect 17555 21981 17589 22015
rect 17969 21981 18003 22015
rect 18245 21981 18279 22015
rect 20269 21981 20303 22015
rect 20453 21981 20487 22015
rect 20821 21981 20855 22015
rect 21189 21981 21223 22015
rect 21281 21981 21315 22015
rect 21373 21981 21407 22015
rect 22477 21981 22511 22015
rect 22937 21981 22971 22015
rect 23397 21981 23431 22015
rect 24041 21981 24075 22015
rect 24869 21981 24903 22015
rect 26065 21981 26099 22015
rect 26801 21981 26835 22015
rect 27077 21981 27111 22015
rect 27445 21981 27479 22015
rect 27537 21981 27571 22015
rect 30113 21981 30147 22015
rect 30573 21981 30607 22015
rect 30757 21981 30791 22015
rect 37933 21981 37967 22015
rect 38945 21981 38979 22015
rect 39129 21981 39163 22015
rect 39313 21981 39347 22015
rect 39405 21981 39439 22015
rect 5181 21913 5215 21947
rect 8309 21913 8343 21947
rect 8401 21913 8435 21947
rect 10425 21913 10459 21947
rect 13277 21913 13311 21947
rect 13369 21913 13403 21947
rect 17417 21913 17451 21947
rect 20545 21913 20579 21947
rect 25145 21913 25179 21947
rect 25350 21913 25384 21947
rect 25605 21913 25639 21947
rect 31861 21913 31895 21947
rect 39037 21913 39071 21947
rect 5365 21845 5399 21879
rect 6653 21845 6687 21879
rect 8953 21845 8987 21879
rect 13645 21845 13679 21879
rect 17693 21845 17727 21879
rect 17785 21845 17819 21879
rect 18153 21845 18187 21879
rect 20643 21845 20677 21879
rect 20729 21845 20763 21879
rect 24409 21845 24443 21879
rect 25513 21845 25547 21879
rect 26249 21845 26283 21879
rect 26985 21845 27019 21879
rect 27169 21845 27203 21879
rect 29929 21845 29963 21879
rect 30389 21845 30423 21879
rect 38025 21845 38059 21879
rect 3985 21641 4019 21675
rect 4353 21641 4387 21675
rect 5181 21641 5215 21675
rect 6193 21641 6227 21675
rect 8585 21641 8619 21675
rect 9781 21641 9815 21675
rect 10149 21641 10183 21675
rect 14105 21641 14139 21675
rect 20821 21641 20855 21675
rect 23863 21641 23897 21675
rect 33701 21641 33735 21675
rect 34069 21641 34103 21675
rect 3433 21573 3467 21607
rect 13185 21573 13219 21607
rect 16773 21573 16807 21607
rect 21097 21573 21131 21607
rect 23949 21573 23983 21607
rect 27537 21573 27571 21607
rect 27629 21573 27663 21607
rect 28089 21573 28123 21607
rect 34713 21573 34747 21607
rect 35587 21573 35621 21607
rect 35817 21573 35851 21607
rect 36369 21573 36403 21607
rect 3617 21505 3651 21539
rect 3801 21505 3835 21539
rect 3893 21505 3927 21539
rect 4445 21505 4479 21539
rect 5733 21505 5767 21539
rect 5917 21505 5951 21539
rect 6009 21505 6043 21539
rect 9229 21505 9263 21539
rect 12812 21505 12846 21539
rect 12909 21505 12943 21539
rect 13001 21505 13035 21539
rect 14289 21505 14323 21539
rect 14473 21505 14507 21539
rect 16681 21505 16715 21539
rect 16865 21505 16899 21539
rect 16957 21505 16991 21539
rect 17141 21505 17175 21539
rect 20959 21505 20993 21539
rect 21189 21505 21223 21539
rect 21372 21505 21406 21539
rect 21465 21505 21499 21539
rect 23765 21505 23799 21539
rect 24041 21505 24075 21539
rect 27261 21505 27295 21539
rect 27354 21505 27388 21539
rect 27726 21505 27760 21539
rect 27997 21505 28031 21539
rect 28273 21505 28307 21539
rect 31861 21505 31895 21539
rect 33517 21505 33551 21539
rect 33885 21505 33919 21539
rect 34529 21505 34563 21539
rect 34805 21505 34839 21539
rect 34897 21505 34931 21539
rect 35449 21505 35483 21539
rect 35725 21505 35759 21539
rect 35909 21505 35943 21539
rect 36185 21505 36219 21539
rect 36461 21505 36495 21539
rect 36553 21505 36587 21539
rect 1501 21437 1535 21471
rect 1777 21437 1811 21471
rect 4629 21437 4663 21471
rect 5273 21437 5307 21471
rect 5365 21437 5399 21471
rect 6837 21437 6871 21471
rect 7113 21437 7147 21471
rect 9597 21437 9631 21471
rect 9689 21437 9723 21471
rect 14565 21437 14599 21471
rect 28365 21437 28399 21471
rect 4813 21369 4847 21403
rect 5825 21369 5859 21403
rect 13185 21369 13219 21403
rect 3249 21301 3283 21335
rect 8677 21301 8711 21335
rect 17049 21301 17083 21335
rect 27905 21301 27939 21335
rect 28365 21301 28399 21335
rect 31677 21301 31711 21335
rect 35081 21301 35115 21335
rect 36093 21301 36127 21335
rect 36737 21301 36771 21335
rect 6653 21097 6687 21131
rect 7665 21097 7699 21131
rect 10885 21097 10919 21131
rect 23397 21097 23431 21131
rect 23581 21097 23615 21131
rect 36553 21097 36587 21131
rect 37013 21097 37047 21131
rect 6561 21029 6595 21063
rect 17325 21029 17359 21063
rect 18705 21029 18739 21063
rect 5089 20961 5123 20995
rect 8309 20961 8343 20995
rect 10977 20961 11011 20995
rect 12725 20961 12759 20995
rect 13369 20961 13403 20995
rect 19809 20961 19843 20995
rect 23765 20961 23799 20995
rect 32505 20961 32539 20995
rect 36737 20961 36771 20995
rect 1869 20893 1903 20927
rect 4905 20893 4939 20927
rect 5917 20893 5951 20927
rect 6009 20893 6043 20927
rect 6101 20893 6135 20927
rect 6212 20893 6246 20927
rect 6377 20893 6411 20927
rect 6837 20893 6871 20927
rect 7205 20893 7239 20927
rect 8033 20893 8067 20927
rect 10241 20893 10275 20927
rect 10334 20893 10368 20927
rect 10706 20893 10740 20927
rect 13737 20893 13771 20927
rect 13829 20893 13863 20927
rect 14473 20893 14507 20927
rect 14657 20893 14691 20927
rect 14749 20893 14783 20927
rect 14933 20893 14967 20927
rect 17049 20893 17083 20927
rect 18429 20893 18463 20927
rect 18521 20893 18555 20927
rect 18705 20893 18739 20927
rect 19901 20893 19935 20927
rect 20269 20893 20303 20927
rect 20453 20893 20487 20927
rect 23581 20893 23615 20927
rect 23857 20893 23891 20927
rect 28825 20893 28859 20927
rect 28917 20893 28951 20927
rect 29009 20893 29043 20927
rect 29929 20893 29963 20927
rect 30113 20893 30147 20927
rect 30205 20893 30239 20927
rect 32229 20893 32263 20927
rect 33701 20893 33735 20927
rect 33793 20893 33827 20927
rect 34161 20893 34195 20927
rect 35725 20893 35759 20927
rect 36829 20893 36863 20927
rect 38761 20893 38795 20927
rect 2145 20825 2179 20859
rect 4813 20825 4847 20859
rect 5273 20825 5307 20859
rect 6929 20825 6963 20859
rect 7021 20825 7055 20859
rect 10517 20825 10551 20859
rect 10609 20825 10643 20859
rect 11253 20825 11287 20859
rect 13553 20825 13587 20859
rect 17325 20825 17359 20859
rect 19257 20825 19291 20859
rect 20821 20825 20855 20859
rect 26249 20825 26283 20859
rect 26433 20825 26467 20859
rect 29193 20825 29227 20859
rect 29285 20825 29319 20859
rect 29745 20825 29779 20859
rect 31217 20825 31251 20859
rect 33885 20825 33919 20859
rect 34023 20825 34057 20859
rect 36553 20825 36587 20859
rect 3617 20757 3651 20791
rect 4445 20757 4479 20791
rect 8125 20757 8159 20791
rect 12817 20757 12851 20791
rect 14289 20757 14323 20791
rect 14749 20757 14783 20791
rect 17141 20757 17175 20791
rect 22109 20757 22143 20791
rect 26617 20757 26651 20791
rect 31309 20757 31343 20791
rect 33517 20757 33551 20791
rect 35909 20757 35943 20791
rect 38485 20757 38519 20791
rect 5273 20553 5307 20587
rect 5917 20553 5951 20587
rect 6377 20553 6411 20587
rect 10333 20553 10367 20587
rect 11805 20553 11839 20587
rect 12173 20553 12207 20587
rect 15853 20553 15887 20587
rect 18613 20553 18647 20587
rect 26709 20553 26743 20587
rect 33793 20553 33827 20587
rect 5549 20485 5583 20519
rect 5641 20485 5675 20519
rect 12265 20485 12299 20519
rect 13921 20485 13955 20519
rect 14105 20485 14139 20519
rect 18245 20485 18279 20519
rect 18445 20485 18479 20519
rect 24961 20485 24995 20519
rect 25421 20485 25455 20519
rect 26536 20485 26570 20519
rect 28733 20485 28767 20519
rect 31375 20485 31409 20519
rect 32781 20485 32815 20519
rect 38393 20485 38427 20519
rect 3065 20417 3099 20451
rect 5365 20417 5399 20451
rect 5733 20417 5767 20451
rect 6561 20417 6595 20451
rect 6745 20417 6779 20451
rect 6837 20417 6871 20451
rect 10977 20417 11011 20451
rect 13369 20417 13403 20451
rect 13553 20417 13587 20451
rect 14381 20417 14415 20451
rect 14749 20417 14783 20451
rect 15485 20417 15519 20451
rect 15669 20417 15703 20451
rect 15761 20417 15795 20451
rect 16313 20417 16347 20451
rect 20913 20417 20947 20451
rect 22753 20417 22787 20451
rect 22845 20417 22879 20451
rect 23029 20417 23063 20451
rect 25053 20417 25087 20451
rect 25513 20417 25547 20451
rect 25789 20417 25823 20451
rect 26249 20417 26283 20451
rect 26617 20417 26651 20451
rect 26801 20417 26835 20451
rect 27353 20417 27387 20451
rect 27445 20417 27479 20451
rect 27629 20417 27663 20451
rect 27721 20417 27755 20451
rect 27905 20417 27939 20451
rect 27997 20417 28031 20451
rect 28273 20417 28307 20451
rect 29009 20417 29043 20451
rect 29837 20417 29871 20451
rect 29929 20417 29963 20451
rect 30113 20417 30147 20451
rect 30205 20417 30239 20451
rect 31493 20417 31527 20451
rect 31585 20417 31619 20451
rect 31677 20417 31711 20451
rect 32505 20417 32539 20451
rect 32689 20417 32723 20451
rect 32873 20417 32907 20451
rect 33977 20417 34011 20451
rect 38117 20417 38151 20451
rect 38210 20417 38244 20451
rect 38485 20417 38519 20451
rect 38582 20417 38616 20451
rect 3157 20349 3191 20383
rect 3341 20349 3375 20383
rect 3525 20349 3559 20383
rect 3801 20349 3835 20383
rect 8585 20349 8619 20383
rect 8861 20349 8895 20383
rect 12357 20349 12391 20383
rect 14197 20349 14231 20383
rect 14841 20349 14875 20383
rect 15117 20349 15151 20383
rect 20637 20349 20671 20383
rect 23213 20349 23247 20383
rect 25329 20349 25363 20383
rect 25605 20349 25639 20383
rect 26433 20349 26467 20383
rect 28089 20349 28123 20383
rect 28641 20349 28675 20383
rect 29193 20349 29227 20383
rect 29653 20349 29687 20383
rect 31217 20349 31251 20383
rect 34161 20349 34195 20383
rect 2697 20281 2731 20315
rect 13277 20281 13311 20315
rect 20361 20281 20395 20315
rect 22937 20281 22971 20315
rect 25237 20281 25271 20315
rect 25973 20281 26007 20315
rect 26065 20281 26099 20315
rect 10425 20213 10459 20247
rect 13737 20213 13771 20247
rect 13921 20213 13955 20247
rect 15577 20213 15611 20247
rect 18429 20213 18463 20247
rect 20545 20213 20579 20247
rect 25513 20213 25547 20247
rect 26249 20213 26283 20247
rect 27997 20213 28031 20247
rect 28457 20213 28491 20247
rect 31861 20213 31895 20247
rect 33057 20213 33091 20247
rect 38761 20213 38795 20247
rect 3801 20009 3835 20043
rect 6101 20009 6135 20043
rect 6745 20009 6779 20043
rect 8033 20009 8067 20043
rect 9321 20009 9355 20043
rect 10149 20009 10183 20043
rect 13553 20009 13587 20043
rect 13737 20009 13771 20043
rect 14381 20009 14415 20043
rect 14473 20009 14507 20043
rect 20085 20009 20119 20043
rect 22845 20009 22879 20043
rect 25053 20009 25087 20043
rect 25329 20009 25363 20043
rect 25513 20009 25547 20043
rect 26065 20009 26099 20043
rect 26525 20009 26559 20043
rect 27905 20009 27939 20043
rect 6837 19941 6871 19975
rect 13185 19941 13219 19975
rect 21281 19941 21315 19975
rect 21373 19941 21407 19975
rect 21649 19941 21683 19975
rect 23213 19941 23247 19975
rect 27813 19941 27847 19975
rect 29101 19941 29135 19975
rect 4353 19873 4387 19907
rect 8769 19873 8803 19907
rect 9781 19873 9815 19907
rect 9873 19873 9907 19907
rect 12541 19873 12575 19907
rect 13277 19873 13311 19907
rect 21005 19873 21039 19907
rect 21097 19873 21131 19907
rect 23305 19873 23339 19907
rect 26433 19873 26467 19907
rect 29837 19873 29871 19907
rect 38945 19873 38979 19907
rect 39313 19873 39347 19907
rect 5089 19805 5123 19839
rect 5549 19805 5583 19839
rect 5733 19805 5767 19839
rect 5917 19805 5951 19839
rect 6193 19805 6227 19839
rect 6377 19805 6411 19839
rect 6469 19805 6503 19839
rect 6561 19805 6595 19839
rect 7021 19805 7055 19839
rect 7297 19805 7331 19839
rect 7573 19805 7607 19839
rect 7849 19805 7883 19839
rect 9689 19805 9723 19839
rect 10333 19805 10367 19839
rect 10701 19805 10735 19839
rect 12449 19805 12483 19839
rect 12817 19805 12851 19839
rect 13001 19805 13035 19839
rect 14105 19805 14139 19839
rect 14197 19805 14231 19839
rect 14611 19805 14645 19839
rect 14841 19805 14875 19839
rect 14969 19805 15003 19839
rect 15117 19805 15151 19839
rect 15393 19805 15427 19839
rect 15485 19805 15519 19839
rect 15669 19805 15703 19839
rect 15761 19805 15795 19839
rect 20269 19805 20303 19839
rect 20361 19805 20395 19839
rect 20545 19805 20579 19839
rect 20637 19805 20671 19839
rect 20821 19805 20855 19839
rect 20913 19805 20947 19839
rect 21557 19805 21591 19839
rect 21741 19805 21775 19839
rect 21833 19805 21867 19839
rect 23029 19805 23063 19839
rect 23765 19805 23799 19839
rect 24409 19805 24443 19839
rect 24593 19805 24627 19839
rect 24685 19805 24719 19839
rect 24777 19805 24811 19839
rect 26249 19805 26283 19839
rect 27353 19805 27387 19839
rect 27629 19805 27663 19839
rect 28273 19805 28307 19839
rect 29285 19805 29319 19839
rect 30113 19805 30147 19839
rect 31125 19805 31159 19839
rect 31309 19805 31343 19839
rect 31493 19805 31527 19839
rect 36829 19805 36863 19839
rect 36922 19805 36956 19839
rect 37294 19805 37328 19839
rect 38853 19805 38887 19839
rect 39129 19805 39163 19839
rect 5825 19737 5859 19771
rect 7665 19737 7699 19771
rect 10425 19737 10459 19771
rect 10517 19737 10551 19771
rect 13737 19737 13771 19771
rect 13933 19737 13967 19771
rect 14381 19737 14415 19771
rect 14749 19737 14783 19771
rect 25145 19737 25179 19771
rect 25361 19737 25395 19771
rect 26525 19737 26559 19771
rect 28089 19737 28123 19771
rect 31401 19737 31435 19771
rect 37105 19737 37139 19771
rect 37197 19737 37231 19771
rect 38577 19737 38611 19771
rect 4537 19669 4571 19703
rect 7205 19669 7239 19703
rect 8125 19669 8159 19703
rect 15209 19669 15243 19703
rect 23581 19669 23615 19703
rect 27445 19669 27479 19703
rect 31677 19669 31711 19703
rect 37473 19669 37507 19703
rect 3433 19465 3467 19499
rect 3893 19465 3927 19499
rect 8677 19465 8711 19499
rect 10517 19465 10551 19499
rect 13737 19465 13771 19499
rect 14289 19465 14323 19499
rect 15209 19465 15243 19499
rect 15669 19465 15703 19499
rect 17141 19465 17175 19499
rect 17233 19465 17267 19499
rect 18429 19465 18463 19499
rect 22017 19465 22051 19499
rect 23397 19465 23431 19499
rect 24041 19465 24075 19499
rect 27445 19465 27479 19499
rect 28917 19465 28951 19499
rect 30297 19465 30331 19499
rect 35173 19465 35207 19499
rect 35449 19465 35483 19499
rect 36737 19465 36771 19499
rect 38660 19465 38694 19499
rect 3985 19397 4019 19431
rect 6745 19397 6779 19431
rect 17693 19397 17727 19431
rect 17969 19397 18003 19431
rect 18245 19397 18279 19431
rect 27613 19397 27647 19431
rect 27813 19397 27847 19431
rect 31585 19397 31619 19431
rect 33951 19397 33985 19431
rect 34161 19397 34195 19431
rect 34529 19397 34563 19431
rect 36277 19397 36311 19431
rect 31355 19363 31389 19397
rect 5825 19329 5859 19363
rect 6561 19329 6595 19363
rect 6837 19329 6871 19363
rect 6929 19329 6963 19363
rect 8769 19329 8803 19363
rect 13829 19329 13863 19363
rect 14013 19329 14047 19363
rect 14473 19329 14507 19363
rect 14657 19329 14691 19363
rect 14749 19329 14783 19363
rect 15393 19329 15427 19363
rect 15945 19329 15979 19363
rect 16221 19329 16255 19363
rect 16405 19329 16439 19363
rect 17049 19329 17083 19363
rect 17417 19329 17451 19363
rect 17596 19329 17630 19363
rect 17785 19329 17819 19363
rect 18521 19329 18555 19363
rect 21833 19329 21867 19363
rect 22109 19329 22143 19363
rect 23581 19329 23615 19363
rect 23857 19329 23891 19363
rect 28733 19329 28767 19363
rect 29285 19329 29319 19363
rect 29561 19329 29595 19363
rect 29929 19329 29963 19363
rect 30481 19329 30515 19363
rect 34069 19329 34103 19363
rect 34253 19329 34287 19363
rect 34437 19329 34471 19363
rect 34713 19329 34747 19363
rect 34989 19329 35023 19363
rect 35633 19329 35667 19363
rect 35725 19329 35759 19363
rect 35817 19329 35851 19363
rect 36001 19329 36035 19363
rect 36461 19329 36495 19363
rect 36553 19329 36587 19363
rect 38393 19329 38427 19363
rect 39037 19329 39071 19363
rect 1685 19261 1719 19295
rect 1961 19261 1995 19295
rect 4077 19261 4111 19295
rect 4905 19261 4939 19295
rect 6377 19261 6411 19295
rect 7205 19261 7239 19295
rect 9045 19261 9079 19295
rect 11161 19261 11195 19295
rect 15577 19261 15611 19295
rect 15669 19261 15703 19295
rect 17877 19261 17911 19295
rect 23765 19261 23799 19295
rect 29101 19261 29135 19295
rect 30113 19261 30147 19295
rect 30205 19261 30239 19295
rect 30665 19261 30699 19295
rect 33793 19261 33827 19295
rect 34897 19261 34931 19295
rect 3525 19193 3559 19227
rect 15853 19193 15887 19227
rect 16865 19193 16899 19227
rect 18245 19193 18279 19227
rect 21833 19193 21867 19227
rect 29377 19193 29411 19227
rect 29469 19193 29503 19227
rect 4353 19125 4387 19159
rect 5181 19125 5215 19159
rect 10609 19125 10643 19159
rect 16405 19125 16439 19159
rect 27629 19125 27663 19159
rect 29745 19125 29779 19159
rect 31217 19125 31251 19159
rect 31401 19125 31435 19159
rect 36277 19125 36311 19159
rect 38669 19125 38703 19159
rect 3341 18921 3375 18955
rect 7665 18921 7699 18955
rect 9505 18921 9539 18955
rect 12633 18921 12667 18955
rect 15853 18921 15887 18955
rect 20821 18921 20855 18955
rect 21649 18921 21683 18955
rect 24685 18921 24719 18955
rect 25145 18921 25179 18955
rect 26157 18921 26191 18955
rect 26893 18921 26927 18955
rect 27077 18921 27111 18955
rect 27445 18921 27479 18955
rect 27629 18921 27663 18955
rect 29745 18921 29779 18955
rect 20453 18853 20487 18887
rect 28181 18853 28215 18887
rect 29285 18853 29319 18887
rect 1593 18785 1627 18819
rect 4905 18785 4939 18819
rect 5181 18785 5215 18819
rect 8309 18785 8343 18819
rect 10149 18785 10183 18819
rect 35081 18785 35115 18819
rect 39313 18785 39347 18819
rect 4721 18717 4755 18751
rect 4813 18717 4847 18751
rect 8033 18717 8067 18751
rect 9229 18717 9263 18751
rect 9413 18717 9447 18751
rect 9873 18717 9907 18751
rect 10885 18717 10919 18751
rect 13277 18717 13311 18751
rect 15945 18717 15979 18751
rect 20361 18717 20395 18751
rect 20637 18717 20671 18751
rect 20913 18717 20947 18751
rect 21097 18717 21131 18751
rect 21925 18717 21959 18751
rect 22017 18717 22051 18751
rect 22109 18717 22143 18751
rect 22293 18717 22327 18751
rect 25697 18717 25731 18751
rect 25789 18717 25823 18751
rect 25881 18717 25915 18751
rect 25973 18717 26007 18751
rect 28549 18717 28583 18751
rect 29101 18717 29135 18751
rect 29377 18717 29411 18751
rect 30205 18717 30239 18751
rect 30297 18717 30331 18751
rect 31033 18717 31067 18751
rect 31217 18717 31251 18751
rect 31401 18717 31435 18751
rect 31677 18717 31711 18751
rect 34897 18717 34931 18751
rect 35633 18717 35667 18751
rect 35817 18717 35851 18751
rect 35909 18717 35943 18751
rect 36001 18717 36035 18751
rect 39037 18717 39071 18751
rect 39221 18717 39255 18751
rect 27031 18683 27065 18717
rect 1869 18649 1903 18683
rect 5457 18649 5491 18683
rect 11161 18649 11195 18683
rect 24869 18649 24903 18683
rect 25329 18649 25363 18683
rect 27261 18649 27295 18683
rect 27813 18649 27847 18683
rect 28365 18649 28399 18683
rect 28917 18649 28951 18683
rect 29653 18649 29687 18683
rect 31309 18649 31343 18683
rect 31861 18649 31895 18683
rect 4353 18581 4387 18615
rect 6929 18581 6963 18615
rect 8125 18581 8159 18615
rect 9321 18581 9355 18615
rect 9965 18581 9999 18615
rect 12725 18581 12759 18615
rect 21281 18581 21315 18615
rect 24501 18581 24535 18615
rect 24685 18581 24719 18615
rect 24961 18581 24995 18615
rect 25129 18581 25163 18615
rect 27603 18581 27637 18615
rect 28733 18581 28767 18615
rect 30481 18581 30515 18615
rect 31585 18581 31619 18615
rect 32045 18581 32079 18615
rect 34713 18581 34747 18615
rect 36185 18581 36219 18615
rect 38853 18581 38887 18615
rect 2697 18377 2731 18411
rect 3157 18377 3191 18411
rect 6377 18377 6411 18411
rect 11713 18377 11747 18411
rect 12081 18377 12115 18411
rect 14289 18377 14323 18411
rect 15945 18377 15979 18411
rect 16773 18377 16807 18411
rect 26801 18377 26835 18411
rect 4077 18309 4111 18343
rect 6837 18309 6871 18343
rect 12173 18309 12207 18343
rect 27905 18309 27939 18343
rect 32321 18309 32355 18343
rect 3065 18241 3099 18275
rect 3801 18241 3835 18275
rect 6745 18241 6779 18275
rect 7205 18241 7239 18275
rect 7757 18241 7791 18275
rect 15577 18241 15611 18275
rect 16129 18241 16163 18275
rect 16405 18241 16439 18275
rect 17049 18241 17083 18275
rect 22109 18241 22143 18275
rect 22201 18241 22235 18275
rect 22385 18241 22419 18275
rect 22477 18241 22511 18275
rect 24409 18241 24443 18275
rect 24685 18241 24719 18275
rect 26157 18241 26191 18275
rect 26341 18241 26375 18275
rect 26433 18241 26467 18275
rect 26525 18241 26559 18275
rect 27169 18241 27203 18275
rect 27353 18241 27387 18275
rect 28089 18241 28123 18275
rect 30573 18241 30607 18275
rect 32137 18241 32171 18275
rect 38209 18241 38243 18275
rect 38393 18241 38427 18275
rect 38577 18241 38611 18275
rect 3341 18173 3375 18207
rect 5549 18173 5583 18207
rect 7021 18173 7055 18207
rect 12265 18173 12299 18207
rect 12541 18173 12575 18207
rect 12817 18173 12851 18207
rect 15393 18173 15427 18207
rect 15853 18173 15887 18207
rect 16221 18173 16255 18207
rect 24501 18173 24535 18207
rect 30757 18173 30791 18207
rect 38485 18173 38519 18207
rect 39313 18173 39347 18207
rect 39405 18173 39439 18207
rect 39681 18173 39715 18207
rect 16313 18105 16347 18139
rect 24593 18105 24627 18139
rect 30389 18105 30423 18139
rect 38669 18105 38703 18139
rect 15761 18037 15795 18071
rect 22661 18037 22695 18071
rect 24225 18037 24259 18071
rect 26985 18037 27019 18071
rect 27813 18037 27847 18071
rect 32505 18037 32539 18071
rect 38945 18037 38979 18071
rect 12817 17833 12851 17867
rect 16589 17833 16623 17867
rect 17049 17833 17083 17867
rect 18429 17833 18463 17867
rect 24869 17833 24903 17867
rect 26525 17833 26559 17867
rect 32965 17833 32999 17867
rect 34069 17833 34103 17867
rect 38577 17833 38611 17867
rect 22937 17765 22971 17799
rect 31677 17765 31711 17799
rect 4445 17697 4479 17731
rect 5273 17697 5307 17731
rect 9413 17697 9447 17731
rect 13461 17697 13495 17731
rect 21649 17697 21683 17731
rect 22845 17697 22879 17731
rect 24961 17697 24995 17731
rect 26433 17697 26467 17731
rect 28365 17697 28399 17731
rect 38577 17697 38611 17731
rect 7389 17629 7423 17663
rect 8585 17629 8619 17663
rect 8769 17629 8803 17663
rect 9229 17629 9263 17663
rect 9689 17629 9723 17663
rect 9873 17629 9907 17663
rect 10977 17629 11011 17663
rect 11161 17629 11195 17663
rect 16773 17629 16807 17663
rect 16865 17629 16899 17663
rect 18245 17629 18279 17663
rect 18521 17629 18555 17663
rect 22201 17629 22235 17663
rect 22385 17629 22419 17663
rect 22661 17629 22695 17663
rect 23121 17629 23155 17663
rect 23489 17629 23523 17663
rect 24685 17629 24719 17663
rect 26525 17629 26559 17663
rect 28549 17629 28583 17663
rect 28641 17629 28675 17663
rect 28825 17629 28859 17663
rect 28917 17629 28951 17663
rect 31125 17629 31159 17663
rect 31493 17629 31527 17663
rect 31861 17629 31895 17663
rect 32321 17629 32355 17663
rect 32505 17629 32539 17663
rect 32781 17629 32815 17663
rect 32965 17629 32999 17663
rect 33333 17629 33367 17663
rect 33701 17629 33735 17663
rect 33977 17629 34011 17663
rect 34161 17629 34195 17663
rect 34253 17629 34287 17663
rect 36093 17629 36127 17663
rect 36186 17629 36220 17663
rect 36558 17629 36592 17663
rect 38393 17629 38427 17663
rect 4169 17561 4203 17595
rect 4629 17561 4663 17595
rect 7205 17561 7239 17595
rect 13185 17561 13219 17595
rect 17049 17561 17083 17595
rect 23213 17561 23247 17595
rect 23305 17561 23339 17595
rect 26249 17561 26283 17595
rect 31309 17561 31343 17595
rect 31401 17561 31435 17595
rect 32413 17561 32447 17595
rect 33517 17561 33551 17595
rect 33609 17561 33643 17595
rect 36369 17561 36403 17595
rect 36461 17561 36495 17595
rect 38669 17561 38703 17595
rect 3801 17493 3835 17527
rect 4261 17493 4295 17527
rect 7021 17493 7055 17527
rect 8677 17493 8711 17527
rect 9045 17493 9079 17527
rect 9873 17493 9907 17527
rect 11161 17493 11195 17527
rect 13277 17493 13311 17527
rect 18061 17493 18095 17527
rect 24501 17493 24535 17527
rect 26709 17493 26743 17527
rect 31953 17493 31987 17527
rect 33149 17493 33183 17527
rect 33885 17493 33919 17527
rect 34437 17493 34471 17527
rect 36737 17493 36771 17527
rect 38209 17493 38243 17527
rect 4261 17289 4295 17323
rect 10977 17289 11011 17323
rect 18429 17289 18463 17323
rect 24409 17289 24443 17323
rect 29009 17289 29043 17323
rect 33793 17289 33827 17323
rect 38393 17289 38427 17323
rect 2789 17221 2823 17255
rect 9781 17221 9815 17255
rect 10885 17221 10919 17255
rect 14013 17221 14047 17255
rect 18613 17221 18647 17255
rect 19041 17221 19075 17255
rect 19257 17221 19291 17255
rect 19625 17221 19659 17255
rect 23949 17221 23983 17255
rect 24501 17221 24535 17255
rect 28733 17221 28767 17255
rect 37933 17221 37967 17255
rect 2513 17153 2547 17187
rect 7113 17153 7147 17187
rect 7297 17153 7331 17187
rect 7573 17153 7607 17187
rect 7757 17153 7791 17187
rect 7941 17153 7975 17187
rect 8125 17153 8159 17187
rect 9597 17153 9631 17187
rect 9873 17153 9907 17187
rect 11805 17153 11839 17187
rect 13829 17153 13863 17187
rect 16957 17153 16991 17187
rect 17049 17153 17083 17187
rect 17325 17153 17359 17187
rect 18797 17153 18831 17187
rect 19441 17153 19475 17187
rect 19717 17153 19751 17187
rect 19809 17153 19843 17187
rect 24225 17153 24259 17187
rect 24685 17153 24719 17187
rect 27169 17153 27203 17187
rect 28354 17153 28388 17187
rect 28485 17153 28519 17187
rect 28641 17153 28675 17187
rect 28849 17153 28883 17187
rect 30113 17153 30147 17187
rect 30297 17153 30331 17187
rect 33701 17153 33735 17187
rect 33885 17153 33919 17187
rect 35081 17153 35115 17187
rect 35229 17153 35263 17187
rect 35357 17153 35391 17187
rect 35449 17153 35483 17187
rect 35587 17153 35621 17187
rect 35909 17153 35943 17187
rect 38117 17153 38151 17187
rect 38209 17153 38243 17187
rect 7205 17085 7239 17119
rect 11069 17085 11103 17119
rect 24041 17085 24075 17119
rect 24961 17085 24995 17119
rect 26985 17085 27019 17119
rect 27445 17085 27479 17119
rect 27997 17085 28031 17119
rect 30389 17085 30423 17119
rect 10517 17017 10551 17051
rect 17233 17017 17267 17051
rect 18889 17017 18923 17051
rect 36093 17017 36127 17051
rect 7389 16949 7423 16983
rect 8033 16949 8067 16983
rect 9413 16949 9447 16983
rect 11897 16949 11931 16983
rect 13645 16949 13679 16983
rect 16773 16949 16807 16983
rect 19073 16949 19107 16983
rect 19993 16949 20027 16983
rect 23949 16949 23983 16983
rect 24869 16949 24903 16983
rect 29929 16949 29963 16983
rect 35725 16949 35759 16983
rect 37933 16949 37967 16983
rect 6561 16745 6595 16779
rect 7297 16745 7331 16779
rect 7849 16745 7883 16779
rect 8217 16745 8251 16779
rect 13001 16745 13035 16779
rect 21189 16745 21223 16779
rect 21281 16745 21315 16779
rect 22293 16745 22327 16779
rect 22753 16745 22787 16779
rect 22937 16745 22971 16779
rect 26801 16745 26835 16779
rect 28181 16745 28215 16779
rect 38393 16745 38427 16779
rect 7021 16677 7055 16711
rect 7113 16677 7147 16711
rect 21649 16677 21683 16711
rect 26525 16677 26559 16711
rect 37105 16677 37139 16711
rect 4813 16609 4847 16643
rect 5089 16609 5123 16643
rect 7665 16609 7699 16643
rect 8125 16609 8159 16643
rect 9413 16609 9447 16643
rect 9505 16609 9539 16643
rect 10517 16609 10551 16643
rect 11345 16609 11379 16643
rect 11713 16609 11747 16643
rect 13737 16609 13771 16643
rect 14381 16609 14415 16643
rect 15025 16609 15059 16643
rect 20545 16609 20579 16643
rect 21373 16609 21407 16643
rect 22385 16609 22419 16643
rect 22937 16609 22971 16643
rect 25697 16609 25731 16643
rect 26341 16609 26375 16643
rect 38485 16609 38519 16643
rect 6745 16541 6779 16575
rect 7941 16541 7975 16575
rect 8033 16541 8067 16575
rect 10241 16541 10275 16575
rect 11161 16541 11195 16575
rect 11897 16541 11931 16575
rect 14105 16541 14139 16575
rect 14565 16541 14599 16575
rect 14657 16541 14691 16575
rect 14841 16541 14875 16575
rect 16773 16541 16807 16575
rect 16865 16541 16899 16575
rect 17049 16541 17083 16575
rect 17141 16541 17175 16575
rect 21005 16541 21039 16575
rect 21281 16541 21315 16575
rect 22569 16541 22603 16575
rect 22845 16541 22879 16575
rect 25329 16541 25363 16575
rect 25513 16541 25547 16575
rect 25789 16531 25823 16565
rect 26065 16541 26099 16575
rect 26249 16541 26283 16575
rect 26433 16541 26467 16575
rect 28360 16541 28394 16575
rect 28677 16541 28711 16575
rect 28825 16541 28859 16575
rect 36461 16541 36495 16575
rect 36609 16541 36643 16575
rect 36737 16541 36771 16575
rect 36967 16541 37001 16575
rect 38393 16541 38427 16575
rect 6837 16473 6871 16507
rect 7021 16473 7055 16507
rect 7481 16473 7515 16507
rect 9321 16473 9355 16507
rect 10333 16473 10367 16507
rect 11069 16473 11103 16507
rect 11805 16473 11839 16507
rect 12449 16473 12483 16507
rect 12725 16473 12759 16507
rect 13645 16473 13679 16507
rect 20703 16473 20737 16507
rect 20821 16473 20855 16507
rect 20913 16473 20947 16507
rect 22293 16473 22327 16507
rect 24777 16473 24811 16507
rect 28457 16473 28491 16507
rect 28549 16473 28583 16507
rect 36829 16473 36863 16507
rect 7281 16405 7315 16439
rect 7665 16405 7699 16439
rect 8401 16405 8435 16439
rect 8953 16405 8987 16439
rect 9873 16405 9907 16439
rect 10701 16405 10735 16439
rect 12265 16405 12299 16439
rect 12541 16405 12575 16439
rect 13185 16405 13219 16439
rect 13553 16405 13587 16439
rect 14197 16405 14231 16439
rect 16589 16405 16623 16439
rect 23213 16405 23247 16439
rect 38761 16405 38795 16439
rect 4721 16201 4755 16235
rect 5273 16201 5307 16235
rect 7481 16201 7515 16235
rect 8309 16201 8343 16235
rect 9505 16201 9539 16235
rect 10977 16201 11011 16235
rect 11897 16201 11931 16235
rect 26985 16201 27019 16235
rect 30021 16201 30055 16235
rect 10885 16133 10919 16167
rect 12541 16133 12575 16167
rect 13997 16133 14031 16167
rect 14197 16133 14231 16167
rect 14841 16133 14875 16167
rect 24133 16133 24167 16167
rect 30389 16133 30423 16167
rect 31309 16133 31343 16167
rect 34299 16133 34333 16167
rect 34437 16133 34471 16167
rect 35173 16133 35207 16167
rect 36829 16133 36863 16167
rect 2973 16065 3007 16099
rect 5181 16065 5215 16099
rect 7481 16065 7515 16099
rect 7665 16065 7699 16099
rect 8493 16065 8527 16099
rect 8677 16065 8711 16099
rect 9413 16065 9447 16099
rect 11989 16065 12023 16099
rect 12725 16065 12759 16099
rect 13369 16065 13403 16099
rect 13645 16065 13679 16099
rect 15025 16065 15059 16099
rect 15209 16065 15243 16099
rect 15853 16065 15887 16099
rect 16037 16065 16071 16099
rect 16129 16065 16163 16099
rect 16313 16065 16347 16099
rect 16405 16065 16439 16099
rect 24317 16065 24351 16099
rect 24501 16065 24535 16099
rect 24593 16065 24627 16099
rect 27169 16065 27203 16099
rect 27445 16065 27479 16099
rect 27629 16065 27663 16099
rect 28181 16065 28215 16099
rect 28365 16065 28399 16099
rect 30205 16065 30239 16099
rect 30297 16065 30331 16099
rect 30573 16065 30607 16099
rect 31171 16065 31205 16099
rect 31401 16065 31435 16099
rect 31493 16065 31527 16099
rect 34161 16065 34195 16099
rect 34529 16065 34563 16099
rect 34621 16065 34655 16099
rect 34897 16065 34931 16099
rect 36553 16065 36587 16099
rect 36737 16065 36771 16099
rect 36921 16065 36955 16099
rect 3249 15997 3283 16031
rect 5365 15997 5399 16031
rect 11069 15997 11103 16031
rect 12081 15997 12115 16031
rect 13553 15997 13587 16031
rect 28089 15997 28123 16031
rect 31033 15997 31067 16031
rect 34805 15997 34839 16031
rect 4813 15929 4847 15963
rect 10517 15929 10551 15963
rect 13461 15929 13495 15963
rect 27353 15929 27387 15963
rect 31677 15929 31711 15963
rect 11529 15861 11563 15895
rect 12357 15861 12391 15895
rect 13185 15861 13219 15895
rect 13829 15861 13863 15895
rect 14013 15861 14047 15895
rect 27905 15861 27939 15895
rect 27997 15861 28031 15895
rect 37105 15861 37139 15895
rect 5457 15657 5491 15691
rect 6193 15657 6227 15691
rect 10241 15657 10275 15691
rect 16405 15657 16439 15691
rect 16865 15657 16899 15691
rect 17049 15657 17083 15691
rect 17417 15657 17451 15691
rect 22017 15657 22051 15691
rect 33057 15657 33091 15691
rect 34989 15657 35023 15691
rect 35357 15657 35391 15691
rect 38301 15657 38335 15691
rect 7021 15589 7055 15623
rect 31401 15589 31435 15623
rect 39221 15589 39255 15623
rect 4905 15521 4939 15555
rect 10333 15521 10367 15555
rect 10517 15521 10551 15555
rect 11345 15521 11379 15555
rect 17141 15521 17175 15555
rect 22293 15521 22327 15555
rect 22385 15521 22419 15555
rect 25145 15521 25179 15555
rect 29653 15521 29687 15555
rect 29929 15521 29963 15555
rect 35081 15521 35115 15555
rect 38485 15521 38519 15555
rect 38853 15521 38887 15555
rect 39313 15521 39347 15555
rect 5549 15453 5583 15487
rect 5642 15453 5676 15487
rect 6055 15453 6089 15487
rect 6285 15453 6319 15487
rect 6469 15453 6503 15487
rect 6837 15453 6871 15487
rect 7021 15453 7055 15487
rect 8033 15453 8067 15487
rect 10057 15453 10091 15487
rect 10425 15453 10459 15487
rect 11621 15453 11655 15487
rect 11713 15453 11747 15487
rect 11805 15453 11839 15487
rect 11989 15453 12023 15487
rect 13185 15453 13219 15487
rect 16589 15453 16623 15487
rect 16681 15453 16715 15487
rect 16865 15453 16899 15487
rect 16957 15453 16991 15487
rect 17233 15453 17267 15487
rect 18153 15453 18187 15487
rect 18337 15453 18371 15487
rect 18429 15453 18463 15487
rect 20361 15453 20395 15487
rect 20637 15453 20671 15487
rect 22201 15453 22235 15487
rect 22477 15453 22511 15487
rect 24225 15453 24259 15487
rect 24409 15453 24443 15487
rect 24777 15453 24811 15487
rect 25513 15453 25547 15487
rect 25697 15453 25731 15487
rect 28917 15453 28951 15487
rect 29009 15453 29043 15487
rect 29193 15453 29227 15487
rect 29285 15453 29319 15487
rect 29837 15453 29871 15487
rect 30021 15453 30055 15487
rect 30113 15453 30147 15487
rect 30481 15453 30515 15487
rect 30849 15453 30883 15487
rect 31033 15453 31067 15487
rect 31217 15453 31251 15487
rect 31493 15453 31527 15487
rect 31586 15453 31620 15487
rect 31958 15453 31992 15487
rect 32413 15453 32447 15487
rect 32506 15453 32540 15487
rect 32878 15453 32912 15487
rect 34989 15453 35023 15487
rect 38577 15453 38611 15487
rect 39037 15453 39071 15487
rect 5825 15385 5859 15419
rect 5917 15385 5951 15419
rect 10701 15385 10735 15419
rect 20177 15385 20211 15419
rect 23857 15385 23891 15419
rect 24041 15385 24075 15419
rect 30665 15385 30699 15419
rect 31125 15385 31159 15419
rect 31769 15385 31803 15419
rect 31861 15385 31895 15419
rect 32689 15385 32723 15419
rect 32781 15385 32815 15419
rect 38301 15385 38335 15419
rect 4997 15317 5031 15351
rect 5089 15317 5123 15351
rect 6469 15317 6503 15351
rect 7941 15317 7975 15351
rect 9873 15317 9907 15351
rect 10425 15317 10459 15351
rect 13369 15317 13403 15351
rect 17969 15317 18003 15351
rect 20545 15317 20579 15351
rect 28733 15317 28767 15351
rect 30297 15317 30331 15351
rect 32137 15317 32171 15351
rect 38761 15317 38795 15351
rect 4629 15113 4663 15147
rect 5273 15113 5307 15147
rect 8677 15113 8711 15147
rect 13829 15113 13863 15147
rect 20545 15113 20579 15147
rect 22753 15113 22787 15147
rect 24593 15113 24627 15147
rect 34437 15113 34471 15147
rect 6745 15045 6779 15079
rect 6929 15045 6963 15079
rect 17325 15045 17359 15079
rect 17877 15045 17911 15079
rect 20177 15045 20211 15079
rect 20393 15045 20427 15079
rect 34161 15045 34195 15079
rect 35725 15045 35759 15079
rect 35909 15045 35943 15079
rect 4261 14977 4295 15011
rect 5181 14977 5215 15011
rect 5365 14977 5399 15011
rect 5825 14977 5859 15011
rect 6009 14977 6043 15011
rect 6561 14977 6595 15011
rect 7389 14977 7423 15011
rect 7665 14977 7699 15011
rect 7757 14977 7791 15011
rect 8309 14977 8343 15011
rect 9413 14977 9447 15011
rect 9689 14977 9723 15011
rect 10057 14977 10091 15011
rect 10793 14977 10827 15011
rect 11897 14977 11931 15011
rect 12449 14977 12483 15011
rect 12633 14977 12667 15011
rect 12725 14977 12759 15011
rect 13093 14977 13127 15011
rect 13185 14977 13219 15011
rect 13553 14977 13587 15011
rect 14197 14977 14231 15011
rect 14933 14977 14967 15011
rect 15117 14977 15151 15011
rect 15393 14977 15427 15011
rect 15853 14977 15887 15011
rect 16313 14977 16347 15011
rect 16865 14977 16899 15011
rect 17601 14977 17635 15011
rect 19717 14977 19751 15011
rect 19809 14977 19843 15011
rect 19993 14977 20027 15011
rect 20085 14977 20119 15011
rect 22477 14977 22511 15011
rect 22845 14977 22879 15011
rect 24777 14977 24811 15011
rect 24869 14977 24903 15011
rect 25053 14977 25087 15011
rect 33885 14977 33919 15011
rect 34069 14977 34103 15011
rect 34253 14977 34287 15011
rect 38669 14977 38703 15011
rect 38853 14977 38887 15011
rect 4353 14909 4387 14943
rect 7205 14909 7239 14943
rect 7849 14909 7883 14943
rect 8217 14909 8251 14943
rect 9321 14909 9355 14943
rect 9781 14909 9815 14943
rect 10149 14909 10183 14943
rect 10241 14909 10275 14943
rect 10333 14909 10367 14943
rect 11805 14909 11839 14943
rect 11989 14909 12023 14943
rect 12081 14909 12115 14943
rect 17049 14909 17083 14943
rect 17785 14909 17819 14943
rect 22385 14909 22419 14943
rect 7021 14841 7055 14875
rect 9137 14841 9171 14875
rect 9873 14841 9907 14875
rect 10609 14841 10643 14875
rect 15393 14841 15427 14875
rect 16681 14841 16715 14875
rect 17417 14841 17451 14875
rect 24961 14841 24995 14875
rect 6193 14773 6227 14807
rect 7205 14773 7239 14807
rect 7297 14773 7331 14807
rect 7481 14773 7515 14807
rect 8033 14773 8067 14807
rect 11621 14773 11655 14807
rect 12909 14773 12943 14807
rect 13645 14773 13679 14807
rect 13829 14773 13863 14807
rect 14749 14773 14783 14807
rect 16865 14773 16899 14807
rect 17785 14773 17819 14807
rect 19533 14773 19567 14807
rect 20361 14773 20395 14807
rect 22109 14773 22143 14807
rect 22569 14773 22603 14807
rect 36093 14773 36127 14807
rect 38669 14773 38703 14807
rect 39037 14773 39071 14807
rect 4537 14569 4571 14603
rect 6285 14569 6319 14603
rect 9321 14569 9355 14603
rect 10241 14569 10275 14603
rect 15669 14569 15703 14603
rect 15853 14569 15887 14603
rect 16037 14569 16071 14603
rect 17417 14569 17451 14603
rect 19533 14569 19567 14603
rect 19809 14569 19843 14603
rect 20361 14569 20395 14603
rect 21005 14569 21039 14603
rect 22201 14569 22235 14603
rect 22661 14569 22695 14603
rect 23305 14569 23339 14603
rect 25605 14569 25639 14603
rect 27905 14569 27939 14603
rect 28549 14569 28583 14603
rect 36645 14569 36679 14603
rect 4629 14501 4663 14535
rect 6193 14501 6227 14535
rect 7849 14501 7883 14535
rect 14933 14501 14967 14535
rect 15301 14501 15335 14535
rect 20821 14501 20855 14535
rect 25237 14501 25271 14535
rect 28917 14501 28951 14535
rect 4261 14433 4295 14467
rect 6469 14433 6503 14467
rect 6561 14433 6595 14467
rect 6745 14433 6779 14467
rect 16129 14433 16163 14467
rect 17233 14433 17267 14467
rect 18705 14433 18739 14467
rect 18889 14433 18923 14467
rect 18981 14433 19015 14467
rect 19533 14433 19567 14467
rect 20453 14433 20487 14467
rect 26065 14433 26099 14467
rect 28825 14433 28859 14467
rect 30113 14433 30147 14467
rect 4169 14365 4203 14399
rect 4843 14365 4877 14399
rect 4997 14365 5031 14399
rect 5917 14365 5951 14399
rect 6653 14365 6687 14399
rect 7205 14365 7239 14399
rect 7298 14365 7332 14399
rect 7481 14365 7515 14399
rect 7711 14365 7745 14399
rect 8401 14365 8435 14399
rect 8493 14365 8527 14399
rect 8585 14365 8619 14399
rect 8677 14365 8711 14399
rect 9500 14365 9534 14399
rect 9689 14365 9723 14399
rect 9872 14365 9906 14399
rect 9965 14365 9999 14399
rect 10057 14365 10091 14399
rect 10241 14365 10275 14399
rect 10333 14365 10367 14399
rect 10517 14365 10551 14399
rect 12541 14365 12575 14399
rect 14841 14365 14875 14399
rect 15025 14365 15059 14399
rect 15485 14365 15519 14399
rect 15577 14365 15611 14399
rect 16405 14365 16439 14399
rect 17141 14365 17175 14399
rect 17417 14365 17451 14399
rect 18797 14365 18831 14399
rect 19625 14365 19659 14399
rect 20269 14365 20303 14399
rect 20545 14365 20579 14399
rect 20729 14365 20763 14399
rect 21649 14365 21683 14399
rect 21741 14365 21775 14399
rect 21925 14365 21959 14399
rect 22017 14365 22051 14399
rect 22753 14365 22787 14399
rect 22845 14365 22879 14399
rect 23029 14365 23063 14399
rect 23121 14365 23155 14399
rect 25053 14365 25087 14399
rect 25237 14365 25271 14399
rect 25789 14365 25823 14399
rect 25973 14365 26007 14399
rect 26433 14365 26467 14399
rect 26617 14365 26651 14399
rect 28089 14365 28123 14399
rect 28181 14365 28215 14399
rect 28273 14365 28307 14399
rect 28365 14365 28399 14399
rect 28733 14365 28767 14399
rect 29009 14365 29043 14399
rect 30297 14365 30331 14399
rect 30573 14365 30607 14399
rect 36093 14365 36127 14399
rect 36277 14365 36311 14399
rect 36461 14365 36495 14399
rect 36737 14365 36771 14399
rect 36921 14365 36955 14399
rect 37013 14365 37047 14399
rect 37105 14365 37139 14399
rect 6193 14297 6227 14331
rect 7573 14297 7607 14331
rect 9597 14297 9631 14331
rect 15761 14297 15795 14331
rect 19349 14297 19383 14331
rect 19993 14297 20027 14331
rect 20989 14297 21023 14331
rect 21189 14297 21223 14331
rect 22293 14297 22327 14331
rect 22477 14297 22511 14331
rect 36369 14297 36403 14331
rect 6009 14229 6043 14263
rect 8217 14229 8251 14263
rect 10425 14229 10459 14263
rect 12633 14229 12667 14263
rect 16957 14229 16991 14263
rect 18521 14229 18555 14263
rect 26433 14229 26467 14263
rect 30481 14229 30515 14263
rect 37289 14229 37323 14263
rect 4169 14025 4203 14059
rect 16037 14025 16071 14059
rect 19717 14025 19751 14059
rect 23673 14025 23707 14059
rect 23857 14025 23891 14059
rect 24041 14025 24075 14059
rect 24317 14025 24351 14059
rect 24485 14025 24519 14059
rect 25789 14025 25823 14059
rect 27077 14025 27111 14059
rect 27997 14025 28031 14059
rect 33057 14025 33091 14059
rect 37105 14025 37139 14059
rect 38853 14025 38887 14059
rect 9597 13957 9631 13991
rect 13645 13957 13679 13991
rect 16221 13957 16255 13991
rect 24685 13957 24719 13991
rect 28457 13957 28491 13991
rect 37289 13957 37323 13991
rect 4353 13889 4387 13923
rect 4445 13889 4479 13923
rect 4629 13889 4663 13923
rect 4721 13889 4755 13923
rect 9413 13889 9447 13923
rect 9689 13889 9723 13923
rect 10517 13889 10551 13923
rect 10609 13889 10643 13923
rect 10701 13889 10735 13923
rect 10879 13889 10913 13923
rect 11069 13889 11103 13923
rect 11253 13889 11287 13923
rect 11805 13889 11839 13923
rect 11989 13889 12023 13923
rect 12633 13889 12667 13923
rect 12817 13889 12851 13923
rect 12909 13889 12943 13923
rect 13185 13889 13219 13923
rect 13369 13889 13403 13923
rect 13921 13889 13955 13923
rect 16405 13889 16439 13923
rect 19625 13889 19659 13923
rect 19809 13889 19843 13923
rect 23949 13889 23983 13923
rect 24225 13889 24259 13923
rect 25697 13889 25731 13923
rect 25881 13889 25915 13923
rect 26433 13889 26467 13923
rect 26985 13889 27019 13923
rect 27169 13889 27203 13923
rect 28181 13889 28215 13923
rect 28917 13889 28951 13923
rect 30573 13889 30607 13923
rect 30665 13889 30699 13923
rect 32597 13889 32631 13923
rect 32781 13889 32815 13923
rect 32873 13889 32907 13923
rect 36737 13889 36771 13923
rect 36921 13889 36955 13923
rect 37473 13889 37507 13923
rect 37565 13889 37599 13923
rect 38393 13889 38427 13923
rect 38669 13889 38703 13923
rect 11161 13821 11195 13855
rect 13737 13821 13771 13855
rect 26249 13821 26283 13855
rect 26525 13821 26559 13855
rect 26617 13821 26651 13855
rect 26709 13821 26743 13855
rect 28365 13821 28399 13855
rect 30849 13821 30883 13855
rect 38485 13821 38519 13855
rect 28733 13753 28767 13787
rect 37749 13753 37783 13787
rect 9229 13685 9263 13719
rect 10241 13685 10275 13719
rect 11989 13685 12023 13719
rect 12449 13685 12483 13719
rect 13001 13685 13035 13719
rect 13185 13685 13219 13719
rect 14105 13685 14139 13719
rect 24501 13685 24535 13719
rect 28181 13685 28215 13719
rect 32597 13685 32631 13719
rect 36921 13685 36955 13719
rect 37289 13685 37323 13719
rect 38577 13685 38611 13719
rect 3525 13481 3559 13515
rect 4353 13481 4387 13515
rect 6745 13481 6779 13515
rect 15945 13481 15979 13515
rect 16313 13481 16347 13515
rect 16865 13481 16899 13515
rect 17049 13481 17083 13515
rect 17233 13481 17267 13515
rect 17969 13481 18003 13515
rect 19901 13481 19935 13515
rect 22109 13481 22143 13515
rect 23029 13481 23063 13515
rect 27077 13481 27111 13515
rect 34713 13481 34747 13515
rect 35173 13481 35207 13515
rect 38945 13481 38979 13515
rect 39129 13481 39163 13515
rect 7665 13413 7699 13447
rect 17601 13413 17635 13447
rect 22845 13413 22879 13447
rect 30021 13413 30055 13447
rect 32321 13413 32355 13447
rect 33425 13413 33459 13447
rect 7297 13345 7331 13379
rect 9229 13345 9263 13379
rect 9781 13345 9815 13379
rect 11253 13345 11287 13379
rect 13185 13345 13219 13379
rect 14105 13345 14139 13379
rect 16221 13345 16255 13379
rect 34897 13345 34931 13379
rect 39221 13345 39255 13379
rect 3433 13277 3467 13311
rect 3617 13277 3651 13311
rect 4537 13277 4571 13311
rect 4721 13277 4755 13311
rect 4813 13277 4847 13311
rect 4997 13277 5031 13311
rect 5181 13277 5215 13311
rect 5273 13277 5307 13311
rect 6929 13277 6963 13311
rect 7113 13277 7147 13311
rect 7205 13277 7239 13311
rect 7849 13277 7883 13311
rect 7942 13277 7976 13311
rect 8125 13277 8159 13311
rect 8355 13277 8389 13311
rect 9965 13277 9999 13311
rect 11161 13277 11195 13311
rect 12541 13277 12575 13311
rect 12817 13277 12851 13311
rect 13001 13277 13035 13311
rect 13093 13277 13127 13311
rect 13369 13277 13403 13311
rect 14381 13277 14415 13311
rect 15209 13277 15243 13311
rect 15301 13277 15335 13311
rect 16313 13277 16347 13311
rect 16681 13277 16715 13311
rect 16957 13277 16991 13311
rect 17233 13277 17267 13311
rect 17325 13277 17359 13311
rect 17785 13277 17819 13311
rect 17877 13277 17911 13311
rect 19257 13277 19291 13311
rect 19349 13277 19383 13311
rect 19533 13277 19567 13311
rect 19625 13277 19659 13311
rect 20085 13277 20119 13311
rect 20361 13277 20395 13311
rect 20913 13277 20947 13311
rect 21097 13277 21131 13311
rect 21189 13277 21223 13311
rect 21281 13277 21315 13311
rect 22385 13277 22419 13311
rect 22477 13277 22511 13311
rect 22569 13277 22603 13311
rect 22753 13277 22787 13311
rect 26157 13277 26191 13311
rect 26249 13277 26283 13311
rect 26617 13277 26651 13311
rect 27169 13277 27203 13311
rect 30113 13277 30147 13311
rect 30297 13277 30331 13311
rect 31769 13277 31803 13311
rect 32137 13277 32171 13311
rect 32689 13277 32723 13311
rect 32781 13277 32815 13311
rect 32874 13277 32908 13311
rect 33149 13277 33183 13311
rect 33287 13277 33321 13311
rect 34713 13277 34747 13311
rect 34989 13277 35023 13311
rect 38761 13277 38795 13311
rect 38853 13277 38887 13311
rect 39129 13277 39163 13311
rect 3801 13209 3835 13243
rect 4169 13209 4203 13243
rect 8217 13209 8251 13243
rect 11529 13209 11563 13243
rect 17509 13209 17543 13243
rect 18061 13209 18095 13243
rect 19809 13209 19843 13243
rect 20269 13209 20303 13243
rect 23213 13209 23247 13243
rect 31953 13209 31987 13243
rect 32045 13209 32079 13243
rect 33057 13209 33091 13243
rect 39037 13209 39071 13243
rect 4905 13141 4939 13175
rect 5457 13141 5491 13175
rect 7757 13141 7791 13175
rect 8493 13141 8527 13175
rect 10333 13141 10367 13175
rect 13553 13141 13587 13175
rect 15025 13141 15059 13175
rect 16405 13141 16439 13175
rect 21557 13141 21591 13175
rect 23013 13141 23047 13175
rect 32505 13141 32539 13175
rect 38577 13141 38611 13175
rect 39497 13141 39531 13175
rect 5181 12937 5215 12971
rect 8493 12937 8527 12971
rect 10609 12937 10643 12971
rect 11897 12937 11931 12971
rect 12541 12937 12575 12971
rect 13185 12937 13219 12971
rect 17509 12937 17543 12971
rect 21005 12937 21039 12971
rect 26985 12937 27019 12971
rect 28917 12937 28951 12971
rect 29101 12937 29135 12971
rect 31217 12937 31251 12971
rect 32689 12937 32723 12971
rect 35449 12937 35483 12971
rect 7389 12869 7423 12903
rect 21833 12869 21867 12903
rect 23397 12869 23431 12903
rect 27353 12869 27387 12903
rect 35173 12869 35207 12903
rect 2145 12801 2179 12835
rect 4353 12801 4387 12835
rect 4445 12801 4479 12835
rect 4629 12801 4663 12835
rect 4721 12801 4755 12835
rect 5456 12801 5490 12835
rect 5549 12801 5583 12835
rect 5641 12801 5675 12835
rect 7113 12801 7147 12835
rect 7665 12801 7699 12835
rect 7757 12801 7791 12835
rect 7849 12801 7883 12835
rect 8033 12801 8067 12835
rect 8309 12801 8343 12835
rect 8585 12801 8619 12835
rect 10793 12801 10827 12835
rect 10885 12801 10919 12835
rect 11253 12801 11287 12835
rect 11713 12801 11747 12835
rect 11989 12801 12023 12835
rect 12909 12801 12943 12835
rect 13277 12801 13311 12835
rect 13737 12801 13771 12835
rect 14105 12801 14139 12835
rect 14565 12801 14599 12835
rect 14749 12801 14783 12835
rect 16957 12801 16991 12835
rect 17417 12801 17451 12835
rect 17693 12801 17727 12835
rect 17785 12801 17819 12835
rect 17969 12801 18003 12835
rect 18061 12801 18095 12835
rect 18521 12801 18555 12835
rect 18981 12801 19015 12835
rect 21189 12801 21223 12835
rect 21557 12801 21591 12835
rect 22109 12801 22143 12835
rect 22293 12801 22327 12835
rect 22385 12801 22419 12835
rect 22569 12801 22603 12835
rect 22845 12801 22879 12835
rect 23213 12801 23247 12835
rect 23857 12801 23891 12835
rect 23949 12801 23983 12835
rect 24133 12801 24167 12835
rect 24593 12801 24627 12835
rect 24685 12801 24719 12835
rect 25053 12801 25087 12835
rect 25329 12801 25363 12835
rect 25605 12801 25639 12835
rect 27169 12801 27203 12835
rect 27261 12801 27295 12835
rect 27537 12801 27571 12835
rect 27629 12801 27663 12835
rect 28089 12801 28123 12835
rect 28181 12801 28215 12835
rect 28365 12801 28399 12835
rect 28549 12801 28583 12835
rect 28733 12801 28767 12835
rect 29009 12801 29043 12835
rect 29193 12801 29227 12835
rect 30021 12801 30055 12835
rect 30205 12801 30239 12835
rect 30481 12801 30515 12835
rect 30573 12801 30607 12835
rect 30757 12801 30791 12835
rect 30849 12801 30883 12835
rect 31033 12801 31067 12835
rect 31131 12801 31165 12835
rect 31309 12801 31343 12835
rect 32137 12801 32171 12835
rect 32321 12801 32355 12835
rect 32413 12801 32447 12835
rect 32505 12801 32539 12835
rect 34805 12801 34839 12835
rect 34898 12801 34932 12835
rect 35081 12801 35115 12835
rect 35270 12801 35304 12835
rect 38669 12801 38703 12835
rect 38945 12801 38979 12835
rect 2421 12733 2455 12767
rect 4169 12733 4203 12767
rect 5733 12733 5767 12767
rect 6745 12733 6779 12767
rect 7021 12733 7055 12767
rect 11161 12733 11195 12767
rect 17141 12733 17175 12767
rect 18705 12733 18739 12767
rect 23121 12733 23155 12767
rect 24777 12733 24811 12767
rect 25421 12733 25455 12767
rect 29745 12733 29779 12767
rect 30941 12733 30975 12767
rect 38761 12733 38795 12767
rect 11529 12665 11563 12699
rect 12817 12665 12851 12699
rect 14289 12665 14323 12699
rect 22661 12665 22695 12699
rect 24041 12665 24075 12699
rect 24317 12665 24351 12699
rect 28273 12665 28307 12699
rect 3893 12597 3927 12631
rect 5825 12597 5859 12631
rect 6009 12597 6043 12631
rect 8125 12597 8159 12631
rect 13001 12597 13035 12631
rect 14105 12597 14139 12631
rect 14473 12597 14507 12631
rect 16681 12597 16715 12631
rect 17049 12597 17083 12631
rect 17233 12597 17267 12631
rect 18337 12597 18371 12631
rect 18889 12597 18923 12631
rect 21465 12597 21499 12631
rect 22201 12597 22235 12631
rect 23029 12597 23063 12631
rect 23673 12597 23707 12631
rect 24869 12597 24903 12631
rect 25145 12597 25179 12631
rect 25605 12597 25639 12631
rect 27905 12597 27939 12631
rect 30113 12597 30147 12631
rect 30297 12597 30331 12631
rect 30757 12597 30791 12631
rect 38945 12597 38979 12631
rect 39129 12597 39163 12631
rect 4445 12393 4479 12427
rect 6377 12393 6411 12427
rect 7021 12393 7055 12427
rect 7665 12393 7699 12427
rect 13001 12393 13035 12427
rect 17969 12393 18003 12427
rect 19349 12393 19383 12427
rect 19533 12393 19567 12427
rect 19809 12393 19843 12427
rect 20177 12393 20211 12427
rect 20269 12393 20303 12427
rect 26249 12393 26283 12427
rect 30113 12393 30147 12427
rect 30757 12393 30791 12427
rect 33425 12393 33459 12427
rect 35357 12393 35391 12427
rect 38117 12393 38151 12427
rect 38577 12393 38611 12427
rect 4353 12325 4387 12359
rect 27905 12325 27939 12359
rect 4077 12257 4111 12291
rect 4813 12257 4847 12291
rect 6101 12257 6135 12291
rect 6561 12257 6595 12291
rect 7205 12257 7239 12291
rect 16773 12257 16807 12291
rect 20361 12257 20395 12291
rect 33793 12257 33827 12291
rect 34713 12257 34747 12291
rect 38301 12257 38335 12291
rect 3985 12189 4019 12223
rect 4629 12189 4663 12223
rect 5641 12189 5675 12223
rect 6193 12189 6227 12223
rect 6653 12189 6687 12223
rect 6929 12189 6963 12223
rect 7573 12189 7607 12223
rect 7757 12189 7791 12223
rect 12817 12189 12851 12223
rect 12910 12189 12944 12223
rect 14105 12189 14139 12223
rect 14749 12189 14783 12223
rect 14841 12189 14875 12223
rect 15209 12189 15243 12223
rect 17049 12189 17083 12223
rect 17509 12189 17543 12223
rect 17877 12189 17911 12223
rect 18153 12189 18187 12223
rect 18613 12189 18647 12223
rect 18797 12189 18831 12223
rect 18981 12189 19015 12223
rect 20085 12189 20119 12223
rect 20545 12189 20579 12223
rect 20637 12189 20671 12223
rect 26065 12189 26099 12223
rect 26249 12189 26283 12223
rect 27905 12189 27939 12223
rect 28089 12189 28123 12223
rect 29929 12189 29963 12223
rect 30113 12189 30147 12223
rect 30665 12189 30699 12223
rect 30757 12189 30791 12223
rect 33149 12189 33183 12223
rect 33609 12189 33643 12223
rect 34871 12189 34905 12223
rect 35173 12189 35207 12223
rect 35725 12189 35759 12223
rect 38393 12189 38427 12223
rect 5733 12121 5767 12155
rect 5825 12121 5859 12155
rect 5943 12121 5977 12155
rect 15025 12121 15059 12155
rect 15117 12121 15151 12155
rect 18337 12121 18371 12155
rect 19717 12121 19751 12155
rect 34989 12121 35023 12155
rect 35081 12121 35115 12155
rect 38117 12121 38151 12155
rect 5457 12053 5491 12087
rect 6837 12053 6871 12087
rect 7481 12053 7515 12087
rect 15393 12053 15427 12087
rect 19533 12053 19567 12087
rect 20821 12053 20855 12087
rect 35541 12053 35575 12087
rect 5273 11849 5307 11883
rect 6377 11849 6411 11883
rect 15669 11849 15703 11883
rect 16865 11849 16899 11883
rect 17233 11849 17267 11883
rect 25513 11849 25547 11883
rect 37105 11849 37139 11883
rect 38485 11849 38519 11883
rect 3801 11781 3835 11815
rect 8861 11781 8895 11815
rect 9505 11781 9539 11815
rect 15209 11781 15243 11815
rect 24041 11781 24075 11815
rect 25881 11781 25915 11815
rect 26065 11781 26099 11815
rect 33333 11781 33367 11815
rect 34687 11781 34721 11815
rect 34897 11781 34931 11815
rect 39037 11781 39071 11815
rect 6652 11713 6686 11747
rect 6745 11713 6779 11747
rect 8493 11713 8527 11747
rect 8586 11713 8620 11747
rect 8769 11713 8803 11747
rect 8999 11713 9033 11747
rect 10057 11713 10091 11747
rect 10150 11713 10184 11747
rect 13093 11713 13127 11747
rect 15485 11713 15519 11747
rect 15761 11713 15795 11747
rect 15945 11713 15979 11747
rect 17049 11713 17083 11747
rect 17325 11713 17359 11747
rect 20085 11713 20119 11747
rect 20177 11713 20211 11747
rect 20361 11713 20395 11747
rect 20545 11713 20579 11747
rect 20821 11713 20855 11747
rect 21097 11713 21131 11747
rect 24133 11713 24167 11747
rect 24501 11713 24535 11747
rect 24961 11713 24995 11747
rect 25145 11713 25179 11747
rect 25237 11713 25271 11747
rect 25513 11713 25547 11747
rect 25697 11713 25731 11747
rect 26157 11713 26191 11747
rect 26433 11713 26467 11747
rect 26617 11713 26651 11747
rect 26709 11713 26743 11747
rect 28641 11713 28675 11747
rect 32505 11713 32539 11747
rect 33609 11713 33643 11747
rect 34805 11713 34839 11747
rect 34989 11713 35023 11747
rect 36461 11713 36495 11747
rect 36554 11713 36588 11747
rect 36737 11713 36771 11747
rect 36829 11713 36863 11747
rect 36926 11713 36960 11747
rect 38025 11713 38059 11747
rect 38301 11713 38335 11747
rect 38761 11713 38795 11747
rect 3525 11645 3559 11679
rect 9965 11645 9999 11679
rect 13185 11645 13219 11679
rect 13737 11645 13771 11679
rect 21005 11645 21039 11679
rect 23213 11645 23247 11679
rect 24685 11645 24719 11679
rect 28549 11645 28583 11679
rect 31677 11645 31711 11679
rect 31953 11645 31987 11679
rect 34529 11645 34563 11679
rect 38117 11645 38151 11679
rect 38945 11645 38979 11679
rect 9781 11577 9815 11611
rect 20269 11577 20303 11611
rect 20637 11577 20671 11611
rect 25053 11577 25087 11611
rect 26433 11577 26467 11611
rect 28273 11577 28307 11611
rect 9137 11509 9171 11543
rect 10241 11509 10275 11543
rect 13461 11509 13495 11543
rect 19901 11509 19935 11543
rect 24225 11509 24259 11543
rect 24777 11509 24811 11543
rect 25881 11509 25915 11543
rect 28641 11509 28675 11543
rect 33701 11509 33735 11543
rect 35173 11509 35207 11543
rect 38025 11509 38059 11543
rect 38577 11509 38611 11543
rect 39037 11509 39071 11543
rect 8677 11305 8711 11339
rect 14197 11305 14231 11339
rect 17325 11305 17359 11339
rect 17601 11305 17635 11339
rect 18245 11305 18279 11339
rect 19901 11305 19935 11339
rect 21741 11305 21775 11339
rect 24409 11305 24443 11339
rect 24593 11305 24627 11339
rect 27077 11305 27111 11339
rect 27997 11305 28031 11339
rect 28089 11305 28123 11339
rect 28457 11305 28491 11339
rect 29561 11305 29595 11339
rect 37197 11305 37231 11339
rect 8125 11237 8159 11271
rect 10241 11237 10275 11271
rect 11713 11237 11747 11271
rect 12265 11237 12299 11271
rect 17141 11237 17175 11271
rect 20085 11237 20119 11271
rect 8769 11169 8803 11203
rect 9045 11169 9079 11203
rect 11069 11169 11103 11203
rect 15485 11169 15519 11203
rect 20269 11169 20303 11203
rect 20361 11169 20395 11203
rect 22293 11169 22327 11203
rect 24685 11169 24719 11203
rect 27537 11169 27571 11203
rect 33149 11169 33183 11203
rect 33241 11169 33275 11203
rect 33333 11169 33367 11203
rect 36277 11169 36311 11203
rect 37105 11169 37139 11203
rect 2053 11101 2087 11135
rect 7849 11101 7883 11135
rect 8033 11101 8067 11135
rect 8306 11101 8340 11135
rect 8953 11101 8987 11135
rect 9137 11101 9171 11135
rect 9781 11101 9815 11135
rect 9873 11101 9907 11135
rect 10057 11101 10091 11135
rect 10149 11101 10183 11135
rect 10420 11101 10454 11135
rect 10517 11101 10551 11135
rect 10737 11101 10771 11135
rect 10885 11101 10919 11135
rect 11161 11101 11195 11135
rect 11345 11101 11379 11135
rect 11529 11101 11563 11135
rect 11805 11101 11839 11135
rect 11989 11101 12023 11135
rect 12403 11101 12437 11135
rect 12541 11101 12575 11135
rect 12633 11101 12667 11135
rect 12816 11101 12850 11135
rect 12909 11101 12943 11135
rect 13001 11101 13035 11135
rect 14105 11101 14139 11135
rect 14289 11101 14323 11135
rect 15669 11101 15703 11135
rect 17785 11101 17819 11135
rect 17877 11101 17911 11135
rect 18061 11101 18095 11135
rect 18153 11101 18187 11135
rect 18245 11101 18279 11135
rect 18521 11101 18555 11135
rect 20545 11101 20579 11135
rect 20729 11101 20763 11135
rect 21557 11101 21591 11135
rect 21741 11101 21775 11135
rect 22477 11101 22511 11135
rect 22661 11101 22695 11135
rect 22937 11101 22971 11135
rect 23213 11101 23247 11135
rect 24777 11101 24811 11135
rect 25881 11101 25915 11135
rect 26157 11101 26191 11135
rect 26801 11101 26835 11135
rect 26893 11101 26927 11135
rect 27813 11101 27847 11135
rect 27905 11101 27939 11135
rect 28273 11101 28307 11135
rect 28457 11101 28491 11135
rect 28733 11101 28767 11135
rect 29009 11101 29043 11135
rect 29193 11101 29227 11135
rect 29561 11101 29595 11135
rect 29745 11101 29779 11135
rect 29837 11101 29871 11135
rect 30573 11101 30607 11135
rect 31769 11101 31803 11135
rect 32045 11101 32079 11135
rect 32873 11101 32907 11135
rect 33425 11101 33459 11135
rect 33701 11101 33735 11135
rect 33859 11101 33893 11135
rect 34069 11101 34103 11135
rect 34161 11101 34195 11135
rect 34345 11101 34379 11135
rect 34897 11101 34931 11135
rect 34989 11101 35023 11135
rect 35265 11101 35299 11135
rect 36415 11101 36449 11135
rect 36645 11101 36679 11135
rect 36737 11101 36771 11135
rect 37289 11101 37323 11135
rect 7941 11033 7975 11067
rect 9597 11033 9631 11067
rect 10609 11033 10643 11067
rect 13093 11033 13127 11067
rect 17309 11033 17343 11067
rect 17509 11033 17543 11067
rect 19717 11033 19751 11067
rect 19933 11033 19967 11067
rect 21281 11033 21315 11067
rect 27077 11033 27111 11067
rect 28641 11033 28675 11067
rect 30297 11033 30331 11067
rect 33977 11033 34011 11067
rect 35081 11033 35115 11067
rect 36553 11033 36587 11067
rect 36921 11033 36955 11067
rect 37013 11033 37047 11067
rect 1869 10965 1903 10999
rect 8309 10965 8343 10999
rect 11897 10965 11931 10999
rect 18429 10965 18463 10999
rect 21925 10965 21959 10999
rect 25973 10965 26007 10999
rect 29285 10965 29319 10999
rect 32965 10965 32999 10999
rect 34713 10965 34747 10999
rect 37473 10965 37507 10999
rect 7389 10761 7423 10795
rect 10149 10761 10183 10795
rect 14473 10761 14507 10795
rect 16957 10761 16991 10795
rect 22569 10761 22603 10795
rect 23121 10761 23155 10795
rect 24041 10761 24075 10795
rect 26065 10761 26099 10795
rect 28089 10761 28123 10795
rect 30665 10761 30699 10795
rect 31217 10761 31251 10795
rect 31769 10761 31803 10795
rect 32873 10761 32907 10795
rect 6653 10693 6687 10727
rect 7573 10693 7607 10727
rect 8401 10693 8435 10727
rect 8601 10693 8635 10727
rect 8953 10693 8987 10727
rect 9137 10693 9171 10727
rect 9597 10693 9631 10727
rect 12725 10693 12759 10727
rect 24225 10693 24259 10727
rect 24409 10693 24443 10727
rect 25421 10693 25455 10727
rect 26249 10693 26283 10727
rect 29653 10693 29687 10727
rect 32413 10693 32447 10727
rect 32505 10693 32539 10727
rect 37289 10693 37323 10727
rect 38853 10693 38887 10727
rect 6561 10625 6595 10659
rect 6745 10625 6779 10659
rect 6929 10625 6963 10659
rect 7205 10625 7239 10659
rect 7481 10625 7515 10659
rect 7757 10625 7791 10659
rect 8033 10625 8067 10659
rect 8217 10625 8251 10659
rect 8861 10625 8895 10659
rect 9872 10625 9906 10659
rect 9965 10625 9999 10659
rect 10057 10625 10091 10659
rect 10241 10625 10275 10659
rect 12449 10625 12483 10659
rect 12633 10625 12667 10659
rect 12817 10625 12851 10659
rect 14841 10625 14875 10659
rect 14933 10625 14967 10659
rect 15117 10625 15151 10659
rect 16957 10625 16991 10659
rect 17141 10625 17175 10659
rect 21005 10625 21039 10659
rect 21189 10625 21223 10659
rect 21281 10625 21315 10659
rect 21373 10625 21407 10659
rect 21833 10625 21867 10659
rect 22017 10625 22051 10659
rect 23029 10625 23063 10659
rect 23305 10625 23339 10659
rect 23489 10625 23523 10659
rect 25789 10625 25823 10659
rect 27537 10625 27571 10659
rect 27721 10625 27755 10659
rect 27813 10625 27847 10659
rect 27905 10625 27939 10659
rect 28181 10625 28215 10659
rect 28365 10625 28399 10659
rect 29837 10625 29871 10659
rect 30297 10625 30331 10659
rect 30849 10625 30883 10659
rect 31401 10625 31435 10659
rect 31953 10625 31987 10659
rect 32321 10625 32355 10659
rect 32689 10625 32723 10659
rect 32781 10625 32815 10659
rect 33057 10625 33091 10659
rect 33333 10625 33367 10659
rect 37565 10625 37599 10659
rect 38301 10625 38335 10659
rect 38485 10625 38519 10659
rect 39037 10625 39071 10659
rect 14749 10557 14783 10591
rect 22293 10557 22327 10591
rect 24685 10557 24719 10591
rect 31033 10557 31067 10591
rect 31585 10557 31619 10591
rect 33149 10557 33183 10591
rect 33241 10557 33275 10591
rect 37473 10557 37507 10591
rect 21649 10489 21683 10523
rect 22201 10489 22235 10523
rect 28365 10489 28399 10523
rect 6377 10421 6411 10455
rect 7021 10421 7055 10455
rect 7941 10421 7975 10455
rect 8125 10421 8159 10455
rect 8585 10421 8619 10455
rect 8769 10421 8803 10455
rect 9137 10421 9171 10455
rect 13001 10421 13035 10455
rect 14749 10421 14783 10455
rect 15117 10421 15151 10455
rect 22109 10421 22143 10455
rect 24225 10421 24259 10455
rect 26065 10421 26099 10455
rect 32137 10421 32171 10455
rect 37289 10421 37323 10455
rect 37749 10421 37783 10455
rect 38485 10421 38519 10455
rect 38669 10421 38703 10455
rect 39221 10421 39255 10455
rect 4248 10217 4282 10251
rect 10149 10217 10183 10251
rect 12633 10217 12667 10251
rect 14473 10217 14507 10251
rect 14933 10217 14967 10251
rect 16865 10217 16899 10251
rect 18705 10217 18739 10251
rect 19073 10217 19107 10251
rect 19533 10217 19567 10251
rect 25697 10217 25731 10251
rect 26709 10217 26743 10251
rect 28549 10217 28583 10251
rect 30849 10217 30883 10251
rect 32321 10217 32355 10251
rect 32781 10217 32815 10251
rect 36737 10217 36771 10251
rect 5733 10149 5767 10183
rect 19717 10149 19751 10183
rect 28917 10149 28951 10183
rect 29009 10149 29043 10183
rect 32505 10149 32539 10183
rect 32965 10149 32999 10183
rect 3985 10081 4019 10115
rect 7297 10081 7331 10115
rect 9965 10081 9999 10115
rect 15117 10081 15151 10115
rect 18981 10081 19015 10115
rect 19349 10081 19383 10115
rect 29377 10081 29411 10115
rect 29653 10081 29687 10115
rect 36921 10081 36955 10115
rect 39681 10081 39715 10115
rect 6101 10013 6135 10047
rect 7113 10013 7147 10047
rect 7389 10013 7423 10047
rect 7481 10013 7515 10047
rect 7573 10013 7607 10047
rect 7757 10013 7791 10047
rect 7849 10013 7883 10047
rect 8309 10013 8343 10047
rect 8953 10013 8987 10047
rect 10241 10013 10275 10047
rect 11345 10013 11379 10047
rect 11529 10013 11563 10047
rect 12725 10013 12759 10047
rect 12909 10013 12943 10047
rect 14657 10013 14691 10047
rect 17233 10013 17267 10047
rect 17601 10013 17635 10047
rect 17693 10013 17727 10047
rect 17877 10013 17911 10047
rect 17969 10013 18003 10047
rect 19073 10013 19107 10047
rect 19533 10013 19567 10047
rect 19993 10013 20027 10047
rect 20085 10013 20119 10047
rect 24869 10013 24903 10047
rect 25329 10013 25363 10047
rect 25605 10013 25639 10047
rect 25973 10013 26007 10047
rect 26065 10013 26099 10047
rect 26341 10013 26375 10047
rect 26433 10013 26467 10047
rect 26525 10013 26559 10047
rect 26709 10013 26743 10047
rect 27721 10013 27755 10047
rect 28089 10013 28123 10047
rect 28457 10013 28491 10047
rect 28733 10013 28767 10047
rect 29837 10013 29871 10047
rect 30021 10013 30055 10047
rect 30573 10013 30607 10047
rect 30665 10013 30699 10047
rect 31125 10013 31159 10047
rect 32597 10013 32631 10047
rect 32781 10013 32815 10047
rect 37013 10013 37047 10047
rect 37841 10013 37875 10047
rect 6837 9945 6871 9979
rect 9689 9945 9723 9979
rect 12265 9945 12299 9979
rect 12449 9945 12483 9979
rect 14749 9945 14783 9979
rect 15393 9945 15427 9979
rect 17325 9945 17359 9979
rect 17417 9945 17451 9979
rect 19257 9945 19291 9979
rect 19809 9945 19843 9979
rect 25513 9945 25547 9979
rect 32137 9945 32171 9979
rect 32353 9945 32387 9979
rect 35633 9945 35667 9979
rect 36737 9945 36771 9979
rect 39405 9945 39439 9979
rect 7205 9877 7239 9911
rect 7665 9877 7699 9911
rect 9965 9877 9999 9911
rect 11437 9877 11471 9911
rect 12817 9877 12851 9911
rect 17049 9877 17083 9911
rect 25145 9877 25179 9911
rect 26157 9877 26191 9911
rect 27905 9877 27939 9911
rect 28273 9877 28307 9911
rect 30941 9877 30975 9911
rect 35725 9877 35759 9911
rect 37197 9877 37231 9911
rect 37657 9877 37691 9911
rect 37933 9877 37967 9911
rect 8217 9673 8251 9707
rect 8953 9673 8987 9707
rect 12541 9673 12575 9707
rect 14473 9673 14507 9707
rect 15669 9673 15703 9707
rect 22661 9673 22695 9707
rect 24317 9673 24351 9707
rect 25329 9673 25363 9707
rect 28641 9673 28675 9707
rect 30849 9673 30883 9707
rect 34897 9673 34931 9707
rect 36737 9673 36771 9707
rect 9321 9605 9355 9639
rect 9505 9605 9539 9639
rect 9689 9605 9723 9639
rect 10701 9605 10735 9639
rect 11897 9605 11931 9639
rect 12449 9605 12483 9639
rect 14565 9605 14599 9639
rect 14765 9605 14799 9639
rect 16221 9605 16255 9639
rect 24961 9605 24995 9639
rect 25161 9605 25195 9639
rect 26985 9605 27019 9639
rect 29193 9605 29227 9639
rect 29837 9605 29871 9639
rect 31401 9605 31435 9639
rect 34621 9605 34655 9639
rect 35219 9605 35253 9639
rect 35449 9605 35483 9639
rect 35725 9605 35759 9639
rect 36093 9605 36127 9639
rect 36185 9605 36219 9639
rect 37749 9605 37783 9639
rect 38025 9605 38059 9639
rect 38301 9605 38335 9639
rect 6837 9537 6871 9571
rect 7021 9537 7055 9571
rect 7205 9537 7239 9571
rect 8125 9537 8159 9571
rect 8381 9537 8415 9571
rect 9137 9537 9171 9571
rect 9413 9537 9447 9571
rect 9781 9537 9815 9571
rect 11069 9537 11103 9571
rect 11161 9537 11195 9571
rect 11713 9537 11747 9571
rect 11989 9537 12023 9571
rect 13277 9537 13311 9571
rect 13461 9537 13495 9571
rect 14289 9537 14323 9571
rect 14473 9537 14507 9571
rect 15117 9537 15151 9571
rect 15209 9537 15243 9571
rect 15393 9537 15427 9571
rect 15485 9537 15519 9571
rect 15945 9537 15979 9571
rect 16037 9537 16071 9571
rect 18153 9537 18187 9571
rect 18337 9537 18371 9571
rect 20545 9537 20579 9571
rect 20729 9537 20763 9571
rect 22109 9537 22143 9571
rect 22385 9537 22419 9571
rect 22845 9537 22879 9571
rect 23029 9537 23063 9571
rect 24133 9537 24167 9571
rect 27813 9537 27847 9571
rect 28825 9537 28859 9571
rect 31033 9537 31067 9571
rect 31125 9537 31159 9571
rect 31217 9537 31251 9571
rect 32137 9537 32171 9571
rect 32321 9537 32355 9571
rect 32505 9537 32539 9571
rect 32689 9537 32723 9571
rect 32873 9537 32907 9571
rect 34253 9537 34287 9571
rect 34401 9537 34435 9571
rect 34529 9537 34563 9571
rect 34718 9537 34752 9571
rect 35081 9537 35115 9571
rect 35357 9537 35391 9571
rect 35541 9537 35575 9571
rect 35975 9537 36009 9571
rect 36277 9537 36311 9571
rect 36645 9537 36679 9571
rect 37657 9537 37691 9571
rect 37841 9537 37875 9571
rect 38669 9537 38703 9571
rect 10793 9469 10827 9503
rect 12357 9469 12391 9503
rect 13185 9469 13219 9503
rect 13369 9469 13403 9503
rect 16221 9469 16255 9503
rect 18429 9469 18463 9503
rect 22201 9469 22235 9503
rect 27353 9469 27387 9503
rect 27905 9469 27939 9503
rect 30205 9469 30239 9503
rect 35817 9469 35851 9503
rect 36461 9469 36495 9503
rect 11345 9401 11379 9435
rect 13001 9401 13035 9435
rect 14933 9401 14967 9435
rect 30297 9401 30331 9435
rect 30757 9401 30791 9435
rect 37473 9401 37507 9435
rect 38485 9401 38519 9435
rect 7389 9333 7423 9367
rect 8585 9333 8619 9367
rect 9597 9333 9631 9367
rect 11529 9333 11563 9367
rect 12909 9333 12943 9367
rect 14749 9333 14783 9367
rect 17969 9333 18003 9367
rect 20637 9333 20671 9367
rect 20913 9333 20947 9367
rect 22385 9333 22419 9367
rect 22569 9333 22603 9367
rect 22845 9333 22879 9367
rect 25145 9333 25179 9367
rect 27445 9333 27479 9367
rect 29101 9333 29135 9367
rect 30389 9333 30423 9367
rect 38209 9333 38243 9367
rect 12817 9129 12851 9163
rect 20361 9129 20395 9163
rect 20545 9129 20579 9163
rect 21005 9129 21039 9163
rect 22293 9129 22327 9163
rect 22477 9129 22511 9163
rect 24041 9129 24075 9163
rect 24593 9129 24627 9163
rect 25053 9129 25087 9163
rect 25513 9129 25547 9163
rect 26525 9129 26559 9163
rect 26893 9129 26927 9163
rect 26985 9129 27019 9163
rect 27721 9129 27755 9163
rect 31493 9129 31527 9163
rect 35541 9129 35575 9163
rect 37381 9129 37415 9163
rect 37657 9129 37691 9163
rect 37841 9129 37875 9163
rect 7941 9061 7975 9095
rect 28917 9061 28951 9095
rect 11897 8993 11931 9027
rect 15485 8993 15519 9027
rect 26801 8993 26835 9027
rect 29101 8993 29135 9027
rect 32965 8993 32999 9027
rect 38301 8993 38335 9027
rect 6929 8925 6963 8959
rect 7297 8925 7331 8959
rect 7481 8925 7515 8959
rect 7665 8925 7699 8959
rect 7757 8925 7791 8959
rect 8217 8925 8251 8959
rect 8401 8925 8435 8959
rect 10517 8925 10551 8959
rect 10609 8925 10643 8959
rect 10701 8925 10735 8959
rect 10885 8925 10919 8959
rect 11161 8925 11195 8959
rect 11437 8925 11471 8959
rect 11713 8925 11747 8959
rect 12173 8925 12207 8959
rect 12357 8925 12391 8959
rect 12449 8925 12483 8959
rect 14565 8925 14599 8959
rect 14749 8925 14783 8959
rect 17693 8925 17727 8959
rect 17877 8925 17911 8959
rect 17969 8925 18003 8959
rect 24225 8925 24259 8959
rect 26157 8925 26191 8959
rect 26341 8925 26375 8959
rect 27353 8925 27387 8959
rect 27629 8925 27663 8959
rect 28273 8925 28307 8959
rect 28733 8925 28767 8959
rect 29009 8925 29043 8959
rect 29285 8925 29319 8959
rect 29745 8925 29779 8959
rect 30113 8925 30147 8959
rect 30665 8925 30699 8959
rect 30849 8925 30883 8959
rect 31125 8925 31159 8959
rect 31309 8925 31343 8959
rect 32781 8925 32815 8959
rect 35725 8925 35759 8959
rect 37197 8925 37231 8959
rect 37381 8925 37415 8959
rect 37933 8925 37967 8959
rect 37703 8891 37737 8925
rect 7021 8857 7055 8891
rect 7205 8857 7239 8891
rect 7941 8857 7975 8891
rect 8309 8857 8343 8891
rect 11345 8857 11379 8891
rect 11529 8857 11563 8891
rect 11989 8857 12023 8891
rect 12633 8857 12667 8891
rect 20513 8857 20547 8891
rect 20729 8857 20763 8891
rect 20973 8857 21007 8891
rect 21189 8857 21223 8891
rect 22661 8857 22695 8891
rect 24409 8857 24443 8891
rect 24625 8857 24659 8891
rect 24869 8857 24903 8891
rect 25329 8857 25363 8891
rect 25545 8857 25579 8891
rect 26249 8857 26283 8891
rect 29561 8857 29595 8891
rect 30389 8857 30423 8891
rect 33333 8857 33367 8891
rect 33517 8857 33551 8891
rect 37473 8857 37507 8891
rect 38485 8857 38519 8891
rect 6929 8789 6963 8823
rect 7389 8789 7423 8823
rect 10333 8789 10367 8823
rect 10977 8789 11011 8823
rect 20821 8789 20855 8823
rect 22461 8789 22495 8823
rect 24777 8789 24811 8823
rect 25074 8789 25108 8823
rect 25237 8789 25271 8823
rect 25697 8789 25731 8823
rect 33425 8789 33459 8823
rect 38117 8789 38151 8823
rect 4261 8585 4295 8619
rect 7205 8585 7239 8619
rect 8953 8585 8987 8619
rect 15853 8585 15887 8619
rect 23121 8585 23155 8619
rect 23397 8585 23431 8619
rect 27077 8585 27111 8619
rect 28181 8585 28215 8619
rect 28641 8585 28675 8619
rect 28733 8585 28767 8619
rect 33793 8585 33827 8619
rect 34253 8585 34287 8619
rect 34529 8585 34563 8619
rect 36093 8585 36127 8619
rect 36185 8585 36219 8619
rect 37933 8585 37967 8619
rect 14841 8517 14875 8551
rect 20177 8517 20211 8551
rect 21833 8517 21867 8551
rect 22043 8517 22077 8551
rect 23565 8517 23599 8551
rect 23765 8517 23799 8551
rect 24133 8517 24167 8551
rect 24225 8517 24259 8551
rect 24777 8517 24811 8551
rect 34621 8517 34655 8551
rect 36645 8517 36679 8551
rect 38761 8517 38795 8551
rect 6009 8449 6043 8483
rect 6653 8449 6687 8483
rect 6837 8449 6871 8483
rect 6929 8449 6963 8483
rect 7389 8449 7423 8483
rect 7481 8449 7515 8483
rect 7573 8449 7607 8483
rect 7757 8449 7791 8483
rect 7849 8449 7883 8483
rect 8217 8449 8251 8483
rect 8401 8449 8435 8483
rect 8769 8449 8803 8483
rect 9045 8449 9079 8483
rect 10333 8449 10367 8483
rect 10517 8449 10551 8483
rect 10609 8449 10643 8483
rect 10885 8449 10919 8483
rect 11897 8449 11931 8483
rect 12357 8449 12391 8483
rect 15209 8449 15243 8483
rect 15301 8449 15335 8483
rect 15485 8449 15519 8483
rect 15577 8449 15611 8483
rect 15669 8449 15703 8483
rect 17601 8449 17635 8483
rect 18613 8449 18647 8483
rect 18705 8449 18739 8483
rect 18889 8449 18923 8483
rect 19073 8449 19107 8483
rect 19625 8449 19659 8483
rect 19901 8449 19935 8483
rect 20085 8449 20119 8483
rect 20453 8449 20487 8483
rect 20545 8449 20579 8483
rect 20637 8449 20671 8483
rect 20821 8449 20855 8483
rect 21373 8449 21407 8483
rect 23305 8449 23339 8483
rect 24041 8449 24075 8483
rect 24409 8449 24443 8483
rect 24869 8449 24903 8483
rect 25237 8449 25271 8483
rect 25697 8449 25731 8483
rect 25973 8449 26007 8483
rect 26709 8449 26743 8483
rect 27261 8449 27295 8483
rect 27629 8449 27663 8483
rect 27905 8449 27939 8483
rect 28273 8449 28307 8483
rect 28365 8449 28399 8483
rect 28917 8449 28951 8483
rect 29193 8449 29227 8483
rect 29653 8449 29687 8483
rect 29745 8449 29779 8483
rect 30665 8449 30699 8483
rect 32321 8449 32355 8483
rect 32597 8449 32631 8483
rect 35909 8449 35943 8483
rect 37749 8449 37783 8483
rect 5733 8381 5767 8415
rect 6745 8381 6779 8415
rect 7941 8381 7975 8415
rect 8125 8381 8159 8415
rect 8300 8381 8334 8415
rect 11529 8381 11563 8415
rect 13369 8381 13403 8415
rect 15117 8381 15151 8415
rect 17693 8381 17727 8415
rect 17877 8381 17911 8415
rect 19809 8381 19843 8415
rect 27721 8381 27755 8415
rect 30021 8381 30055 8415
rect 33333 8381 33367 8415
rect 34412 8381 34446 8415
rect 34897 8381 34931 8415
rect 38485 8381 38519 8415
rect 40233 8381 40267 8415
rect 8585 8313 8619 8347
rect 10425 8313 10459 8347
rect 10701 8313 10735 8347
rect 11069 8313 11103 8347
rect 18797 8313 18831 8347
rect 19349 8313 19383 8347
rect 22201 8313 22235 8347
rect 29009 8313 29043 8347
rect 29101 8313 29135 8347
rect 33701 8313 33735 8347
rect 36645 8313 36679 8347
rect 6469 8245 6503 8279
rect 17233 8245 17267 8279
rect 18429 8245 18463 8279
rect 19717 8245 19751 8279
rect 21281 8245 21315 8279
rect 22017 8245 22051 8279
rect 23581 8245 23615 8279
rect 23857 8245 23891 8279
rect 27261 8245 27295 8279
rect 27997 8245 28031 8279
rect 29469 8245 29503 8279
rect 32137 8245 32171 8279
rect 32413 8245 32447 8279
rect 5181 8041 5215 8075
rect 11253 8041 11287 8075
rect 14565 8041 14599 8075
rect 15301 8041 15335 8075
rect 18797 8041 18831 8075
rect 19441 8041 19475 8075
rect 23397 8041 23431 8075
rect 24685 8041 24719 8075
rect 25513 8041 25547 8075
rect 26341 8041 26375 8075
rect 27261 8041 27295 8075
rect 28273 8041 28307 8075
rect 28641 8041 28675 8075
rect 30205 8041 30239 8075
rect 30389 8041 30423 8075
rect 30849 8041 30883 8075
rect 36553 8041 36587 8075
rect 7113 7973 7147 8007
rect 7849 7973 7883 8007
rect 8033 7973 8067 8007
rect 11161 7973 11195 8007
rect 15117 7973 15151 8007
rect 20269 7973 20303 8007
rect 25237 7973 25271 8007
rect 25973 7973 26007 8007
rect 26801 7973 26835 8007
rect 28457 7973 28491 8007
rect 5641 7905 5675 7939
rect 5825 7905 5859 7939
rect 6837 7905 6871 7939
rect 7389 7905 7423 7939
rect 7941 7905 7975 7939
rect 8217 7905 8251 7939
rect 8401 7905 8435 7939
rect 9781 7905 9815 7939
rect 9873 7905 9907 7939
rect 9965 7905 9999 7939
rect 10793 7905 10827 7939
rect 16037 7905 16071 7939
rect 20913 7905 20947 7939
rect 23029 7905 23063 7939
rect 25605 7905 25639 7939
rect 26249 7905 26283 7939
rect 27077 7905 27111 7939
rect 31401 7905 31435 7939
rect 31493 7905 31527 7939
rect 32413 7905 32447 7939
rect 32597 7905 32631 7939
rect 33333 7905 33367 7939
rect 33517 7905 33551 7939
rect 34897 7905 34931 7939
rect 35817 7905 35851 7939
rect 36737 7905 36771 7939
rect 5549 7837 5583 7871
rect 6745 7837 6779 7871
rect 7297 7837 7331 7871
rect 7481 7837 7515 7871
rect 7573 7837 7607 7871
rect 7849 7837 7883 7871
rect 8493 7837 8527 7871
rect 9689 7837 9723 7871
rect 13921 7837 13955 7871
rect 14105 7837 14139 7871
rect 14381 7837 14415 7871
rect 14565 7837 14599 7871
rect 14841 7837 14875 7871
rect 15577 7837 15611 7871
rect 15669 7837 15703 7871
rect 15853 7837 15887 7871
rect 15945 7837 15979 7871
rect 18705 7837 18739 7871
rect 18889 7837 18923 7871
rect 19257 7837 19291 7871
rect 19441 7837 19475 7871
rect 20177 7837 20211 7871
rect 20361 7837 20395 7871
rect 20453 7837 20487 7871
rect 21189 7837 21223 7871
rect 22109 7837 22143 7871
rect 22201 7837 22235 7871
rect 22293 7837 22327 7871
rect 22385 7837 22419 7871
rect 22569 7837 22603 7871
rect 22753 7837 22787 7871
rect 22937 7837 22971 7871
rect 23121 7837 23155 7871
rect 23213 7837 23247 7871
rect 24133 7837 24167 7871
rect 25881 7837 25915 7871
rect 26341 7837 26375 7871
rect 26985 7837 27019 7871
rect 27261 7837 27295 7871
rect 28733 7837 28767 7871
rect 28825 7837 28859 7871
rect 29193 7837 29227 7871
rect 29377 7837 29411 7871
rect 29745 7837 29779 7871
rect 29837 7837 29871 7871
rect 30205 7837 30239 7871
rect 30573 7837 30607 7871
rect 30849 7837 30883 7871
rect 31217 7837 31251 7871
rect 31861 7837 31895 7871
rect 31953 7837 31987 7871
rect 32965 7837 32999 7871
rect 33977 7837 34011 7871
rect 35265 7837 35299 7871
rect 35357 7837 35391 7871
rect 40141 7837 40175 7871
rect 7757 7769 7791 7803
rect 8309 7769 8343 7803
rect 15393 7769 15427 7803
rect 16313 7769 16347 7803
rect 18061 7769 18095 7803
rect 24961 7769 24995 7803
rect 28089 7769 28123 7803
rect 32045 7769 32079 7803
rect 33149 7769 33183 7803
rect 34069 7769 34103 7803
rect 34805 7769 34839 7803
rect 36461 7769 36495 7803
rect 37013 7769 37047 7803
rect 38761 7769 38795 7803
rect 9505 7701 9539 7735
rect 13829 7701 13863 7735
rect 14197 7701 14231 7735
rect 19993 7701 20027 7735
rect 21925 7701 21959 7735
rect 24041 7701 24075 7735
rect 24869 7701 24903 7735
rect 25053 7701 25087 7735
rect 25329 7701 25363 7735
rect 28289 7701 28323 7735
rect 31033 7701 31067 7735
rect 33057 7701 33091 7735
rect 33885 7701 33919 7735
rect 39957 7701 39991 7735
rect 8033 7497 8067 7531
rect 12081 7497 12115 7531
rect 14473 7497 14507 7531
rect 16773 7497 16807 7531
rect 17509 7497 17543 7531
rect 17969 7497 18003 7531
rect 18137 7497 18171 7531
rect 22017 7497 22051 7531
rect 22185 7497 22219 7531
rect 24961 7497 24995 7531
rect 25053 7497 25087 7531
rect 27445 7497 27479 7531
rect 29653 7497 29687 7531
rect 31309 7497 31343 7531
rect 32413 7497 32447 7531
rect 33885 7497 33919 7531
rect 37381 7497 37415 7531
rect 40049 7497 40083 7531
rect 9505 7429 9539 7463
rect 15117 7429 15151 7463
rect 16497 7429 16531 7463
rect 17325 7429 17359 7463
rect 18337 7429 18371 7463
rect 21649 7429 21683 7463
rect 22385 7429 22419 7463
rect 26249 7429 26283 7463
rect 29561 7429 29595 7463
rect 31125 7429 31159 7463
rect 38577 7429 38611 7463
rect 21419 7395 21453 7429
rect 8217 7361 8251 7395
rect 8309 7361 8343 7395
rect 9229 7361 9263 7395
rect 11989 7361 12023 7395
rect 12449 7361 12483 7395
rect 12725 7361 12759 7395
rect 14749 7361 14783 7395
rect 15301 7361 15335 7395
rect 15393 7361 15427 7395
rect 16681 7361 16715 7395
rect 16865 7361 16899 7395
rect 18429 7361 18463 7395
rect 21005 7361 21039 7395
rect 21097 7361 21131 7395
rect 24409 7361 24443 7395
rect 25605 7361 25639 7395
rect 26525 7361 26559 7395
rect 26617 7361 26651 7395
rect 26985 7361 27019 7395
rect 27353 7361 27387 7395
rect 27537 7361 27571 7395
rect 27813 7361 27847 7395
rect 31217 7361 31251 7395
rect 32781 7361 32815 7395
rect 33793 7361 33827 7395
rect 33977 7361 34011 7395
rect 34345 7361 34379 7395
rect 34529 7361 34563 7395
rect 35265 7361 35299 7395
rect 35449 7361 35483 7395
rect 35817 7361 35851 7395
rect 37289 7361 37323 7395
rect 37473 7361 37507 7395
rect 38301 7361 38335 7395
rect 10977 7293 11011 7327
rect 13001 7293 13035 7327
rect 15025 7293 15059 7327
rect 15117 7293 15151 7327
rect 15761 7293 15795 7327
rect 18521 7293 18555 7327
rect 20821 7293 20855 7327
rect 20913 7293 20947 7327
rect 24685 7293 24719 7327
rect 25329 7293 25363 7327
rect 26433 7293 26467 7327
rect 26709 7293 26743 7327
rect 31585 7293 31619 7327
rect 32296 7293 32330 7327
rect 32505 7293 32539 7327
rect 35173 7293 35207 7327
rect 16957 7225 16991 7259
rect 20637 7225 20671 7259
rect 34897 7225 34931 7259
rect 12541 7157 12575 7191
rect 14565 7157 14599 7191
rect 14933 7157 14967 7191
rect 17325 7157 17359 7191
rect 18153 7157 18187 7191
rect 18429 7157 18463 7191
rect 18797 7157 18831 7191
rect 21281 7157 21315 7191
rect 21465 7157 21499 7191
rect 22201 7157 22235 7191
rect 24777 7157 24811 7191
rect 25237 7157 25271 7191
rect 30941 7157 30975 7191
rect 32137 7157 32171 7191
rect 12357 6953 12391 6987
rect 13277 6953 13311 6987
rect 36369 6953 36403 6987
rect 37853 6953 37887 6987
rect 14197 6885 14231 6919
rect 15669 6885 15703 6919
rect 21189 6885 21223 6919
rect 30389 6885 30423 6919
rect 33977 6885 34011 6919
rect 11621 6817 11655 6851
rect 12173 6817 12207 6851
rect 13461 6817 13495 6851
rect 13553 6817 13587 6851
rect 14933 6817 14967 6851
rect 17233 6817 17267 6851
rect 17417 6817 17451 6851
rect 33793 6817 33827 6851
rect 38117 6817 38151 6851
rect 11529 6749 11563 6783
rect 11805 6749 11839 6783
rect 12357 6749 12391 6783
rect 13645 6749 13679 6783
rect 13737 6749 13771 6783
rect 14749 6749 14783 6783
rect 15485 6749 15519 6783
rect 15669 6749 15703 6783
rect 20913 6749 20947 6783
rect 29561 6749 29595 6783
rect 29929 6749 29963 6783
rect 30205 6749 30239 6783
rect 34253 6749 34287 6783
rect 11897 6681 11931 6715
rect 12081 6681 12115 6715
rect 14197 6681 14231 6715
rect 15778 6681 15812 6715
rect 29745 6681 29779 6715
rect 29837 6681 29871 6715
rect 12541 6613 12575 6647
rect 14657 6613 14691 6647
rect 16773 6613 16807 6647
rect 17141 6613 17175 6647
rect 30113 6613 30147 6647
rect 11897 6409 11931 6443
rect 16405 6409 16439 6443
rect 17877 6409 17911 6443
rect 21465 6409 21499 6443
rect 26617 6409 26651 6443
rect 29469 6409 29503 6443
rect 19349 6341 19383 6375
rect 27629 6341 27663 6375
rect 30941 6341 30975 6375
rect 11989 6273 12023 6307
rect 12357 6273 12391 6307
rect 14657 6273 14691 6307
rect 24961 6273 24995 6307
rect 26801 6273 26835 6307
rect 27169 6273 27203 6307
rect 27261 6273 27295 6307
rect 27353 6273 27387 6307
rect 27537 6273 27571 6307
rect 27997 6273 28031 6307
rect 31217 6273 31251 6307
rect 12173 6205 12207 6239
rect 12909 6205 12943 6239
rect 14933 6205 14967 6239
rect 19625 6205 19659 6239
rect 19717 6205 19751 6239
rect 19993 6205 20027 6239
rect 22845 6205 22879 6239
rect 22477 6137 22511 6171
rect 11529 6069 11563 6103
rect 22385 6069 22419 6103
rect 25145 6069 25179 6103
rect 26985 6069 27019 6103
rect 19993 5865 20027 5899
rect 20453 5865 20487 5899
rect 28733 5865 28767 5899
rect 29561 5865 29595 5899
rect 19073 5797 19107 5831
rect 29377 5797 29411 5831
rect 10425 5729 10459 5763
rect 17693 5729 17727 5763
rect 19717 5729 19751 5763
rect 20913 5729 20947 5763
rect 22201 5729 22235 5763
rect 24225 5729 24259 5763
rect 26985 5729 27019 5763
rect 27261 5729 27295 5763
rect 31033 5729 31067 5763
rect 31309 5729 31343 5763
rect 18521 5661 18555 5695
rect 18797 5661 18831 5695
rect 19349 5661 19383 5695
rect 19533 5661 19567 5695
rect 19625 5661 19659 5695
rect 19809 5661 19843 5695
rect 20085 5661 20119 5695
rect 20269 5661 20303 5695
rect 20453 5661 20487 5695
rect 20545 5661 20579 5695
rect 21097 5661 21131 5695
rect 21373 5661 21407 5695
rect 21557 5661 21591 5695
rect 21649 5661 21683 5695
rect 21833 5661 21867 5695
rect 24501 5661 24535 5695
rect 24869 5661 24903 5695
rect 25329 5661 25363 5695
rect 25697 5661 25731 5695
rect 25789 5661 25823 5695
rect 26249 5661 26283 5695
rect 26617 5661 26651 5695
rect 28825 5661 28859 5695
rect 29101 5661 29135 5695
rect 29193 5661 29227 5695
rect 10701 5593 10735 5627
rect 17417 5593 17451 5627
rect 19073 5593 19107 5627
rect 20637 5593 20671 5627
rect 22477 5593 22511 5627
rect 24685 5593 24719 5627
rect 24777 5593 24811 5627
rect 25421 5593 25455 5627
rect 25513 5593 25547 5627
rect 26433 5593 26467 5627
rect 26525 5593 26559 5627
rect 29009 5593 29043 5627
rect 12173 5525 12207 5559
rect 17049 5525 17083 5559
rect 17509 5525 17543 5559
rect 17969 5525 18003 5559
rect 18889 5525 18923 5559
rect 19441 5525 19475 5559
rect 21833 5525 21867 5559
rect 25053 5525 25087 5559
rect 25145 5525 25179 5559
rect 25973 5525 26007 5559
rect 26801 5525 26835 5559
rect 13553 5321 13587 5355
rect 18429 5321 18463 5355
rect 21373 5321 21407 5355
rect 22569 5321 22603 5355
rect 23581 5321 23615 5355
rect 26985 5321 27019 5355
rect 30297 5321 30331 5355
rect 16957 5253 16991 5287
rect 22937 5253 22971 5287
rect 24961 5253 24995 5287
rect 11805 5185 11839 5219
rect 18521 5185 18555 5219
rect 18797 5185 18831 5219
rect 19349 5185 19383 5219
rect 20361 5185 20395 5219
rect 20729 5185 20763 5219
rect 21281 5185 21315 5219
rect 21465 5185 21499 5219
rect 22753 5185 22787 5219
rect 22845 5185 22879 5219
rect 23121 5185 23155 5219
rect 23213 5185 23247 5219
rect 23397 5185 23431 5219
rect 24685 5185 24719 5219
rect 28733 5185 28767 5219
rect 29009 5185 29043 5219
rect 29193 5185 29227 5219
rect 30205 5185 30239 5219
rect 12081 5117 12115 5151
rect 13645 5117 13679 5151
rect 13921 5117 13955 5151
rect 16037 5117 16071 5151
rect 16681 5117 16715 5151
rect 22385 5117 22419 5151
rect 26709 5117 26743 5151
rect 28457 5117 28491 5151
rect 15485 5049 15519 5083
rect 19073 5049 19107 5083
rect 20545 5049 20579 5083
rect 15393 4981 15427 5015
rect 18613 4981 18647 5015
rect 19993 4981 20027 5015
rect 20269 4981 20303 5015
rect 20913 4981 20947 5015
rect 21833 4981 21867 5015
rect 28825 4981 28859 5015
rect 12357 4777 12391 4811
rect 14289 4777 14323 4811
rect 19073 4777 19107 4811
rect 21189 4777 21223 4811
rect 13001 4641 13035 4675
rect 14749 4641 14783 4675
rect 14841 4641 14875 4675
rect 15301 4641 15335 4675
rect 15577 4641 15611 4675
rect 19257 4641 19291 4675
rect 19533 4641 19567 4675
rect 21005 4641 21039 4675
rect 22937 4641 22971 4675
rect 24777 4641 24811 4675
rect 12265 4573 12299 4607
rect 12725 4573 12759 4607
rect 13829 4573 13863 4607
rect 17325 4573 17359 4607
rect 26801 4573 26835 4607
rect 14657 4505 14691 4539
rect 17601 4505 17635 4539
rect 22661 4505 22695 4539
rect 25053 4505 25087 4539
rect 11621 4437 11655 4471
rect 12817 4437 12851 4471
rect 13185 4437 13219 4471
rect 17049 4437 17083 4471
rect 11989 4233 12023 4267
rect 12725 4233 12759 4267
rect 16221 4233 16255 4267
rect 21097 4233 21131 4267
rect 22661 4233 22695 4267
rect 11897 4165 11931 4199
rect 16129 4165 16163 4199
rect 19809 4165 19843 4199
rect 20269 4165 20303 4199
rect 21281 4165 21315 4199
rect 21373 4165 21407 4199
rect 12817 4097 12851 4131
rect 14105 4097 14139 4131
rect 16681 4097 16715 4131
rect 18521 4097 18555 4131
rect 18705 4097 18739 4131
rect 18981 4097 19015 4131
rect 19717 4097 19751 4131
rect 19993 4097 20027 4131
rect 20085 4097 20119 4131
rect 21005 4097 21039 4131
rect 21557 4097 21591 4131
rect 21649 4097 21683 4131
rect 23121 4097 23155 4131
rect 23213 4097 23247 4131
rect 23305 4097 23339 4131
rect 23489 4097 23523 4131
rect 28181 4097 28215 4131
rect 28549 4097 28583 4131
rect 12173 4029 12207 4063
rect 13001 4029 13035 4063
rect 13921 4029 13955 4063
rect 14657 4029 14691 4063
rect 15761 4029 15795 4063
rect 17693 4029 17727 4063
rect 18337 4029 18371 4063
rect 18613 4029 18647 4063
rect 18797 4029 18831 4063
rect 19073 4029 19107 4063
rect 22017 4029 22051 4063
rect 22845 4029 22879 4063
rect 19809 3961 19843 3995
rect 21281 3961 21315 3995
rect 29929 3961 29963 3995
rect 11529 3893 11563 3927
rect 12357 3893 12391 3927
rect 13369 3893 13403 3927
rect 15209 3893 15243 3927
rect 16773 3893 16807 3927
rect 17141 3893 17175 3927
rect 20361 3893 20395 3927
rect 21373 3893 21407 3927
rect 12449 3689 12483 3723
rect 19901 3689 19935 3723
rect 21649 3689 21683 3723
rect 22740 3689 22774 3723
rect 39957 3621 39991 3655
rect 10701 3553 10735 3587
rect 13001 3553 13035 3587
rect 13139 3553 13173 3587
rect 14841 3553 14875 3587
rect 15025 3553 15059 3587
rect 17325 3553 17359 3587
rect 17969 3553 18003 3587
rect 22477 3553 22511 3587
rect 26157 3553 26191 3587
rect 12909 3485 12943 3519
rect 13737 3485 13771 3519
rect 14749 3485 14783 3519
rect 15577 3485 15611 3519
rect 19257 3485 19291 3519
rect 21373 3485 21407 3519
rect 22201 3485 22235 3519
rect 26801 3485 26835 3519
rect 10977 3417 11011 3451
rect 13369 3417 13403 3451
rect 15853 3417 15887 3451
rect 21465 3417 21499 3451
rect 25881 3417 25915 3451
rect 26249 3417 26283 3451
rect 40141 3417 40175 3451
rect 12541 3349 12575 3383
rect 14381 3349 14415 3383
rect 17417 3349 17451 3383
rect 24225 3349 24259 3383
rect 24409 3349 24443 3383
rect 17049 3145 17083 3179
rect 17141 3145 17175 3179
rect 21649 3145 21683 3179
rect 22753 3145 22787 3179
rect 25789 3145 25823 3179
rect 12265 3077 12299 3111
rect 14105 3077 14139 3111
rect 15761 3077 15795 3111
rect 23949 3077 23983 3111
rect 24501 3077 24535 3111
rect 11621 3009 11655 3043
rect 13829 3009 13863 3043
rect 15669 3009 15703 3043
rect 18061 3009 18095 3043
rect 19901 3009 19935 3043
rect 21833 3009 21867 3043
rect 22569 3009 22603 3043
rect 22845 3009 22879 3043
rect 23213 3009 23247 3043
rect 24317 3009 24351 3043
rect 24593 3009 24627 3043
rect 11989 2941 12023 2975
rect 17325 2941 17359 2975
rect 18337 2941 18371 2975
rect 20177 2941 20211 2975
rect 22201 2941 22235 2975
rect 23489 2941 23523 2975
rect 25329 2941 25363 2975
rect 13737 2873 13771 2907
rect 15577 2873 15611 2907
rect 16681 2873 16715 2907
rect 25237 2873 25271 2907
rect 25605 2873 25639 2907
rect 11805 2805 11839 2839
rect 19809 2805 19843 2839
rect 18889 2601 18923 2635
rect 19349 2601 19383 2635
rect 20637 2601 20671 2635
rect 13461 2533 13495 2567
rect 15485 2533 15519 2567
rect 21189 2533 21223 2567
rect 11529 2465 11563 2499
rect 13277 2465 13311 2499
rect 17141 2465 17175 2499
rect 17417 2465 17451 2499
rect 19993 2465 20027 2499
rect 23213 2465 23247 2499
rect 11345 2397 11379 2431
rect 13645 2397 13679 2431
rect 14289 2397 14323 2431
rect 15209 2397 15243 2431
rect 15301 2397 15335 2431
rect 16221 2397 16255 2431
rect 17049 2397 17083 2431
rect 19441 2397 19475 2431
rect 21005 2397 21039 2431
rect 21373 2397 21407 2431
rect 23397 2397 23431 2431
rect 11805 2329 11839 2363
rect 21097 2329 21131 2363
rect 21281 2329 21315 2363
rect 11161 2261 11195 2295
rect 14473 2261 14507 2295
rect 15025 2261 15059 2295
rect 16405 2261 16439 2295
rect 16865 2261 16899 2295
rect 21557 2261 21591 2295
rect 23581 2261 23615 2295
<< metal1 >>
rect 1104 41370 40572 41392
rect 1104 41318 4874 41370
rect 4926 41318 4938 41370
rect 4990 41318 5002 41370
rect 5054 41318 5066 41370
rect 5118 41318 5130 41370
rect 5182 41318 35594 41370
rect 35646 41318 35658 41370
rect 35710 41318 35722 41370
rect 35774 41318 35786 41370
rect 35838 41318 35850 41370
rect 35902 41318 40572 41370
rect 1104 41296 40572 41318
rect 30926 41080 30932 41132
rect 30984 41120 30990 41132
rect 31021 41123 31079 41129
rect 31021 41120 31033 41123
rect 30984 41092 31033 41120
rect 30984 41080 30990 41092
rect 31021 41089 31033 41092
rect 31067 41089 31079 41123
rect 31021 41083 31079 41089
rect 31202 41012 31208 41064
rect 31260 41012 31266 41064
rect 1104 40826 40572 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 40572 40826
rect 1104 40752 40572 40774
rect 16301 40647 16359 40653
rect 16301 40613 16313 40647
rect 16347 40644 16359 40647
rect 17034 40644 17040 40656
rect 16347 40616 17040 40644
rect 16347 40613 16359 40616
rect 16301 40607 16359 40613
rect 17034 40604 17040 40616
rect 17092 40604 17098 40656
rect 15010 40536 15016 40588
rect 15068 40576 15074 40588
rect 15841 40579 15899 40585
rect 15841 40576 15853 40579
rect 15068 40548 15853 40576
rect 15068 40536 15074 40548
rect 15841 40545 15853 40548
rect 15887 40545 15899 40579
rect 15841 40539 15899 40545
rect 15746 40468 15752 40520
rect 15804 40468 15810 40520
rect 16025 40511 16083 40517
rect 16025 40477 16037 40511
rect 16071 40508 16083 40511
rect 16390 40508 16396 40520
rect 16071 40480 16396 40508
rect 16071 40477 16083 40480
rect 16025 40471 16083 40477
rect 16390 40468 16396 40480
rect 16448 40468 16454 40520
rect 16574 40468 16580 40520
rect 16632 40468 16638 40520
rect 16301 40443 16359 40449
rect 16301 40409 16313 40443
rect 16347 40409 16359 40443
rect 16301 40403 16359 40409
rect 15930 40332 15936 40384
rect 15988 40372 15994 40384
rect 16209 40375 16267 40381
rect 16209 40372 16221 40375
rect 15988 40344 16221 40372
rect 15988 40332 15994 40344
rect 16209 40341 16221 40344
rect 16255 40372 16267 40375
rect 16316 40372 16344 40403
rect 16255 40344 16344 40372
rect 16255 40341 16267 40344
rect 16209 40335 16267 40341
rect 16482 40332 16488 40384
rect 16540 40332 16546 40384
rect 1104 40282 40572 40304
rect 1104 40230 4874 40282
rect 4926 40230 4938 40282
rect 4990 40230 5002 40282
rect 5054 40230 5066 40282
rect 5118 40230 5130 40282
rect 5182 40230 35594 40282
rect 35646 40230 35658 40282
rect 35710 40230 35722 40282
rect 35774 40230 35786 40282
rect 35838 40230 35850 40282
rect 35902 40230 40572 40282
rect 1104 40208 40572 40230
rect 13534 40171 13592 40177
rect 13534 40137 13546 40171
rect 13580 40168 13592 40171
rect 15470 40168 15476 40180
rect 13580 40140 13860 40168
rect 13580 40137 13592 40140
rect 13534 40131 13592 40137
rect 13446 40100 13452 40112
rect 11992 40072 13452 40100
rect 11992 40041 12020 40072
rect 13446 40060 13452 40072
rect 13504 40060 13510 40112
rect 13832 40100 13860 40140
rect 14844 40140 15476 40168
rect 14844 40100 14872 40140
rect 15470 40128 15476 40140
rect 15528 40128 15534 40180
rect 13832 40072 13952 40100
rect 11977 40035 12035 40041
rect 11977 40001 11989 40035
rect 12023 40001 12035 40035
rect 11977 39995 12035 40001
rect 13357 40035 13415 40041
rect 13357 40001 13369 40035
rect 13403 40001 13415 40035
rect 13357 39995 13415 40001
rect 12069 39967 12127 39973
rect 12069 39933 12081 39967
rect 12115 39964 12127 39967
rect 12250 39964 12256 39976
rect 12115 39936 12256 39964
rect 12115 39933 12127 39936
rect 12069 39927 12127 39933
rect 12250 39924 12256 39936
rect 12308 39924 12314 39976
rect 12158 39788 12164 39840
rect 12216 39828 12222 39840
rect 12345 39831 12403 39837
rect 12345 39828 12357 39831
rect 12216 39800 12357 39828
rect 12216 39788 12222 39800
rect 12345 39797 12357 39800
rect 12391 39797 12403 39831
rect 12345 39791 12403 39797
rect 12526 39788 12532 39840
rect 12584 39828 12590 39840
rect 13372 39828 13400 39995
rect 13630 39992 13636 40044
rect 13688 39992 13694 40044
rect 13924 40041 13952 40072
rect 14752 40072 14872 40100
rect 15289 40103 15347 40109
rect 14752 40041 14780 40072
rect 15289 40069 15301 40103
rect 15335 40100 15347 40103
rect 15335 40072 16436 40100
rect 15335 40069 15347 40072
rect 15289 40063 15347 40069
rect 13909 40035 13967 40041
rect 13909 40001 13921 40035
rect 13955 40001 13967 40035
rect 13909 39995 13967 40001
rect 14737 40035 14795 40041
rect 14737 40001 14749 40035
rect 14783 40001 14795 40035
rect 14737 39995 14795 40001
rect 15010 39992 15016 40044
rect 15068 39992 15074 40044
rect 14001 39967 14059 39973
rect 14001 39933 14013 39967
rect 14047 39964 14059 39967
rect 14369 39967 14427 39973
rect 14369 39964 14381 39967
rect 14047 39936 14381 39964
rect 14047 39933 14059 39936
rect 14001 39927 14059 39933
rect 14369 39933 14381 39936
rect 14415 39964 14427 39967
rect 14458 39964 14464 39976
rect 14415 39936 14464 39964
rect 14415 39933 14427 39936
rect 14369 39927 14427 39933
rect 14458 39924 14464 39936
rect 14516 39924 14522 39976
rect 15396 39973 15424 40072
rect 16408 40044 16436 40072
rect 15562 39992 15568 40044
rect 15620 40032 15626 40044
rect 15749 40035 15807 40041
rect 15749 40032 15761 40035
rect 15620 40004 15761 40032
rect 15620 39992 15626 40004
rect 15749 40001 15761 40004
rect 15795 40001 15807 40035
rect 15749 39995 15807 40001
rect 16209 40035 16267 40041
rect 16209 40001 16221 40035
rect 16255 40001 16267 40035
rect 16209 39995 16267 40001
rect 14645 39967 14703 39973
rect 14645 39933 14657 39967
rect 14691 39933 14703 39967
rect 14645 39927 14703 39933
rect 15381 39967 15439 39973
rect 15381 39933 15393 39967
rect 15427 39933 15439 39967
rect 15381 39927 15439 39933
rect 15841 39967 15899 39973
rect 15841 39933 15853 39967
rect 15887 39964 15899 39967
rect 16224 39964 16252 39995
rect 16390 39992 16396 40044
rect 16448 40032 16454 40044
rect 16669 40035 16727 40041
rect 16669 40032 16681 40035
rect 16448 40004 16681 40032
rect 16448 39992 16454 40004
rect 16669 40001 16681 40004
rect 16715 40001 16727 40035
rect 16669 39995 16727 40001
rect 16853 40035 16911 40041
rect 16853 40001 16865 40035
rect 16899 40032 16911 40035
rect 17126 40032 17132 40044
rect 16899 40004 17132 40032
rect 16899 40001 16911 40004
rect 16853 39995 16911 40001
rect 17126 39992 17132 40004
rect 17184 39992 17190 40044
rect 15887 39936 16252 39964
rect 15887 39933 15899 39936
rect 15841 39927 15899 39933
rect 14274 39856 14280 39908
rect 14332 39856 14338 39908
rect 14660 39828 14688 39927
rect 15105 39899 15163 39905
rect 15105 39865 15117 39899
rect 15151 39896 15163 39899
rect 15746 39896 15752 39908
rect 15151 39868 15752 39896
rect 15151 39865 15163 39868
rect 15105 39859 15163 39865
rect 15746 39856 15752 39868
rect 15804 39896 15810 39908
rect 16025 39899 16083 39905
rect 16025 39896 16037 39899
rect 15804 39868 16037 39896
rect 15804 39856 15810 39868
rect 16025 39865 16037 39868
rect 16071 39865 16083 39899
rect 16224 39896 16252 39936
rect 16298 39924 16304 39976
rect 16356 39964 16362 39976
rect 16485 39967 16543 39973
rect 16485 39964 16497 39967
rect 16356 39936 16497 39964
rect 16356 39924 16362 39936
rect 16485 39933 16497 39936
rect 16531 39933 16543 39967
rect 16485 39927 16543 39933
rect 16850 39896 16856 39908
rect 16224 39868 16856 39896
rect 16025 39859 16083 39865
rect 16850 39856 16856 39868
rect 16908 39896 16914 39908
rect 17862 39896 17868 39908
rect 16908 39868 17868 39896
rect 16908 39856 16914 39868
rect 17862 39856 17868 39868
rect 17920 39856 17926 39908
rect 12584 39800 14688 39828
rect 12584 39788 12590 39800
rect 15194 39788 15200 39840
rect 15252 39788 15258 39840
rect 16390 39788 16396 39840
rect 16448 39788 16454 39840
rect 16942 39788 16948 39840
rect 17000 39828 17006 39840
rect 17037 39831 17095 39837
rect 17037 39828 17049 39831
rect 17000 39800 17049 39828
rect 17000 39788 17006 39800
rect 17037 39797 17049 39800
rect 17083 39797 17095 39831
rect 17037 39791 17095 39797
rect 1104 39738 40572 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 40572 39738
rect 1104 39664 40572 39686
rect 11974 39624 11980 39636
rect 11440 39596 11980 39624
rect 8297 39491 8355 39497
rect 8297 39457 8309 39491
rect 8343 39488 8355 39491
rect 8478 39488 8484 39500
rect 8343 39460 8484 39488
rect 8343 39457 8355 39460
rect 8297 39451 8355 39457
rect 8478 39448 8484 39460
rect 8536 39488 8542 39500
rect 8536 39460 11284 39488
rect 8536 39448 8542 39460
rect 11256 39432 11284 39460
rect 8386 39380 8392 39432
rect 8444 39420 8450 39432
rect 8573 39423 8631 39429
rect 8573 39420 8585 39423
rect 8444 39392 8585 39420
rect 8444 39380 8450 39392
rect 8573 39389 8585 39392
rect 8619 39389 8631 39423
rect 8573 39383 8631 39389
rect 8757 39423 8815 39429
rect 8757 39389 8769 39423
rect 8803 39420 8815 39423
rect 9398 39420 9404 39432
rect 8803 39392 9404 39420
rect 8803 39389 8815 39392
rect 8757 39383 8815 39389
rect 9398 39380 9404 39392
rect 9456 39380 9462 39432
rect 11238 39380 11244 39432
rect 11296 39380 11302 39432
rect 11440 39429 11468 39596
rect 11974 39584 11980 39596
rect 12032 39584 12038 39636
rect 12345 39627 12403 39633
rect 12345 39593 12357 39627
rect 12391 39624 12403 39627
rect 12391 39596 13032 39624
rect 12391 39593 12403 39596
rect 12345 39587 12403 39593
rect 12066 39556 12072 39568
rect 11900 39528 12072 39556
rect 11900 39497 11928 39528
rect 12066 39516 12072 39528
rect 12124 39556 12130 39568
rect 12529 39559 12587 39565
rect 12529 39556 12541 39559
rect 12124 39528 12541 39556
rect 12124 39516 12130 39528
rect 12529 39525 12541 39528
rect 12575 39525 12587 39559
rect 12529 39519 12587 39525
rect 11885 39491 11943 39497
rect 11885 39488 11897 39491
rect 11716 39460 11897 39488
rect 11425 39423 11483 39429
rect 11425 39389 11437 39423
rect 11471 39389 11483 39423
rect 11425 39383 11483 39389
rect 11514 39380 11520 39432
rect 11572 39380 11578 39432
rect 11716 39429 11744 39460
rect 11885 39457 11897 39460
rect 11931 39457 11943 39491
rect 12713 39491 12771 39497
rect 12713 39488 12725 39491
rect 11885 39451 11943 39457
rect 12176 39460 12725 39488
rect 12176 39432 12204 39460
rect 12713 39457 12725 39460
rect 12759 39457 12771 39491
rect 12713 39451 12771 39457
rect 11701 39423 11759 39429
rect 11701 39389 11713 39423
rect 11747 39389 11759 39423
rect 11701 39383 11759 39389
rect 12158 39380 12164 39432
rect 12216 39380 12222 39432
rect 13004 39429 13032 39596
rect 15286 39584 15292 39636
rect 15344 39624 15350 39636
rect 16209 39627 16267 39633
rect 16209 39624 16221 39627
rect 15344 39596 16221 39624
rect 15344 39584 15350 39596
rect 16209 39593 16221 39596
rect 16255 39624 16267 39627
rect 16390 39624 16396 39636
rect 16255 39596 16396 39624
rect 16255 39593 16267 39596
rect 16209 39587 16267 39593
rect 16390 39584 16396 39596
rect 16448 39584 16454 39636
rect 15562 39516 15568 39568
rect 15620 39556 15626 39568
rect 16117 39559 16175 39565
rect 16117 39556 16129 39559
rect 15620 39528 16129 39556
rect 15620 39516 15626 39528
rect 16117 39525 16129 39528
rect 16163 39556 16175 39559
rect 16482 39556 16488 39568
rect 16163 39528 16488 39556
rect 16163 39525 16175 39528
rect 16117 39519 16175 39525
rect 16482 39516 16488 39528
rect 16540 39516 16546 39568
rect 13630 39448 13636 39500
rect 13688 39488 13694 39500
rect 14277 39491 14335 39497
rect 14277 39488 14289 39491
rect 13688 39460 14289 39488
rect 13688 39448 13694 39460
rect 14277 39457 14289 39460
rect 14323 39457 14335 39491
rect 15930 39488 15936 39500
rect 14277 39451 14335 39457
rect 15764 39460 15936 39488
rect 12437 39423 12495 39429
rect 12437 39420 12449 39423
rect 12268 39392 12449 39420
rect 8294 39244 8300 39296
rect 8352 39284 8358 39296
rect 8481 39287 8539 39293
rect 8481 39284 8493 39287
rect 8352 39256 8493 39284
rect 8352 39244 8358 39256
rect 8481 39253 8493 39256
rect 8527 39253 8539 39287
rect 8481 39247 8539 39253
rect 11054 39244 11060 39296
rect 11112 39284 11118 39296
rect 11333 39287 11391 39293
rect 11333 39284 11345 39287
rect 11112 39256 11345 39284
rect 11112 39244 11118 39256
rect 11333 39253 11345 39256
rect 11379 39253 11391 39287
rect 11333 39247 11391 39253
rect 11606 39244 11612 39296
rect 11664 39244 11670 39296
rect 11974 39244 11980 39296
rect 12032 39284 12038 39296
rect 12268 39284 12296 39392
rect 12437 39389 12449 39392
rect 12483 39389 12495 39423
rect 12437 39383 12495 39389
rect 12805 39423 12863 39429
rect 12805 39389 12817 39423
rect 12851 39389 12863 39423
rect 12805 39383 12863 39389
rect 12989 39423 13047 39429
rect 12989 39389 13001 39423
rect 13035 39420 13047 39423
rect 13648 39420 13676 39448
rect 13035 39392 13676 39420
rect 13035 39389 13047 39392
rect 12989 39383 13047 39389
rect 12032 39256 12296 39284
rect 12437 39287 12495 39293
rect 12032 39244 12038 39256
rect 12437 39253 12449 39287
rect 12483 39284 12495 39287
rect 12820 39284 12848 39383
rect 14458 39380 14464 39432
rect 14516 39380 14522 39432
rect 15194 39380 15200 39432
rect 15252 39420 15258 39432
rect 15764 39429 15792 39460
rect 15930 39448 15936 39460
rect 15988 39448 15994 39500
rect 17034 39448 17040 39500
rect 17092 39448 17098 39500
rect 17589 39491 17647 39497
rect 17589 39457 17601 39491
rect 17635 39457 17647 39491
rect 17589 39451 17647 39457
rect 15565 39423 15623 39429
rect 15565 39420 15577 39423
rect 15252 39392 15577 39420
rect 15252 39380 15258 39392
rect 15565 39389 15577 39392
rect 15611 39389 15623 39423
rect 15565 39383 15623 39389
rect 15749 39423 15807 39429
rect 15749 39389 15761 39423
rect 15795 39389 15807 39423
rect 15749 39383 15807 39389
rect 15838 39380 15844 39432
rect 15896 39380 15902 39432
rect 16025 39423 16083 39429
rect 16025 39389 16037 39423
rect 16071 39420 16083 39423
rect 16206 39420 16212 39432
rect 16071 39392 16212 39420
rect 16071 39389 16083 39392
rect 16025 39383 16083 39389
rect 15470 39312 15476 39364
rect 15528 39352 15534 39364
rect 16040 39352 16068 39383
rect 16206 39380 16212 39392
rect 16264 39380 16270 39432
rect 16301 39423 16359 39429
rect 16301 39389 16313 39423
rect 16347 39420 16359 39423
rect 16574 39420 16580 39432
rect 16347 39392 16580 39420
rect 16347 39389 16359 39392
rect 16301 39383 16359 39389
rect 16574 39380 16580 39392
rect 16632 39380 16638 39432
rect 17126 39380 17132 39432
rect 17184 39420 17190 39432
rect 17604 39420 17632 39451
rect 17862 39448 17868 39500
rect 17920 39488 17926 39500
rect 18049 39491 18107 39497
rect 18049 39488 18061 39491
rect 17920 39460 18061 39488
rect 17920 39448 17926 39460
rect 18049 39457 18061 39460
rect 18095 39457 18107 39491
rect 18049 39451 18107 39457
rect 17184 39392 17632 39420
rect 17957 39423 18015 39429
rect 17184 39380 17190 39392
rect 17957 39389 17969 39423
rect 18003 39389 18015 39423
rect 17957 39383 18015 39389
rect 17972 39352 18000 39383
rect 18046 39352 18052 39364
rect 15528 39324 16068 39352
rect 16500 39324 18052 39352
rect 15528 39312 15534 39324
rect 12483 39256 12848 39284
rect 12897 39287 12955 39293
rect 12483 39253 12495 39256
rect 12437 39247 12495 39253
rect 12897 39253 12909 39287
rect 12943 39284 12955 39287
rect 12986 39284 12992 39296
rect 12943 39256 12992 39284
rect 12943 39253 12955 39256
rect 12897 39247 12955 39253
rect 12986 39244 12992 39256
rect 13044 39244 13050 39296
rect 14642 39244 14648 39296
rect 14700 39244 14706 39296
rect 15657 39287 15715 39293
rect 15657 39253 15669 39287
rect 15703 39284 15715 39287
rect 15838 39284 15844 39296
rect 15703 39256 15844 39284
rect 15703 39253 15715 39256
rect 15657 39247 15715 39253
rect 15838 39244 15844 39256
rect 15896 39244 15902 39296
rect 15930 39244 15936 39296
rect 15988 39284 15994 39296
rect 16500 39284 16528 39324
rect 18046 39312 18052 39324
rect 18104 39312 18110 39364
rect 15988 39256 16528 39284
rect 16577 39287 16635 39293
rect 15988 39244 15994 39256
rect 16577 39253 16589 39287
rect 16623 39284 16635 39287
rect 16666 39284 16672 39296
rect 16623 39256 16672 39284
rect 16623 39253 16635 39256
rect 16577 39247 16635 39253
rect 16666 39244 16672 39256
rect 16724 39244 16730 39296
rect 17497 39287 17555 39293
rect 17497 39253 17509 39287
rect 17543 39284 17555 39287
rect 17954 39284 17960 39296
rect 17543 39256 17960 39284
rect 17543 39253 17555 39256
rect 17497 39247 17555 39253
rect 17954 39244 17960 39256
rect 18012 39244 18018 39296
rect 1104 39194 40572 39216
rect 1104 39142 4874 39194
rect 4926 39142 4938 39194
rect 4990 39142 5002 39194
rect 5054 39142 5066 39194
rect 5118 39142 5130 39194
rect 5182 39142 35594 39194
rect 35646 39142 35658 39194
rect 35710 39142 35722 39194
rect 35774 39142 35786 39194
rect 35838 39142 35850 39194
rect 35902 39142 40572 39194
rect 1104 39120 40572 39142
rect 10870 39080 10876 39092
rect 10704 39052 10876 39080
rect 10704 39012 10732 39052
rect 10870 39040 10876 39052
rect 10928 39040 10934 39092
rect 11974 39040 11980 39092
rect 12032 39040 12038 39092
rect 12066 39040 12072 39092
rect 12124 39040 12130 39092
rect 14642 39040 14648 39092
rect 14700 39080 14706 39092
rect 15010 39080 15016 39092
rect 14700 39052 15016 39080
rect 14700 39040 14706 39052
rect 15010 39040 15016 39052
rect 15068 39080 15074 39092
rect 16853 39083 16911 39089
rect 16853 39080 16865 39083
rect 15068 39052 16865 39080
rect 15068 39040 15074 39052
rect 16853 39049 16865 39052
rect 16899 39049 16911 39083
rect 16853 39043 16911 39049
rect 20714 39040 20720 39092
rect 20772 39080 20778 39092
rect 25777 39083 25835 39089
rect 25777 39080 25789 39083
rect 20772 39052 25789 39080
rect 20772 39040 20778 39052
rect 25777 39049 25789 39052
rect 25823 39049 25835 39083
rect 25777 39043 25835 39049
rect 11606 39012 11612 39024
rect 9798 38984 10732 39012
rect 10796 38984 11612 39012
rect 10226 38904 10232 38956
rect 10284 38904 10290 38956
rect 10796 38953 10824 38984
rect 11606 38972 11612 38984
rect 11664 39012 11670 39024
rect 11664 38984 11836 39012
rect 11664 38972 11670 38984
rect 10413 38947 10471 38953
rect 10413 38913 10425 38947
rect 10459 38913 10471 38947
rect 10413 38907 10471 38913
rect 10781 38947 10839 38953
rect 10781 38913 10793 38947
rect 10827 38913 10839 38947
rect 10781 38907 10839 38913
rect 6822 38836 6828 38888
rect 6880 38876 6886 38888
rect 8297 38879 8355 38885
rect 8297 38876 8309 38879
rect 6880 38848 8309 38876
rect 6880 38836 6886 38848
rect 8297 38845 8309 38848
rect 8343 38845 8355 38879
rect 8297 38839 8355 38845
rect 8312 38740 8340 38839
rect 8570 38836 8576 38888
rect 8628 38836 8634 38888
rect 9306 38836 9312 38888
rect 9364 38876 9370 38888
rect 10428 38876 10456 38907
rect 11054 38904 11060 38956
rect 11112 38904 11118 38956
rect 11808 38953 11836 38984
rect 16666 38972 16672 39024
rect 16724 38972 16730 39024
rect 18046 38972 18052 39024
rect 18104 39012 18110 39024
rect 18322 39012 18328 39024
rect 18104 38984 18328 39012
rect 18104 38972 18110 38984
rect 18322 38972 18328 38984
rect 18380 38972 18386 39024
rect 20806 39012 20812 39024
rect 19366 38984 20812 39012
rect 20806 38972 20812 38984
rect 20864 38972 20870 39024
rect 22925 39015 22983 39021
rect 22925 38981 22937 39015
rect 22971 39012 22983 39015
rect 23198 39012 23204 39024
rect 22971 38984 23204 39012
rect 22971 38981 22983 38984
rect 22925 38975 22983 38981
rect 23198 38972 23204 38984
rect 23256 38972 23262 39024
rect 24486 38972 24492 39024
rect 24544 39012 24550 39024
rect 24673 39015 24731 39021
rect 24673 39012 24685 39015
rect 24544 38984 24685 39012
rect 24544 38972 24550 38984
rect 24673 38981 24685 38984
rect 24719 38981 24731 39015
rect 24673 38975 24731 38981
rect 25685 39015 25743 39021
rect 25685 38981 25697 39015
rect 25731 39012 25743 39015
rect 27062 39012 27068 39024
rect 25731 38984 27068 39012
rect 25731 38981 25743 38984
rect 25685 38975 25743 38981
rect 27062 38972 27068 38984
rect 27120 38972 27126 39024
rect 11793 38947 11851 38953
rect 11793 38913 11805 38947
rect 11839 38913 11851 38947
rect 11793 38907 11851 38913
rect 12250 38904 12256 38956
rect 12308 38904 12314 38956
rect 16942 38904 16948 38956
rect 17000 38904 17006 38956
rect 25222 38944 25228 38956
rect 24058 38916 25228 38944
rect 25222 38904 25228 38916
rect 25280 38904 25286 38956
rect 10502 38876 10508 38888
rect 9364 38848 10364 38876
rect 10428 38848 10508 38876
rect 9364 38836 9370 38848
rect 9582 38768 9588 38820
rect 9640 38808 9646 38820
rect 10229 38811 10287 38817
rect 10229 38808 10241 38811
rect 9640 38780 10241 38808
rect 9640 38768 9646 38780
rect 10229 38777 10241 38780
rect 10275 38777 10287 38811
rect 10336 38808 10364 38848
rect 10502 38836 10508 38848
rect 10560 38876 10566 38888
rect 10873 38879 10931 38885
rect 10873 38876 10885 38879
rect 10560 38848 10885 38876
rect 10560 38836 10566 38848
rect 10873 38845 10885 38848
rect 10919 38876 10931 38879
rect 11517 38879 11575 38885
rect 11517 38876 11529 38879
rect 10919 38848 11529 38876
rect 10919 38845 10931 38848
rect 10873 38839 10931 38845
rect 11517 38845 11529 38848
rect 11563 38845 11575 38879
rect 11517 38839 11575 38845
rect 12434 38836 12440 38888
rect 12492 38836 12498 38888
rect 19794 38836 19800 38888
rect 19852 38836 19858 38888
rect 20070 38836 20076 38888
rect 20128 38836 20134 38888
rect 22649 38879 22707 38885
rect 22649 38845 22661 38879
rect 22695 38876 22707 38879
rect 23014 38876 23020 38888
rect 22695 38848 23020 38876
rect 22695 38845 22707 38848
rect 22649 38839 22707 38845
rect 23014 38836 23020 38848
rect 23072 38836 23078 38888
rect 25498 38836 25504 38888
rect 25556 38836 25562 38888
rect 10965 38811 11023 38817
rect 10965 38808 10977 38811
rect 10336 38780 10977 38808
rect 10229 38771 10287 38777
rect 10965 38777 10977 38780
rect 11011 38808 11023 38811
rect 11609 38811 11667 38817
rect 11609 38808 11621 38811
rect 11011 38780 11621 38808
rect 11011 38777 11023 38780
rect 10965 38771 11023 38777
rect 11609 38777 11621 38780
rect 11655 38777 11667 38811
rect 11609 38771 11667 38777
rect 9950 38740 9956 38752
rect 8312 38712 9956 38740
rect 9950 38700 9956 38712
rect 10008 38700 10014 38752
rect 10045 38743 10103 38749
rect 10045 38709 10057 38743
rect 10091 38740 10103 38743
rect 10134 38740 10140 38752
rect 10091 38712 10140 38740
rect 10091 38709 10103 38712
rect 10045 38703 10103 38709
rect 10134 38700 10140 38712
rect 10192 38700 10198 38752
rect 10594 38700 10600 38752
rect 10652 38700 10658 38752
rect 16669 38743 16727 38749
rect 16669 38709 16681 38743
rect 16715 38740 16727 38743
rect 19058 38740 19064 38752
rect 16715 38712 19064 38740
rect 16715 38709 16727 38712
rect 16669 38703 16727 38709
rect 19058 38700 19064 38712
rect 19116 38700 19122 38752
rect 26145 38743 26203 38749
rect 26145 38709 26157 38743
rect 26191 38740 26203 38743
rect 27430 38740 27436 38752
rect 26191 38712 27436 38740
rect 26191 38709 26203 38712
rect 26145 38703 26203 38709
rect 27430 38700 27436 38712
rect 27488 38700 27494 38752
rect 1104 38650 40572 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 40572 38650
rect 1104 38576 40572 38598
rect 8021 38539 8079 38545
rect 8021 38505 8033 38539
rect 8067 38536 8079 38539
rect 8386 38536 8392 38548
rect 8067 38508 8392 38536
rect 8067 38505 8079 38508
rect 8021 38499 8079 38505
rect 8386 38496 8392 38508
rect 8444 38496 8450 38548
rect 8570 38496 8576 38548
rect 8628 38536 8634 38548
rect 8757 38539 8815 38545
rect 8757 38536 8769 38539
rect 8628 38508 8769 38536
rect 8628 38496 8634 38508
rect 8757 38505 8769 38508
rect 8803 38505 8815 38539
rect 8757 38499 8815 38505
rect 9398 38496 9404 38548
rect 9456 38496 9462 38548
rect 9953 38539 10011 38545
rect 9953 38505 9965 38539
rect 9999 38536 10011 38539
rect 10226 38536 10232 38548
rect 9999 38508 10232 38536
rect 9999 38505 10011 38508
rect 9953 38499 10011 38505
rect 10226 38496 10232 38508
rect 10284 38496 10290 38548
rect 10502 38496 10508 38548
rect 10560 38496 10566 38548
rect 11514 38496 11520 38548
rect 11572 38496 11578 38548
rect 13446 38496 13452 38548
rect 13504 38536 13510 38548
rect 15194 38536 15200 38548
rect 13504 38508 15200 38536
rect 13504 38496 13510 38508
rect 15194 38496 15200 38508
rect 15252 38496 15258 38548
rect 18509 38539 18567 38545
rect 18509 38505 18521 38539
rect 18555 38536 18567 38539
rect 19794 38536 19800 38548
rect 18555 38508 19800 38536
rect 18555 38505 18567 38508
rect 18509 38499 18567 38505
rect 19794 38496 19800 38508
rect 19852 38496 19858 38548
rect 19886 38496 19892 38548
rect 19944 38536 19950 38548
rect 19944 38508 22968 38536
rect 19944 38496 19950 38508
rect 7929 38471 7987 38477
rect 7929 38437 7941 38471
rect 7975 38468 7987 38471
rect 7975 38440 8708 38468
rect 7975 38437 7987 38440
rect 7929 38431 7987 38437
rect 7745 38403 7803 38409
rect 7745 38369 7757 38403
rect 7791 38400 7803 38403
rect 8570 38400 8576 38412
rect 7791 38372 8576 38400
rect 7791 38369 7803 38372
rect 7745 38363 7803 38369
rect 8570 38360 8576 38372
rect 8628 38360 8634 38412
rect 8680 38344 8708 38440
rect 8846 38428 8852 38480
rect 8904 38468 8910 38480
rect 8904 38440 9260 38468
rect 8904 38428 8910 38440
rect 5442 38292 5448 38344
rect 5500 38292 5506 38344
rect 5718 38292 5724 38344
rect 5776 38292 5782 38344
rect 8018 38292 8024 38344
rect 8076 38292 8082 38344
rect 8110 38292 8116 38344
rect 8168 38292 8174 38344
rect 8294 38292 8300 38344
rect 8352 38292 8358 38344
rect 8386 38292 8392 38344
rect 8444 38292 8450 38344
rect 8481 38335 8539 38341
rect 8481 38301 8493 38335
rect 8527 38332 8539 38335
rect 8527 38304 8616 38332
rect 8527 38301 8539 38304
rect 8481 38295 8539 38301
rect 5629 38267 5687 38273
rect 5629 38233 5641 38267
rect 5675 38264 5687 38267
rect 7006 38264 7012 38276
rect 5675 38236 7012 38264
rect 5675 38233 5687 38236
rect 5629 38227 5687 38233
rect 7006 38224 7012 38236
rect 7064 38224 7070 38276
rect 8588 38264 8616 38304
rect 8662 38292 8668 38344
rect 8720 38332 8726 38344
rect 8941 38335 8999 38341
rect 8941 38332 8953 38335
rect 8720 38304 8953 38332
rect 8720 38292 8726 38304
rect 8941 38301 8953 38304
rect 8987 38301 8999 38335
rect 8941 38295 8999 38301
rect 9030 38292 9036 38344
rect 9088 38292 9094 38344
rect 9232 38341 9260 38440
rect 12820 38440 16528 38468
rect 9306 38360 9312 38412
rect 9364 38400 9370 38412
rect 9364 38372 11560 38400
rect 9364 38360 9370 38372
rect 9217 38335 9275 38341
rect 9217 38301 9229 38335
rect 9263 38332 9275 38335
rect 9582 38332 9588 38344
rect 9263 38304 9588 38332
rect 9263 38301 9275 38304
rect 9217 38295 9275 38301
rect 9582 38292 9588 38304
rect 9640 38292 9646 38344
rect 9968 38341 9996 38372
rect 9769 38335 9827 38341
rect 9769 38301 9781 38335
rect 9815 38301 9827 38335
rect 9769 38295 9827 38301
rect 9953 38335 10011 38341
rect 9953 38301 9965 38335
rect 9999 38301 10011 38335
rect 9953 38295 10011 38301
rect 9784 38264 9812 38295
rect 10226 38292 10232 38344
rect 10284 38292 10290 38344
rect 10336 38341 10364 38372
rect 10321 38335 10379 38341
rect 10321 38301 10333 38335
rect 10367 38301 10379 38335
rect 10321 38295 10379 38301
rect 11330 38292 11336 38344
rect 11388 38292 11394 38344
rect 11532 38341 11560 38372
rect 11517 38335 11575 38341
rect 11517 38301 11529 38335
rect 11563 38332 11575 38335
rect 12250 38332 12256 38344
rect 11563 38304 12256 38332
rect 11563 38301 11575 38304
rect 11517 38295 11575 38301
rect 12250 38292 12256 38304
rect 12308 38292 12314 38344
rect 12618 38292 12624 38344
rect 12676 38292 12682 38344
rect 12820 38341 12848 38440
rect 12986 38360 12992 38412
rect 13044 38360 13050 38412
rect 13446 38400 13452 38412
rect 13096 38372 13452 38400
rect 12805 38335 12863 38341
rect 12805 38301 12817 38335
rect 12851 38301 12863 38335
rect 12805 38295 12863 38301
rect 12897 38335 12955 38341
rect 12897 38301 12909 38335
rect 12943 38332 12955 38335
rect 13096 38332 13124 38372
rect 13446 38360 13452 38372
rect 13504 38360 13510 38412
rect 12943 38304 13124 38332
rect 12943 38301 12955 38304
rect 12897 38295 12955 38301
rect 13170 38292 13176 38344
rect 13228 38292 13234 38344
rect 10244 38264 10272 38292
rect 8588 38236 9674 38264
rect 4430 38156 4436 38208
rect 4488 38196 4494 38208
rect 5261 38199 5319 38205
rect 5261 38196 5273 38199
rect 4488 38168 5273 38196
rect 4488 38156 4494 38168
rect 5261 38165 5273 38168
rect 5307 38165 5319 38199
rect 9646 38196 9674 38236
rect 9784 38236 10272 38264
rect 11348 38264 11376 38292
rect 12434 38264 12440 38276
rect 11348 38236 12440 38264
rect 9784 38196 9812 38236
rect 12434 38224 12440 38236
rect 12492 38224 12498 38276
rect 16500 38264 16528 38440
rect 20622 38428 20628 38480
rect 20680 38468 20686 38480
rect 20806 38468 20812 38480
rect 20680 38440 20812 38468
rect 20680 38428 20686 38440
rect 20806 38428 20812 38440
rect 20864 38428 20870 38480
rect 21266 38468 21272 38480
rect 20916 38440 21272 38468
rect 16574 38360 16580 38412
rect 16632 38400 16638 38412
rect 20916 38400 20944 38440
rect 21266 38428 21272 38440
rect 21324 38428 21330 38480
rect 16632 38372 20944 38400
rect 16632 38360 16638 38372
rect 17770 38292 17776 38344
rect 17828 38292 17834 38344
rect 17954 38292 17960 38344
rect 18012 38292 18018 38344
rect 18046 38292 18052 38344
rect 18104 38292 18110 38344
rect 18141 38335 18199 38341
rect 18141 38301 18153 38335
rect 18187 38301 18199 38335
rect 18141 38295 18199 38301
rect 18156 38264 18184 38295
rect 18322 38292 18328 38344
rect 18380 38292 18386 38344
rect 19242 38292 19248 38344
rect 19300 38332 19306 38344
rect 20916 38341 20944 38372
rect 20717 38335 20775 38341
rect 20717 38332 20729 38335
rect 19300 38304 20729 38332
rect 19300 38292 19306 38304
rect 20717 38301 20729 38304
rect 20763 38301 20775 38335
rect 20717 38295 20775 38301
rect 20901 38335 20959 38341
rect 20901 38301 20913 38335
rect 20947 38301 20959 38335
rect 20901 38295 20959 38301
rect 18506 38264 18512 38276
rect 16500 38236 18512 38264
rect 18506 38224 18512 38236
rect 18564 38224 18570 38276
rect 9646 38168 9812 38196
rect 5261 38159 5319 38165
rect 11238 38156 11244 38208
rect 11296 38196 11302 38208
rect 12802 38196 12808 38208
rect 11296 38168 12808 38196
rect 11296 38156 11302 38168
rect 12802 38156 12808 38168
rect 12860 38156 12866 38208
rect 13262 38156 13268 38208
rect 13320 38196 13326 38208
rect 13357 38199 13415 38205
rect 13357 38196 13369 38199
rect 13320 38168 13369 38196
rect 13320 38156 13326 38168
rect 13357 38165 13369 38168
rect 13403 38165 13415 38199
rect 13357 38159 13415 38165
rect 14826 38156 14832 38208
rect 14884 38196 14890 38208
rect 18322 38196 18328 38208
rect 14884 38168 18328 38196
rect 14884 38156 14890 38168
rect 18322 38156 18328 38168
rect 18380 38196 18386 38208
rect 19334 38196 19340 38208
rect 18380 38168 19340 38196
rect 18380 38156 18386 38168
rect 19334 38156 19340 38168
rect 19392 38156 19398 38208
rect 20732 38196 20760 38295
rect 21174 38292 21180 38344
rect 21232 38332 21238 38344
rect 21453 38335 21511 38341
rect 21453 38332 21465 38335
rect 21232 38304 21465 38332
rect 21232 38292 21238 38304
rect 21453 38301 21465 38304
rect 21499 38301 21511 38335
rect 21453 38295 21511 38301
rect 21545 38335 21603 38341
rect 21545 38301 21557 38335
rect 21591 38301 21603 38335
rect 21545 38295 21603 38301
rect 21729 38335 21787 38341
rect 21729 38301 21741 38335
rect 21775 38332 21787 38335
rect 22094 38332 22100 38344
rect 21775 38304 22100 38332
rect 21775 38301 21787 38304
rect 21729 38295 21787 38301
rect 21085 38267 21143 38273
rect 21085 38233 21097 38267
rect 21131 38264 21143 38267
rect 21560 38264 21588 38295
rect 22094 38292 22100 38304
rect 22152 38292 22158 38344
rect 22940 38341 22968 38508
rect 23198 38496 23204 38548
rect 23256 38496 23262 38548
rect 23845 38403 23903 38409
rect 23845 38369 23857 38403
rect 23891 38400 23903 38403
rect 25498 38400 25504 38412
rect 23891 38372 25504 38400
rect 23891 38369 23903 38372
rect 23845 38363 23903 38369
rect 25498 38360 25504 38372
rect 25556 38360 25562 38412
rect 26418 38360 26424 38412
rect 26476 38400 26482 38412
rect 26605 38403 26663 38409
rect 26605 38400 26617 38403
rect 26476 38372 26617 38400
rect 26476 38360 26482 38372
rect 26605 38369 26617 38372
rect 26651 38369 26663 38403
rect 26605 38363 26663 38369
rect 26697 38403 26755 38409
rect 26697 38369 26709 38403
rect 26743 38400 26755 38403
rect 27062 38400 27068 38412
rect 26743 38372 27068 38400
rect 26743 38369 26755 38372
rect 26697 38363 26755 38369
rect 27062 38360 27068 38372
rect 27120 38360 27126 38412
rect 27430 38360 27436 38412
rect 27488 38400 27494 38412
rect 28445 38403 28503 38409
rect 28445 38400 28457 38403
rect 27488 38372 28457 38400
rect 27488 38360 27494 38372
rect 28445 38369 28457 38372
rect 28491 38369 28503 38403
rect 28445 38363 28503 38369
rect 22925 38335 22983 38341
rect 22925 38301 22937 38335
rect 22971 38301 22983 38335
rect 22925 38295 22983 38301
rect 23014 38292 23020 38344
rect 23072 38332 23078 38344
rect 24581 38335 24639 38341
rect 24581 38332 24593 38335
rect 23072 38304 24593 38332
rect 23072 38292 23078 38304
rect 24581 38301 24593 38304
rect 24627 38301 24639 38335
rect 24581 38295 24639 38301
rect 28721 38335 28779 38341
rect 28721 38301 28733 38335
rect 28767 38332 28779 38335
rect 28902 38332 28908 38344
rect 28767 38304 28908 38332
rect 28767 38301 28779 38304
rect 28721 38295 28779 38301
rect 28902 38292 28908 38304
rect 28960 38292 28966 38344
rect 23569 38267 23627 38273
rect 23569 38264 23581 38267
rect 21131 38236 21588 38264
rect 23032 38236 23581 38264
rect 21131 38233 21143 38236
rect 21085 38227 21143 38233
rect 21450 38196 21456 38208
rect 20732 38168 21456 38196
rect 21450 38156 21456 38168
rect 21508 38156 21514 38208
rect 21634 38156 21640 38208
rect 21692 38156 21698 38208
rect 23032 38205 23060 38236
rect 23569 38233 23581 38236
rect 23615 38233 23627 38267
rect 23569 38227 23627 38233
rect 23661 38267 23719 38273
rect 23661 38233 23673 38267
rect 23707 38264 23719 38267
rect 24486 38264 24492 38276
rect 23707 38236 24492 38264
rect 23707 38233 23719 38236
rect 23661 38227 23719 38233
rect 24486 38224 24492 38236
rect 24544 38224 24550 38276
rect 24857 38267 24915 38273
rect 24857 38233 24869 38267
rect 24903 38264 24915 38267
rect 24946 38264 24952 38276
rect 24903 38236 24952 38264
rect 24903 38233 24915 38236
rect 24857 38227 24915 38233
rect 24946 38224 24952 38236
rect 25004 38224 25010 38276
rect 25314 38264 25320 38276
rect 25240 38236 25320 38264
rect 23017 38199 23075 38205
rect 23017 38165 23029 38199
rect 23063 38165 23075 38199
rect 25240 38196 25268 38236
rect 25314 38224 25320 38236
rect 25372 38224 25378 38276
rect 26344 38236 27278 38264
rect 26344 38196 26372 38236
rect 25240 38168 26372 38196
rect 23017 38159 23075 38165
rect 1104 38106 40572 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 35594 38106
rect 35646 38054 35658 38106
rect 35710 38054 35722 38106
rect 35774 38054 35786 38106
rect 35838 38054 35850 38106
rect 35902 38054 40572 38106
rect 1104 38032 40572 38054
rect 7006 37992 7012 38004
rect 6196 37964 7012 37992
rect 4430 37884 4436 37936
rect 4488 37884 4494 37936
rect 6196 37933 6224 37964
rect 7006 37952 7012 37964
rect 7064 37952 7070 38004
rect 8662 37952 8668 38004
rect 8720 37952 8726 38004
rect 12802 37952 12808 38004
rect 12860 37992 12866 38004
rect 13170 37992 13176 38004
rect 12860 37964 13176 37992
rect 12860 37952 12866 37964
rect 13170 37952 13176 37964
rect 13228 37992 13234 38004
rect 13228 37964 15976 37992
rect 13228 37952 13234 37964
rect 6181 37927 6239 37933
rect 6181 37893 6193 37927
rect 6227 37893 6239 37927
rect 8680 37924 8708 37952
rect 6181 37887 6239 37893
rect 6288 37896 7130 37924
rect 8680 37896 9628 37924
rect 5902 37856 5908 37868
rect 5566 37828 5908 37856
rect 5902 37816 5908 37828
rect 5960 37856 5966 37868
rect 6288 37856 6316 37896
rect 5960 37828 6316 37856
rect 8849 37859 8907 37865
rect 5960 37816 5966 37828
rect 8849 37825 8861 37859
rect 8895 37856 8907 37859
rect 8938 37856 8944 37868
rect 8895 37828 8944 37856
rect 8895 37825 8907 37828
rect 8849 37819 8907 37825
rect 8938 37816 8944 37828
rect 8996 37816 9002 37868
rect 9125 37859 9183 37865
rect 9125 37856 9137 37859
rect 9048 37828 9137 37856
rect 4157 37791 4215 37797
rect 4157 37757 4169 37791
rect 4203 37757 4215 37791
rect 4157 37751 4215 37757
rect 6365 37791 6423 37797
rect 6365 37757 6377 37791
rect 6411 37757 6423 37791
rect 6365 37751 6423 37757
rect 4172 37652 4200 37751
rect 5534 37652 5540 37664
rect 4172 37624 5540 37652
rect 5534 37612 5540 37624
rect 5592 37652 5598 37664
rect 6380 37652 6408 37751
rect 6638 37748 6644 37800
rect 6696 37748 6702 37800
rect 9048 37797 9076 37828
rect 9125 37825 9137 37828
rect 9171 37825 9183 37859
rect 9125 37819 9183 37825
rect 9306 37816 9312 37868
rect 9364 37816 9370 37868
rect 9600 37865 9628 37896
rect 13262 37884 13268 37936
rect 13320 37884 13326 37936
rect 15010 37924 15016 37936
rect 14490 37896 15016 37924
rect 15010 37884 15016 37896
rect 15068 37884 15074 37936
rect 15473 37927 15531 37933
rect 15473 37893 15485 37927
rect 15519 37924 15531 37927
rect 15948 37924 15976 37964
rect 17770 37952 17776 38004
rect 17828 37992 17834 38004
rect 18049 37995 18107 38001
rect 18049 37992 18061 37995
rect 17828 37964 18061 37992
rect 17828 37952 17834 37964
rect 18049 37961 18061 37964
rect 18095 37961 18107 37995
rect 20070 37992 20076 38004
rect 18049 37955 18107 37961
rect 19812 37964 20076 37992
rect 15519 37896 15792 37924
rect 15519 37893 15531 37896
rect 15473 37887 15531 37893
rect 9401 37859 9459 37865
rect 9401 37825 9413 37859
rect 9447 37825 9459 37859
rect 9401 37819 9459 37825
rect 9585 37859 9643 37865
rect 9585 37825 9597 37859
rect 9631 37825 9643 37859
rect 9585 37819 9643 37825
rect 9033 37791 9091 37797
rect 9033 37757 9045 37791
rect 9079 37757 9091 37791
rect 9033 37751 9091 37757
rect 9217 37791 9275 37797
rect 9217 37757 9229 37791
rect 9263 37788 9275 37791
rect 9416 37788 9444 37819
rect 14826 37816 14832 37868
rect 14884 37856 14890 37868
rect 15105 37859 15163 37865
rect 15105 37856 15117 37859
rect 14884 37828 15117 37856
rect 14884 37816 14890 37828
rect 15105 37825 15117 37828
rect 15151 37825 15163 37859
rect 15105 37819 15163 37825
rect 15289 37859 15347 37865
rect 15289 37825 15301 37859
rect 15335 37825 15347 37859
rect 15289 37819 15347 37825
rect 9263 37760 9444 37788
rect 12989 37791 13047 37797
rect 9263 37757 9275 37760
rect 9217 37751 9275 37757
rect 12989 37757 13001 37791
rect 13035 37757 13047 37791
rect 12989 37751 13047 37757
rect 15013 37791 15071 37797
rect 15013 37757 15025 37791
rect 15059 37788 15071 37791
rect 15194 37788 15200 37800
rect 15059 37760 15200 37788
rect 15059 37757 15071 37760
rect 15013 37751 15071 37757
rect 6822 37652 6828 37664
rect 5592 37624 6828 37652
rect 5592 37612 5598 37624
rect 6822 37612 6828 37624
rect 6880 37612 6886 37664
rect 7926 37612 7932 37664
rect 7984 37652 7990 37664
rect 8113 37655 8171 37661
rect 8113 37652 8125 37655
rect 7984 37624 8125 37652
rect 7984 37612 7990 37624
rect 8113 37621 8125 37624
rect 8159 37652 8171 37655
rect 9048 37652 9076 37751
rect 8159 37624 9076 37652
rect 8159 37621 8171 37624
rect 8113 37615 8171 37621
rect 9122 37612 9128 37664
rect 9180 37652 9186 37664
rect 9401 37655 9459 37661
rect 9401 37652 9413 37655
rect 9180 37624 9413 37652
rect 9180 37612 9186 37624
rect 9401 37621 9413 37624
rect 9447 37621 9459 37655
rect 13004 37652 13032 37751
rect 15194 37748 15200 37760
rect 15252 37748 15258 37800
rect 15304 37788 15332 37819
rect 15378 37816 15384 37868
rect 15436 37856 15442 37868
rect 15764 37865 15792 37896
rect 15948 37896 18092 37924
rect 15565 37859 15623 37865
rect 15565 37856 15577 37859
rect 15436 37828 15577 37856
rect 15436 37816 15442 37828
rect 15565 37825 15577 37828
rect 15611 37825 15623 37859
rect 15565 37819 15623 37825
rect 15749 37859 15807 37865
rect 15749 37825 15761 37859
rect 15795 37825 15807 37859
rect 15749 37819 15807 37825
rect 15838 37816 15844 37868
rect 15896 37816 15902 37868
rect 15948 37865 15976 37896
rect 15933 37859 15991 37865
rect 15933 37825 15945 37859
rect 15979 37825 15991 37859
rect 15933 37819 15991 37825
rect 17402 37816 17408 37868
rect 17460 37856 17466 37868
rect 17589 37859 17647 37865
rect 17589 37856 17601 37859
rect 17460 37828 17601 37856
rect 17460 37816 17466 37828
rect 17589 37825 17601 37828
rect 17635 37825 17647 37859
rect 17589 37819 17647 37825
rect 17678 37816 17684 37868
rect 17736 37816 17742 37868
rect 17865 37859 17923 37865
rect 17865 37825 17877 37859
rect 17911 37825 17923 37859
rect 17865 37819 17923 37825
rect 15304 37760 15608 37788
rect 15580 37732 15608 37760
rect 17310 37748 17316 37800
rect 17368 37788 17374 37800
rect 17880 37788 17908 37819
rect 18064 37800 18092 37896
rect 19242 37884 19248 37936
rect 19300 37924 19306 37936
rect 19300 37896 19564 37924
rect 19300 37884 19306 37896
rect 18138 37816 18144 37868
rect 18196 37856 18202 37868
rect 18417 37859 18475 37865
rect 18417 37856 18429 37859
rect 18196 37828 18429 37856
rect 18196 37816 18202 37828
rect 18417 37825 18429 37828
rect 18463 37825 18475 37859
rect 18417 37819 18475 37825
rect 18966 37816 18972 37868
rect 19024 37816 19030 37868
rect 19150 37816 19156 37868
rect 19208 37816 19214 37868
rect 19334 37816 19340 37868
rect 19392 37816 19398 37868
rect 19536 37865 19564 37896
rect 19812 37865 19840 37964
rect 20070 37952 20076 37964
rect 20128 37992 20134 38004
rect 22370 37992 22376 38004
rect 20128 37964 22376 37992
rect 20128 37952 20134 37964
rect 22370 37952 22376 37964
rect 22428 37952 22434 38004
rect 22480 37964 23980 37992
rect 20622 37884 20628 37936
rect 20680 37884 20686 37936
rect 22480 37924 22508 37964
rect 22296 37896 22508 37924
rect 23952 37924 23980 37964
rect 24946 37952 24952 38004
rect 25004 37952 25010 38004
rect 25409 37995 25467 38001
rect 25409 37961 25421 37995
rect 25455 37992 25467 37995
rect 26418 37992 26424 38004
rect 25455 37964 26424 37992
rect 25455 37961 25467 37964
rect 25409 37955 25467 37961
rect 26418 37952 26424 37964
rect 26476 37952 26482 38004
rect 25317 37927 25375 37933
rect 25317 37924 25329 37927
rect 23952 37896 25329 37924
rect 19521 37859 19579 37865
rect 19521 37825 19533 37859
rect 19567 37825 19579 37859
rect 19521 37819 19579 37825
rect 19797 37859 19855 37865
rect 19797 37825 19809 37859
rect 19843 37825 19855 37859
rect 19797 37819 19855 37825
rect 17368 37760 17908 37788
rect 17368 37748 17374 37760
rect 18046 37748 18052 37800
rect 18104 37788 18110 37800
rect 19242 37788 19248 37800
rect 18104 37760 19248 37788
rect 18104 37748 18110 37760
rect 19242 37748 19248 37760
rect 19300 37748 19306 37800
rect 15562 37680 15568 37732
rect 15620 37680 15626 37732
rect 16758 37680 16764 37732
rect 16816 37720 16822 37732
rect 19536 37720 19564 37819
rect 21542 37816 21548 37868
rect 21600 37856 21606 37868
rect 22005 37859 22063 37865
rect 22005 37856 22017 37859
rect 21600 37828 22017 37856
rect 21600 37816 21606 37828
rect 22005 37825 22017 37828
rect 22051 37825 22063 37859
rect 22005 37819 22063 37825
rect 22094 37816 22100 37868
rect 22152 37816 22158 37868
rect 19705 37791 19763 37797
rect 19705 37757 19717 37791
rect 19751 37788 19763 37791
rect 20073 37791 20131 37797
rect 20073 37788 20085 37791
rect 19751 37760 20085 37788
rect 19751 37757 19763 37760
rect 19705 37751 19763 37757
rect 20073 37757 20085 37760
rect 20119 37757 20131 37791
rect 20073 37751 20131 37757
rect 21818 37748 21824 37800
rect 21876 37748 21882 37800
rect 22296 37720 22324 37896
rect 25317 37893 25329 37896
rect 25363 37893 25375 37927
rect 25317 37887 25375 37893
rect 25222 37856 25228 37868
rect 23782 37828 25228 37856
rect 25222 37816 25228 37828
rect 25280 37816 25286 37868
rect 22370 37748 22376 37800
rect 22428 37748 22434 37800
rect 22646 37748 22652 37800
rect 22704 37748 22710 37800
rect 23842 37748 23848 37800
rect 23900 37788 23906 37800
rect 24397 37791 24455 37797
rect 24397 37788 24409 37791
rect 23900 37760 24409 37788
rect 23900 37748 23906 37760
rect 24397 37757 24409 37760
rect 24443 37757 24455 37791
rect 24397 37751 24455 37757
rect 25498 37748 25504 37800
rect 25556 37748 25562 37800
rect 16816 37692 19564 37720
rect 21100 37692 22324 37720
rect 16816 37680 16822 37692
rect 13722 37652 13728 37664
rect 13004 37624 13728 37652
rect 9401 37615 9459 37621
rect 13722 37612 13728 37624
rect 13780 37612 13786 37664
rect 15286 37612 15292 37664
rect 15344 37652 15350 37664
rect 16209 37655 16267 37661
rect 16209 37652 16221 37655
rect 15344 37624 16221 37652
rect 15344 37612 15350 37624
rect 16209 37621 16221 37624
rect 16255 37621 16267 37655
rect 16209 37615 16267 37621
rect 18509 37655 18567 37661
rect 18509 37621 18521 37655
rect 18555 37652 18567 37655
rect 18598 37652 18604 37664
rect 18555 37624 18604 37652
rect 18555 37621 18567 37624
rect 18509 37615 18567 37621
rect 18598 37612 18604 37624
rect 18656 37652 18662 37664
rect 21100 37652 21128 37692
rect 18656 37624 21128 37652
rect 18656 37612 18662 37624
rect 21450 37612 21456 37664
rect 21508 37652 21514 37664
rect 21545 37655 21603 37661
rect 21545 37652 21557 37655
rect 21508 37624 21557 37652
rect 21508 37612 21514 37624
rect 21545 37621 21557 37624
rect 21591 37621 21603 37655
rect 21545 37615 21603 37621
rect 21910 37612 21916 37664
rect 21968 37612 21974 37664
rect 22388 37652 22416 37748
rect 23014 37652 23020 37664
rect 22388 37624 23020 37652
rect 23014 37612 23020 37624
rect 23072 37612 23078 37664
rect 1104 37562 40572 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 40572 37562
rect 1104 37488 40572 37510
rect 6457 37451 6515 37457
rect 6457 37417 6469 37451
rect 6503 37448 6515 37451
rect 6638 37448 6644 37460
rect 6503 37420 6644 37448
rect 6503 37417 6515 37420
rect 6457 37411 6515 37417
rect 6638 37408 6644 37420
rect 6696 37408 6702 37460
rect 7837 37451 7895 37457
rect 7837 37417 7849 37451
rect 7883 37448 7895 37451
rect 8110 37448 8116 37460
rect 7883 37420 8116 37448
rect 7883 37417 7895 37420
rect 7837 37411 7895 37417
rect 8110 37408 8116 37420
rect 8168 37408 8174 37460
rect 8846 37408 8852 37460
rect 8904 37448 8910 37460
rect 8941 37451 8999 37457
rect 8941 37448 8953 37451
rect 8904 37420 8953 37448
rect 8904 37408 8910 37420
rect 8941 37417 8953 37420
rect 8987 37417 8999 37451
rect 8941 37411 8999 37417
rect 12618 37408 12624 37460
rect 12676 37448 12682 37460
rect 12713 37451 12771 37457
rect 12713 37448 12725 37451
rect 12676 37420 12725 37448
rect 12676 37408 12682 37420
rect 12713 37417 12725 37420
rect 12759 37417 12771 37451
rect 12713 37411 12771 37417
rect 14921 37451 14979 37457
rect 14921 37417 14933 37451
rect 14967 37448 14979 37451
rect 15378 37448 15384 37460
rect 14967 37420 15384 37448
rect 14967 37417 14979 37420
rect 14921 37411 14979 37417
rect 15378 37408 15384 37420
rect 15436 37408 15442 37460
rect 17310 37408 17316 37460
rect 17368 37408 17374 37460
rect 17589 37451 17647 37457
rect 17589 37417 17601 37451
rect 17635 37448 17647 37451
rect 17678 37448 17684 37460
rect 17635 37420 17684 37448
rect 17635 37417 17647 37420
rect 17589 37411 17647 37417
rect 17678 37408 17684 37420
rect 17736 37408 17742 37460
rect 19150 37408 19156 37460
rect 19208 37448 19214 37460
rect 20533 37451 20591 37457
rect 20533 37448 20545 37451
rect 19208 37420 20545 37448
rect 19208 37408 19214 37420
rect 20533 37417 20545 37420
rect 20579 37417 20591 37451
rect 20533 37411 20591 37417
rect 21361 37451 21419 37457
rect 21361 37417 21373 37451
rect 21407 37448 21419 37451
rect 21818 37448 21824 37460
rect 21407 37420 21824 37448
rect 21407 37417 21419 37420
rect 21361 37411 21419 37417
rect 21818 37408 21824 37420
rect 21876 37408 21882 37460
rect 22646 37408 22652 37460
rect 22704 37448 22710 37460
rect 23017 37451 23075 37457
rect 23017 37448 23029 37451
rect 22704 37420 23029 37448
rect 22704 37408 22710 37420
rect 23017 37417 23029 37420
rect 23063 37417 23075 37451
rect 23017 37411 23075 37417
rect 7006 37380 7012 37392
rect 6104 37352 7012 37380
rect 6104 37321 6132 37352
rect 7006 37340 7012 37352
rect 7064 37380 7070 37392
rect 8202 37380 8208 37392
rect 7064 37352 8208 37380
rect 7064 37340 7070 37352
rect 8202 37340 8208 37352
rect 8260 37380 8266 37392
rect 14826 37380 14832 37392
rect 8260 37352 14832 37380
rect 8260 37340 8266 37352
rect 14826 37340 14832 37352
rect 14884 37340 14890 37392
rect 17402 37340 17408 37392
rect 17460 37380 17466 37392
rect 18046 37380 18052 37392
rect 17460 37352 18052 37380
rect 17460 37340 17466 37352
rect 18046 37340 18052 37352
rect 18104 37340 18110 37392
rect 21542 37380 21548 37392
rect 20732 37352 21548 37380
rect 5169 37315 5227 37321
rect 5169 37281 5181 37315
rect 5215 37312 5227 37315
rect 6089 37315 6147 37321
rect 5215 37284 5948 37312
rect 5215 37281 5227 37284
rect 5169 37275 5227 37281
rect 5353 37247 5411 37253
rect 5353 37213 5365 37247
rect 5399 37244 5411 37247
rect 5442 37244 5448 37256
rect 5399 37216 5448 37244
rect 5399 37213 5411 37216
rect 5353 37207 5411 37213
rect 5442 37204 5448 37216
rect 5500 37204 5506 37256
rect 5537 37247 5595 37253
rect 5537 37213 5549 37247
rect 5583 37213 5595 37247
rect 5537 37207 5595 37213
rect 5552 37108 5580 37207
rect 5626 37204 5632 37256
rect 5684 37204 5690 37256
rect 5920 37253 5948 37284
rect 6089 37281 6101 37315
rect 6135 37281 6147 37315
rect 8018 37312 8024 37324
rect 6089 37275 6147 37281
rect 7668 37284 8024 37312
rect 5721 37247 5779 37253
rect 5721 37213 5733 37247
rect 5767 37213 5779 37247
rect 5721 37207 5779 37213
rect 5905 37247 5963 37253
rect 5905 37213 5917 37247
rect 5951 37213 5963 37247
rect 5905 37207 5963 37213
rect 5736 37176 5764 37207
rect 5994 37204 6000 37256
rect 6052 37204 6058 37256
rect 6273 37247 6331 37253
rect 6273 37213 6285 37247
rect 6319 37244 6331 37247
rect 7668 37244 7696 37284
rect 8018 37272 8024 37284
rect 8076 37272 8082 37324
rect 8113 37315 8171 37321
rect 8113 37281 8125 37315
rect 8159 37312 8171 37315
rect 8478 37312 8484 37324
rect 8159 37284 8484 37312
rect 8159 37281 8171 37284
rect 8113 37275 8171 37281
rect 8478 37272 8484 37284
rect 8536 37312 8542 37324
rect 8662 37312 8668 37324
rect 8536 37284 8668 37312
rect 8536 37272 8542 37284
rect 8662 37272 8668 37284
rect 8720 37272 8726 37324
rect 12158 37272 12164 37324
rect 12216 37312 12222 37324
rect 12253 37315 12311 37321
rect 12253 37312 12265 37315
rect 12216 37284 12265 37312
rect 12216 37272 12222 37284
rect 12253 37281 12265 37284
rect 12299 37281 12311 37315
rect 12253 37275 12311 37281
rect 6319 37216 7696 37244
rect 7745 37247 7803 37253
rect 6319 37213 6331 37216
rect 6273 37207 6331 37213
rect 7745 37213 7757 37247
rect 7791 37244 7803 37247
rect 7834 37244 7840 37256
rect 7791 37216 7840 37244
rect 7791 37213 7803 37216
rect 7745 37207 7803 37213
rect 7834 37204 7840 37216
rect 7892 37204 7898 37256
rect 7929 37247 7987 37253
rect 7929 37213 7941 37247
rect 7975 37244 7987 37247
rect 7975 37216 8064 37244
rect 7975 37213 7987 37216
rect 7929 37207 7987 37213
rect 8036 37188 8064 37216
rect 8386 37204 8392 37256
rect 8444 37204 8450 37256
rect 8573 37247 8631 37253
rect 8573 37213 8585 37247
rect 8619 37244 8631 37247
rect 8846 37244 8852 37256
rect 8619 37216 8852 37244
rect 8619 37213 8631 37216
rect 8573 37207 8631 37213
rect 8846 37204 8852 37216
rect 8904 37204 8910 37256
rect 9122 37204 9128 37256
rect 9180 37204 9186 37256
rect 9309 37247 9367 37253
rect 9309 37213 9321 37247
rect 9355 37213 9367 37247
rect 9309 37207 9367 37213
rect 5736 37148 7880 37176
rect 5810 37108 5816 37120
rect 5552 37080 5816 37108
rect 5810 37068 5816 37080
rect 5868 37068 5874 37120
rect 7852 37108 7880 37148
rect 8018 37136 8024 37188
rect 8076 37136 8082 37188
rect 8478 37136 8484 37188
rect 8536 37176 8542 37188
rect 9324 37176 9352 37207
rect 9398 37204 9404 37256
rect 9456 37204 9462 37256
rect 8536 37148 9352 37176
rect 12268 37176 12296 37275
rect 12434 37272 12440 37324
rect 12492 37272 12498 37324
rect 15286 37272 15292 37324
rect 15344 37272 15350 37324
rect 15654 37272 15660 37324
rect 15712 37312 15718 37324
rect 15712 37284 16528 37312
rect 15712 37272 15718 37284
rect 12342 37204 12348 37256
rect 12400 37244 12406 37256
rect 12526 37244 12532 37256
rect 12400 37216 12532 37244
rect 12400 37204 12406 37216
rect 12526 37204 12532 37216
rect 12584 37204 12590 37256
rect 12618 37204 12624 37256
rect 12676 37204 12682 37256
rect 12805 37247 12863 37253
rect 12805 37213 12817 37247
rect 12851 37244 12863 37247
rect 14182 37244 14188 37256
rect 12851 37216 14188 37244
rect 12851 37213 12863 37216
rect 12805 37207 12863 37213
rect 14182 37204 14188 37216
rect 14240 37204 14246 37256
rect 14461 37247 14519 37253
rect 14461 37213 14473 37247
rect 14507 37244 14519 37247
rect 14642 37244 14648 37256
rect 14507 37216 14648 37244
rect 14507 37213 14519 37216
rect 14461 37207 14519 37213
rect 14642 37204 14648 37216
rect 14700 37204 14706 37256
rect 14734 37204 14740 37256
rect 14792 37204 14798 37256
rect 15013 37247 15071 37253
rect 15013 37213 15025 37247
rect 15059 37213 15071 37247
rect 16500 37244 16528 37284
rect 17218 37272 17224 37324
rect 17276 37272 17282 37324
rect 18509 37315 18567 37321
rect 18509 37312 18521 37315
rect 18064 37284 18521 37312
rect 17037 37247 17095 37253
rect 17037 37244 17049 37247
rect 16500 37216 17049 37244
rect 15013 37207 15071 37213
rect 17037 37213 17049 37216
rect 17083 37213 17095 37247
rect 17037 37207 17095 37213
rect 17497 37247 17555 37253
rect 17497 37213 17509 37247
rect 17543 37244 17555 37247
rect 17678 37244 17684 37256
rect 17543 37216 17684 37244
rect 17543 37213 17555 37216
rect 17497 37207 17555 37213
rect 12268 37148 12434 37176
rect 8536 37136 8542 37148
rect 8297 37111 8355 37117
rect 8297 37108 8309 37111
rect 7852 37080 8309 37108
rect 8297 37077 8309 37080
rect 8343 37077 8355 37111
rect 8297 37071 8355 37077
rect 12250 37068 12256 37120
rect 12308 37068 12314 37120
rect 12406 37108 12434 37148
rect 13814 37136 13820 37188
rect 13872 37176 13878 37188
rect 15028 37176 15056 37207
rect 17678 37204 17684 37216
rect 17736 37204 17742 37256
rect 17770 37204 17776 37256
rect 17828 37204 17834 37256
rect 17954 37204 17960 37256
rect 18012 37244 18018 37256
rect 18064 37253 18092 37284
rect 18509 37281 18521 37284
rect 18555 37281 18567 37315
rect 18509 37275 18567 37281
rect 18049 37247 18107 37253
rect 18049 37244 18061 37247
rect 18012 37216 18061 37244
rect 18012 37204 18018 37216
rect 18049 37213 18061 37216
rect 18095 37213 18107 37247
rect 18049 37207 18107 37213
rect 18230 37204 18236 37256
rect 18288 37244 18294 37256
rect 18325 37247 18383 37253
rect 18325 37244 18337 37247
rect 18288 37216 18337 37244
rect 18288 37204 18294 37216
rect 18325 37213 18337 37216
rect 18371 37213 18383 37247
rect 18325 37207 18383 37213
rect 18417 37247 18475 37253
rect 18417 37213 18429 37247
rect 18463 37213 18475 37247
rect 18417 37207 18475 37213
rect 17862 37176 17868 37188
rect 13872 37148 15056 37176
rect 16514 37148 17868 37176
rect 13872 37136 13878 37148
rect 17862 37136 17868 37148
rect 17920 37136 17926 37188
rect 18432 37176 18460 37207
rect 17972 37148 18460 37176
rect 18524 37176 18552 37275
rect 18598 37272 18604 37324
rect 18656 37272 18662 37324
rect 19058 37272 19064 37324
rect 19116 37312 19122 37324
rect 20732 37321 20760 37352
rect 21542 37340 21548 37352
rect 21600 37340 21606 37392
rect 21729 37383 21787 37389
rect 21729 37349 21741 37383
rect 21775 37380 21787 37383
rect 22094 37380 22100 37392
rect 21775 37352 22100 37380
rect 21775 37349 21787 37352
rect 21729 37343 21787 37349
rect 22094 37340 22100 37352
rect 22152 37340 22158 37392
rect 23842 37380 23848 37392
rect 23492 37352 23848 37380
rect 20717 37315 20775 37321
rect 20717 37312 20729 37315
rect 19116 37284 20729 37312
rect 19116 37272 19122 37284
rect 20717 37281 20729 37284
rect 20763 37281 20775 37315
rect 21634 37312 21640 37324
rect 20717 37275 20775 37281
rect 20824 37284 21640 37312
rect 19245 37247 19303 37253
rect 19245 37213 19257 37247
rect 19291 37244 19303 37247
rect 19334 37244 19340 37256
rect 19291 37216 19340 37244
rect 19291 37213 19303 37216
rect 19245 37207 19303 37213
rect 19334 37204 19340 37216
rect 19392 37244 19398 37256
rect 19392 37216 19656 37244
rect 19392 37204 19398 37216
rect 19628 37176 19656 37216
rect 19702 37204 19708 37256
rect 19760 37204 19766 37256
rect 20824 37253 20852 37284
rect 21634 37272 21640 37284
rect 21692 37272 21698 37324
rect 23492 37321 23520 37352
rect 23842 37340 23848 37352
rect 23900 37340 23906 37392
rect 23477 37315 23535 37321
rect 23477 37281 23489 37315
rect 23523 37281 23535 37315
rect 23477 37275 23535 37281
rect 23661 37315 23719 37321
rect 23661 37281 23673 37315
rect 23707 37312 23719 37315
rect 25498 37312 25504 37324
rect 23707 37284 25504 37312
rect 23707 37281 23719 37284
rect 23661 37275 23719 37281
rect 25498 37272 25504 37284
rect 25556 37312 25562 37324
rect 25958 37312 25964 37324
rect 25556 37284 25964 37312
rect 25556 37272 25562 37284
rect 25958 37272 25964 37284
rect 26016 37272 26022 37324
rect 20809 37247 20867 37253
rect 20809 37213 20821 37247
rect 20855 37213 20867 37247
rect 20809 37207 20867 37213
rect 21266 37204 21272 37256
rect 21324 37204 21330 37256
rect 21450 37204 21456 37256
rect 21508 37244 21514 37256
rect 21545 37247 21603 37253
rect 21545 37244 21557 37247
rect 21508 37216 21557 37244
rect 21508 37204 21514 37216
rect 21545 37213 21557 37216
rect 21591 37213 21603 37247
rect 21545 37207 21603 37213
rect 21729 37247 21787 37253
rect 21729 37213 21741 37247
rect 21775 37213 21787 37247
rect 21729 37207 21787 37213
rect 25869 37247 25927 37253
rect 25869 37213 25881 37247
rect 25915 37244 25927 37247
rect 27706 37244 27712 37256
rect 25915 37216 27712 37244
rect 25915 37213 25927 37216
rect 25869 37207 25927 37213
rect 19886 37176 19892 37188
rect 18524 37148 19564 37176
rect 19628 37148 19892 37176
rect 13998 37108 14004 37120
rect 12406 37080 14004 37108
rect 13998 37068 14004 37080
rect 14056 37068 14062 37120
rect 14553 37111 14611 37117
rect 14553 37077 14565 37111
rect 14599 37108 14611 37111
rect 15654 37108 15660 37120
rect 14599 37080 15660 37108
rect 14599 37077 14611 37080
rect 14553 37071 14611 37077
rect 15654 37068 15660 37080
rect 15712 37068 15718 37120
rect 16022 37068 16028 37120
rect 16080 37108 16086 37120
rect 17972 37117 18000 37148
rect 17957 37111 18015 37117
rect 17957 37108 17969 37111
rect 16080 37080 17969 37108
rect 16080 37068 16086 37080
rect 17957 37077 17969 37080
rect 18003 37077 18015 37111
rect 17957 37071 18015 37077
rect 18690 37068 18696 37120
rect 18748 37108 18754 37120
rect 18785 37111 18843 37117
rect 18785 37108 18797 37111
rect 18748 37080 18797 37108
rect 18748 37068 18754 37080
rect 18785 37077 18797 37080
rect 18831 37108 18843 37111
rect 19337 37111 19395 37117
rect 19337 37108 19349 37111
rect 18831 37080 19349 37108
rect 18831 37077 18843 37080
rect 18785 37071 18843 37077
rect 19337 37077 19349 37080
rect 19383 37077 19395 37111
rect 19337 37071 19395 37077
rect 19426 37068 19432 37120
rect 19484 37068 19490 37120
rect 19536 37108 19564 37148
rect 19886 37136 19892 37148
rect 19944 37136 19950 37188
rect 21284 37176 21312 37204
rect 21744 37176 21772 37207
rect 27706 37204 27712 37216
rect 27764 37204 27770 37256
rect 21284 37148 21772 37176
rect 22554 37136 22560 37188
rect 22612 37176 22618 37188
rect 25777 37179 25835 37185
rect 25777 37176 25789 37179
rect 22612 37148 25789 37176
rect 22612 37136 22618 37148
rect 25777 37145 25789 37148
rect 25823 37145 25835 37179
rect 25777 37139 25835 37145
rect 23385 37111 23443 37117
rect 23385 37108 23397 37111
rect 19536 37080 23397 37108
rect 23385 37077 23397 37080
rect 23431 37077 23443 37111
rect 23385 37071 23443 37077
rect 25038 37068 25044 37120
rect 25096 37108 25102 37120
rect 25409 37111 25467 37117
rect 25409 37108 25421 37111
rect 25096 37080 25421 37108
rect 25096 37068 25102 37080
rect 25409 37077 25421 37080
rect 25455 37077 25467 37111
rect 25409 37071 25467 37077
rect 1104 37018 40572 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 40572 37018
rect 1104 36944 40572 36966
rect 5994 36864 6000 36916
rect 6052 36864 6058 36916
rect 8386 36864 8392 36916
rect 8444 36904 8450 36916
rect 8481 36907 8539 36913
rect 8481 36904 8493 36907
rect 8444 36876 8493 36904
rect 8444 36864 8450 36876
rect 8481 36873 8493 36876
rect 8527 36873 8539 36907
rect 8481 36867 8539 36873
rect 9766 36864 9772 36916
rect 9824 36904 9830 36916
rect 10870 36904 10876 36916
rect 9824 36876 10876 36904
rect 9824 36864 9830 36876
rect 10870 36864 10876 36876
rect 10928 36864 10934 36916
rect 11698 36864 11704 36916
rect 11756 36904 11762 36916
rect 11793 36907 11851 36913
rect 11793 36904 11805 36907
rect 11756 36876 11805 36904
rect 11756 36864 11762 36876
rect 11793 36873 11805 36876
rect 11839 36904 11851 36907
rect 12342 36904 12348 36916
rect 11839 36876 12348 36904
rect 11839 36873 11851 36876
rect 11793 36867 11851 36873
rect 12342 36864 12348 36876
rect 12400 36864 12406 36916
rect 12529 36907 12587 36913
rect 12529 36873 12541 36907
rect 12575 36904 12587 36907
rect 12618 36904 12624 36916
rect 12575 36876 12624 36904
rect 12575 36873 12587 36876
rect 12529 36867 12587 36873
rect 12618 36864 12624 36876
rect 12676 36864 12682 36916
rect 15194 36904 15200 36916
rect 13924 36876 15200 36904
rect 6457 36839 6515 36845
rect 6457 36836 6469 36839
rect 5828 36808 6469 36836
rect 5828 36780 5856 36808
rect 6457 36805 6469 36808
rect 6503 36805 6515 36839
rect 6457 36799 6515 36805
rect 8757 36839 8815 36845
rect 8757 36805 8769 36839
rect 8803 36836 8815 36839
rect 9122 36836 9128 36848
rect 8803 36808 9128 36836
rect 8803 36805 8815 36808
rect 8757 36799 8815 36805
rect 9122 36796 9128 36808
rect 9180 36796 9186 36848
rect 10594 36796 10600 36848
rect 10652 36836 10658 36848
rect 12710 36836 12716 36848
rect 10652 36808 11008 36836
rect 10652 36796 10658 36808
rect 5442 36728 5448 36780
rect 5500 36768 5506 36780
rect 5537 36771 5595 36777
rect 5537 36768 5549 36771
rect 5500 36740 5549 36768
rect 5500 36728 5506 36740
rect 5537 36737 5549 36740
rect 5583 36737 5595 36771
rect 5537 36731 5595 36737
rect 5810 36728 5816 36780
rect 5868 36728 5874 36780
rect 5997 36771 6055 36777
rect 5997 36737 6009 36771
rect 6043 36737 6055 36771
rect 5997 36731 6055 36737
rect 6012 36700 6040 36731
rect 6362 36728 6368 36780
rect 6420 36728 6426 36780
rect 6549 36771 6607 36777
rect 6549 36737 6561 36771
rect 6595 36768 6607 36771
rect 8294 36768 8300 36780
rect 6595 36740 8300 36768
rect 6595 36737 6607 36740
rect 6549 36731 6607 36737
rect 8294 36728 8300 36740
rect 8352 36728 8358 36780
rect 8478 36728 8484 36780
rect 8536 36728 8542 36780
rect 8573 36771 8631 36777
rect 8573 36737 8585 36771
rect 8619 36768 8631 36771
rect 8846 36768 8852 36780
rect 8619 36740 8852 36768
rect 8619 36737 8631 36740
rect 8573 36731 8631 36737
rect 8846 36728 8852 36740
rect 8904 36768 8910 36780
rect 9398 36768 9404 36780
rect 8904 36740 9404 36768
rect 8904 36728 8910 36740
rect 9398 36728 9404 36740
rect 9456 36728 9462 36780
rect 10686 36728 10692 36780
rect 10744 36728 10750 36780
rect 10980 36777 11008 36808
rect 12406 36808 12716 36836
rect 10781 36771 10839 36777
rect 10781 36737 10793 36771
rect 10827 36737 10839 36771
rect 10781 36731 10839 36737
rect 10965 36771 11023 36777
rect 10965 36737 10977 36771
rect 11011 36737 11023 36771
rect 10965 36731 11023 36737
rect 11057 36771 11115 36777
rect 11057 36737 11069 36771
rect 11103 36768 11115 36771
rect 11146 36768 11152 36780
rect 11103 36740 11152 36768
rect 11103 36737 11115 36740
rect 11057 36731 11115 36737
rect 6086 36700 6092 36712
rect 6012 36672 6092 36700
rect 6086 36660 6092 36672
rect 6144 36700 6150 36712
rect 8018 36700 8024 36712
rect 6144 36672 8024 36700
rect 6144 36660 6150 36672
rect 8018 36660 8024 36672
rect 8076 36660 8082 36712
rect 10796 36700 10824 36731
rect 11146 36728 11152 36740
rect 11204 36728 11210 36780
rect 11701 36771 11759 36777
rect 11701 36737 11713 36771
rect 11747 36768 11759 36771
rect 12161 36771 12219 36777
rect 11747 36740 12112 36768
rect 11747 36737 11759 36740
rect 11701 36731 11759 36737
rect 11330 36700 11336 36712
rect 10796 36672 11336 36700
rect 11330 36660 11336 36672
rect 11388 36700 11394 36712
rect 11974 36700 11980 36712
rect 11388 36672 11980 36700
rect 11388 36660 11394 36672
rect 11974 36660 11980 36672
rect 12032 36660 12038 36712
rect 3970 36592 3976 36644
rect 4028 36632 4034 36644
rect 9214 36632 9220 36644
rect 4028 36604 9220 36632
rect 4028 36592 4034 36604
rect 9214 36592 9220 36604
rect 9272 36592 9278 36644
rect 12084 36632 12112 36740
rect 12161 36737 12173 36771
rect 12207 36768 12219 36771
rect 12406 36768 12434 36808
rect 12710 36796 12716 36808
rect 12768 36836 12774 36848
rect 13170 36836 13176 36848
rect 12768 36808 13176 36836
rect 12768 36796 12774 36808
rect 13170 36796 13176 36808
rect 13228 36836 13234 36848
rect 13924 36836 13952 36876
rect 15194 36864 15200 36876
rect 15252 36864 15258 36916
rect 15654 36864 15660 36916
rect 15712 36864 15718 36916
rect 16114 36864 16120 36916
rect 16172 36904 16178 36916
rect 16172 36876 17080 36904
rect 16172 36864 16178 36876
rect 13228 36808 13952 36836
rect 13228 36796 13234 36808
rect 12207 36740 12434 36768
rect 12897 36771 12955 36777
rect 12207 36737 12219 36740
rect 12161 36731 12219 36737
rect 12897 36737 12909 36771
rect 12943 36768 12955 36771
rect 13078 36768 13084 36780
rect 12943 36740 13084 36768
rect 12943 36737 12955 36740
rect 12897 36731 12955 36737
rect 13078 36728 13084 36740
rect 13136 36728 13142 36780
rect 13538 36728 13544 36780
rect 13596 36728 13602 36780
rect 13817 36771 13875 36777
rect 13817 36737 13829 36771
rect 13863 36768 13875 36771
rect 13924 36768 13952 36808
rect 14274 36796 14280 36848
rect 14332 36836 14338 36848
rect 14461 36839 14519 36845
rect 14461 36836 14473 36839
rect 14332 36808 14473 36836
rect 14332 36796 14338 36808
rect 14461 36805 14473 36808
rect 14507 36805 14519 36839
rect 15381 36839 15439 36845
rect 15381 36836 15393 36839
rect 14461 36799 14519 36805
rect 14568 36808 15393 36836
rect 13863 36740 13952 36768
rect 13863 36737 13875 36740
rect 13817 36731 13875 36737
rect 13998 36728 14004 36780
rect 14056 36768 14062 36780
rect 14568 36768 14596 36808
rect 15381 36805 15393 36808
rect 15427 36805 15439 36839
rect 15381 36799 15439 36805
rect 15565 36839 15623 36845
rect 15565 36805 15577 36839
rect 15611 36836 15623 36839
rect 17052 36836 17080 36876
rect 18230 36864 18236 36916
rect 18288 36864 18294 36916
rect 18966 36864 18972 36916
rect 19024 36864 19030 36916
rect 24946 36864 24952 36916
rect 25004 36904 25010 36916
rect 25314 36904 25320 36916
rect 25004 36876 25320 36904
rect 25004 36864 25010 36876
rect 25314 36864 25320 36876
rect 25372 36904 25378 36916
rect 25372 36876 25537 36904
rect 25372 36864 25378 36876
rect 20714 36836 20720 36848
rect 15611 36808 16344 36836
rect 15611 36805 15623 36808
rect 15565 36799 15623 36805
rect 14056 36740 14596 36768
rect 14056 36728 14062 36740
rect 15194 36728 15200 36780
rect 15252 36728 15258 36780
rect 15286 36728 15292 36780
rect 15344 36768 15350 36780
rect 15841 36771 15899 36777
rect 15841 36768 15853 36771
rect 15344 36740 15853 36768
rect 15344 36728 15350 36740
rect 15841 36737 15853 36740
rect 15887 36768 15899 36771
rect 16022 36768 16028 36780
rect 15887 36740 16028 36768
rect 15887 36737 15899 36740
rect 15841 36731 15899 36737
rect 16022 36728 16028 36740
rect 16080 36728 16086 36780
rect 16114 36728 16120 36780
rect 16172 36728 16178 36780
rect 16316 36777 16344 36808
rect 17052 36808 20720 36836
rect 17052 36777 17080 36808
rect 20714 36796 20720 36808
rect 20772 36796 20778 36848
rect 25038 36796 25044 36848
rect 25096 36796 25102 36848
rect 25509 36808 25537 36876
rect 26789 36839 26847 36845
rect 26789 36805 26801 36839
rect 26835 36836 26847 36839
rect 27706 36836 27712 36848
rect 26835 36808 27712 36836
rect 26835 36805 26847 36808
rect 26789 36799 26847 36805
rect 27706 36796 27712 36808
rect 27764 36796 27770 36848
rect 16301 36771 16359 36777
rect 16301 36737 16313 36771
rect 16347 36768 16359 36771
rect 16853 36771 16911 36777
rect 16853 36768 16865 36771
rect 16347 36740 16865 36768
rect 16347 36737 16359 36740
rect 16301 36731 16359 36737
rect 16853 36737 16865 36740
rect 16899 36737 16911 36771
rect 16853 36731 16911 36737
rect 17037 36771 17095 36777
rect 17037 36737 17049 36771
rect 17083 36737 17095 36771
rect 17037 36731 17095 36737
rect 17126 36728 17132 36780
rect 17184 36768 17190 36780
rect 17954 36768 17960 36780
rect 17184 36740 17960 36768
rect 17184 36728 17190 36740
rect 17954 36728 17960 36740
rect 18012 36728 18018 36780
rect 18046 36728 18052 36780
rect 18104 36728 18110 36780
rect 18690 36728 18696 36780
rect 18748 36728 18754 36780
rect 23750 36728 23756 36780
rect 23808 36728 23814 36780
rect 12250 36660 12256 36712
rect 12308 36660 12314 36712
rect 12989 36703 13047 36709
rect 12989 36669 13001 36703
rect 13035 36700 13047 36703
rect 13357 36703 13415 36709
rect 13357 36700 13369 36703
rect 13035 36672 13369 36700
rect 13035 36669 13047 36672
rect 12989 36663 13047 36669
rect 13357 36669 13369 36672
rect 13403 36669 13415 36703
rect 13357 36663 13415 36669
rect 14182 36660 14188 36712
rect 14240 36660 14246 36712
rect 14369 36703 14427 36709
rect 14369 36669 14381 36703
rect 14415 36669 14427 36703
rect 14369 36663 14427 36669
rect 12894 36632 12900 36644
rect 10428 36604 10732 36632
rect 12084 36604 12900 36632
rect 5626 36524 5632 36576
rect 5684 36573 5690 36576
rect 5684 36567 5733 36573
rect 5684 36533 5687 36567
rect 5721 36533 5733 36567
rect 5684 36527 5733 36533
rect 5684 36524 5690 36527
rect 9122 36524 9128 36576
rect 9180 36564 9186 36576
rect 10428 36564 10456 36604
rect 9180 36536 10456 36564
rect 10505 36567 10563 36573
rect 9180 36524 9186 36536
rect 10505 36533 10517 36567
rect 10551 36564 10563 36567
rect 10594 36564 10600 36576
rect 10551 36536 10600 36564
rect 10551 36533 10563 36536
rect 10505 36527 10563 36533
rect 10594 36524 10600 36536
rect 10652 36524 10658 36576
rect 10704 36564 10732 36604
rect 12894 36592 12900 36604
rect 12952 36592 12958 36644
rect 11514 36564 11520 36576
rect 10704 36536 11520 36564
rect 11514 36524 11520 36536
rect 11572 36524 11578 36576
rect 13173 36567 13231 36573
rect 13173 36533 13185 36567
rect 13219 36564 13231 36567
rect 14384 36564 14412 36663
rect 17770 36660 17776 36712
rect 17828 36700 17834 36712
rect 17865 36703 17923 36709
rect 17865 36700 17877 36703
rect 17828 36672 17877 36700
rect 17828 36660 17834 36672
rect 17865 36669 17877 36672
rect 17911 36669 17923 36703
rect 17865 36663 17923 36669
rect 18969 36703 19027 36709
rect 18969 36669 18981 36703
rect 19015 36700 19027 36703
rect 19426 36700 19432 36712
rect 19015 36672 19432 36700
rect 19015 36669 19027 36672
rect 18969 36663 19027 36669
rect 17129 36635 17187 36641
rect 17129 36601 17141 36635
rect 17175 36632 17187 36635
rect 17880 36632 17908 36663
rect 19426 36660 19432 36672
rect 19484 36660 19490 36712
rect 23014 36660 23020 36712
rect 23072 36660 23078 36712
rect 24762 36660 24768 36712
rect 24820 36660 24826 36712
rect 17175 36604 17908 36632
rect 17175 36601 17187 36604
rect 17129 36595 17187 36601
rect 17954 36592 17960 36644
rect 18012 36632 18018 36644
rect 20622 36632 20628 36644
rect 18012 36604 20628 36632
rect 18012 36592 18018 36604
rect 20622 36592 20628 36604
rect 20680 36592 20686 36644
rect 13219 36536 14412 36564
rect 13219 36533 13231 36536
rect 13173 36527 13231 36533
rect 14550 36524 14556 36576
rect 14608 36564 14614 36576
rect 14829 36567 14887 36573
rect 14829 36564 14841 36567
rect 14608 36536 14841 36564
rect 14608 36524 14614 36536
rect 14829 36533 14841 36536
rect 14875 36533 14887 36567
rect 14829 36527 14887 36533
rect 15010 36524 15016 36576
rect 15068 36564 15074 36576
rect 17972 36564 18000 36592
rect 15068 36536 18000 36564
rect 15068 36524 15074 36536
rect 18782 36524 18788 36576
rect 18840 36564 18846 36576
rect 19334 36564 19340 36576
rect 18840 36536 19340 36564
rect 18840 36524 18846 36536
rect 19334 36524 19340 36536
rect 19392 36524 19398 36576
rect 1104 36474 40572 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 40572 36474
rect 1104 36400 40572 36422
rect 5442 36320 5448 36372
rect 5500 36360 5506 36372
rect 6457 36363 6515 36369
rect 6457 36360 6469 36363
rect 5500 36332 6469 36360
rect 5500 36320 5506 36332
rect 3970 36116 3976 36168
rect 4028 36116 4034 36168
rect 4249 36159 4307 36165
rect 4249 36125 4261 36159
rect 4295 36156 4307 36159
rect 4614 36156 4620 36168
rect 4295 36128 4620 36156
rect 4295 36125 4307 36128
rect 4249 36119 4307 36125
rect 4614 36116 4620 36128
rect 4672 36156 4678 36168
rect 5718 36156 5724 36168
rect 4672 36128 5724 36156
rect 4672 36116 4678 36128
rect 5718 36116 5724 36128
rect 5776 36116 5782 36168
rect 5828 36156 5856 36332
rect 6457 36329 6469 36332
rect 6503 36360 6515 36363
rect 7466 36360 7472 36372
rect 6503 36332 7472 36360
rect 6503 36329 6515 36332
rect 6457 36323 6515 36329
rect 7466 36320 7472 36332
rect 7524 36320 7530 36372
rect 7834 36320 7840 36372
rect 7892 36320 7898 36372
rect 7929 36363 7987 36369
rect 7929 36329 7941 36363
rect 7975 36360 7987 36363
rect 8570 36360 8576 36372
rect 7975 36332 8576 36360
rect 7975 36329 7987 36332
rect 7929 36323 7987 36329
rect 5905 36295 5963 36301
rect 5905 36261 5917 36295
rect 5951 36261 5963 36295
rect 5905 36255 5963 36261
rect 5920 36224 5948 36255
rect 5920 36196 6868 36224
rect 6089 36159 6147 36165
rect 6089 36156 6101 36159
rect 5828 36128 6101 36156
rect 6089 36125 6101 36128
rect 6135 36125 6147 36159
rect 6089 36119 6147 36125
rect 6181 36159 6239 36165
rect 6181 36125 6193 36159
rect 6227 36156 6239 36159
rect 6362 36156 6368 36168
rect 6227 36128 6368 36156
rect 6227 36125 6239 36128
rect 6181 36119 6239 36125
rect 6362 36116 6368 36128
rect 6420 36116 6426 36168
rect 3789 36091 3847 36097
rect 3789 36057 3801 36091
rect 3835 36088 3847 36091
rect 3835 36060 4292 36088
rect 3835 36057 3847 36060
rect 3789 36051 3847 36057
rect 4264 36032 4292 36060
rect 5810 36048 5816 36100
rect 5868 36088 5874 36100
rect 5905 36091 5963 36097
rect 5905 36088 5917 36091
rect 5868 36060 5917 36088
rect 5868 36048 5874 36060
rect 5905 36057 5917 36060
rect 5951 36088 5963 36091
rect 6270 36088 6276 36100
rect 5951 36060 6276 36088
rect 5951 36057 5963 36060
rect 5905 36051 5963 36057
rect 6270 36048 6276 36060
rect 6328 36048 6334 36100
rect 6380 36088 6408 36116
rect 6840 36097 6868 36196
rect 7282 36116 7288 36168
rect 7340 36116 7346 36168
rect 7653 36159 7711 36165
rect 7653 36125 7665 36159
rect 7699 36156 7711 36159
rect 7944 36156 7972 36323
rect 8570 36320 8576 36332
rect 8628 36320 8634 36372
rect 9217 36363 9275 36369
rect 9217 36329 9229 36363
rect 9263 36329 9275 36363
rect 9217 36323 9275 36329
rect 9401 36363 9459 36369
rect 9401 36329 9413 36363
rect 9447 36360 9459 36363
rect 12158 36360 12164 36372
rect 9447 36332 12164 36360
rect 9447 36329 9459 36332
rect 9401 36323 9459 36329
rect 9232 36292 9260 36323
rect 12158 36320 12164 36332
rect 12216 36320 12222 36372
rect 14734 36320 14740 36372
rect 14792 36360 14798 36372
rect 15749 36363 15807 36369
rect 15749 36360 15761 36363
rect 14792 36332 15761 36360
rect 14792 36320 14798 36332
rect 15749 36329 15761 36332
rect 15795 36329 15807 36363
rect 15749 36323 15807 36329
rect 18046 36320 18052 36372
rect 18104 36360 18110 36372
rect 18104 36332 21680 36360
rect 18104 36320 18110 36332
rect 9490 36292 9496 36304
rect 8404 36264 9496 36292
rect 8297 36227 8355 36233
rect 8297 36224 8309 36227
rect 7699 36128 7972 36156
rect 8036 36196 8309 36224
rect 7699 36125 7711 36128
rect 7653 36119 7711 36125
rect 6473 36091 6531 36097
rect 6473 36088 6485 36091
rect 6380 36060 6485 36088
rect 6473 36057 6485 36060
rect 6519 36057 6531 36091
rect 6473 36051 6531 36057
rect 6825 36091 6883 36097
rect 6825 36057 6837 36091
rect 6871 36057 6883 36091
rect 6825 36051 6883 36057
rect 7009 36091 7067 36097
rect 7009 36057 7021 36091
rect 7055 36057 7067 36091
rect 7009 36051 7067 36057
rect 7193 36091 7251 36097
rect 7193 36057 7205 36091
rect 7239 36088 7251 36091
rect 7469 36091 7527 36097
rect 7469 36088 7481 36091
rect 7239 36060 7481 36088
rect 7239 36057 7251 36060
rect 7193 36051 7251 36057
rect 7469 36057 7481 36060
rect 7515 36057 7527 36091
rect 7469 36051 7527 36057
rect 2958 35980 2964 36032
rect 3016 36020 3022 36032
rect 4157 36023 4215 36029
rect 4157 36020 4169 36023
rect 3016 35992 4169 36020
rect 3016 35980 3022 35992
rect 4157 35989 4169 35992
rect 4203 35989 4215 36023
rect 4157 35983 4215 35989
rect 4246 35980 4252 36032
rect 4304 35980 4310 36032
rect 6641 36023 6699 36029
rect 6641 35989 6653 36023
rect 6687 36020 6699 36023
rect 7024 36020 7052 36051
rect 7558 36048 7564 36100
rect 7616 36048 7622 36100
rect 7742 36048 7748 36100
rect 7800 36088 7806 36100
rect 8036 36088 8064 36196
rect 8297 36193 8309 36196
rect 8343 36193 8355 36227
rect 8297 36187 8355 36193
rect 8113 36159 8171 36165
rect 8113 36125 8125 36159
rect 8159 36156 8171 36159
rect 8202 36156 8208 36168
rect 8159 36128 8208 36156
rect 8159 36125 8171 36128
rect 8113 36119 8171 36125
rect 8202 36116 8208 36128
rect 8260 36116 8266 36168
rect 8404 36165 8432 36264
rect 9490 36252 9496 36264
rect 9548 36252 9554 36304
rect 13078 36252 13084 36304
rect 13136 36292 13142 36304
rect 13136 36264 14964 36292
rect 13136 36252 13142 36264
rect 8570 36184 8576 36236
rect 8628 36224 8634 36236
rect 8628 36196 9812 36224
rect 8628 36184 8634 36196
rect 8389 36159 8447 36165
rect 8389 36125 8401 36159
rect 8435 36125 8447 36159
rect 8389 36119 8447 36125
rect 9122 36116 9128 36168
rect 9180 36116 9186 36168
rect 9214 36116 9220 36168
rect 9272 36156 9278 36168
rect 9674 36156 9680 36168
rect 9272 36128 9680 36156
rect 9272 36116 9278 36128
rect 9674 36116 9680 36128
rect 9732 36116 9738 36168
rect 9784 36165 9812 36196
rect 9950 36184 9956 36236
rect 10008 36224 10014 36236
rect 10321 36227 10379 36233
rect 10321 36224 10333 36227
rect 10008 36196 10333 36224
rect 10008 36184 10014 36196
rect 10321 36193 10333 36196
rect 10367 36224 10379 36227
rect 10686 36224 10692 36236
rect 10367 36196 10692 36224
rect 10367 36193 10379 36196
rect 10321 36187 10379 36193
rect 10686 36184 10692 36196
rect 10744 36184 10750 36236
rect 11606 36184 11612 36236
rect 11664 36224 11670 36236
rect 11664 36196 11836 36224
rect 11664 36184 11670 36196
rect 9769 36159 9827 36165
rect 9769 36125 9781 36159
rect 9815 36125 9827 36159
rect 9769 36119 9827 36125
rect 10045 36159 10103 36165
rect 10045 36125 10057 36159
rect 10091 36125 10103 36159
rect 10045 36119 10103 36125
rect 10229 36159 10287 36165
rect 10229 36125 10241 36159
rect 10275 36125 10287 36159
rect 11808 36156 11836 36196
rect 11882 36184 11888 36236
rect 11940 36224 11946 36236
rect 11940 36196 12848 36224
rect 11940 36184 11946 36196
rect 11808 36128 11928 36156
rect 10229 36119 10287 36125
rect 8941 36091 8999 36097
rect 8941 36088 8953 36091
rect 7800 36060 8953 36088
rect 7800 36048 7806 36060
rect 8941 36057 8953 36060
rect 8987 36057 8999 36091
rect 10060 36088 10088 36119
rect 10134 36088 10140 36100
rect 8941 36051 8999 36057
rect 9508 36060 10140 36088
rect 9508 36020 9536 36060
rect 10134 36048 10140 36060
rect 10192 36048 10198 36100
rect 10244 36088 10272 36119
rect 10244 36060 10548 36088
rect 6687 35992 9536 36020
rect 9585 36023 9643 36029
rect 6687 35989 6699 35992
rect 6641 35983 6699 35989
rect 9585 35989 9597 36023
rect 9631 36020 9643 36023
rect 10410 36020 10416 36032
rect 9631 35992 10416 36020
rect 9631 35989 9643 35992
rect 9585 35983 9643 35989
rect 10410 35980 10416 35992
rect 10468 35980 10474 36032
rect 10520 36020 10548 36060
rect 10594 36048 10600 36100
rect 10652 36048 10658 36100
rect 10870 36048 10876 36100
rect 10928 36088 10934 36100
rect 10928 36060 11086 36088
rect 10928 36048 10934 36060
rect 11606 36020 11612 36032
rect 10520 35992 11612 36020
rect 11606 35980 11612 35992
rect 11664 35980 11670 36032
rect 11900 36020 11928 36128
rect 11974 36116 11980 36168
rect 12032 36156 12038 36168
rect 12345 36159 12403 36165
rect 12345 36156 12357 36159
rect 12032 36128 12357 36156
rect 12032 36116 12038 36128
rect 12345 36125 12357 36128
rect 12391 36156 12403 36159
rect 12391 36128 12664 36156
rect 12391 36125 12403 36128
rect 12345 36119 12403 36125
rect 12434 36048 12440 36100
rect 12492 36048 12498 36100
rect 12636 36088 12664 36128
rect 12710 36116 12716 36168
rect 12768 36116 12774 36168
rect 12820 36165 12848 36196
rect 14550 36184 14556 36236
rect 14608 36184 14614 36236
rect 14737 36227 14795 36233
rect 14737 36193 14749 36227
rect 14783 36224 14795 36227
rect 14826 36224 14832 36236
rect 14783 36196 14832 36224
rect 14783 36193 14795 36196
rect 14737 36187 14795 36193
rect 14826 36184 14832 36196
rect 14884 36184 14890 36236
rect 14936 36233 14964 36264
rect 15286 36252 15292 36304
rect 15344 36252 15350 36304
rect 15654 36292 15660 36304
rect 15580 36264 15660 36292
rect 14921 36227 14979 36233
rect 14921 36193 14933 36227
rect 14967 36224 14979 36227
rect 15194 36224 15200 36236
rect 14967 36196 15200 36224
rect 14967 36193 14979 36196
rect 14921 36187 14979 36193
rect 15194 36184 15200 36196
rect 15252 36224 15258 36236
rect 15252 36196 15516 36224
rect 15252 36184 15258 36196
rect 12805 36159 12863 36165
rect 12805 36125 12817 36159
rect 12851 36125 12863 36159
rect 12805 36119 12863 36125
rect 15105 36159 15163 36165
rect 15105 36125 15117 36159
rect 15151 36125 15163 36159
rect 15105 36119 15163 36125
rect 12989 36091 13047 36097
rect 12636 36060 12940 36088
rect 12621 36023 12679 36029
rect 12621 36020 12633 36023
rect 11900 35992 12633 36020
rect 12621 35989 12633 35992
rect 12667 35989 12679 36023
rect 12912 36020 12940 36060
rect 12989 36057 13001 36091
rect 13035 36088 13047 36091
rect 13538 36088 13544 36100
rect 13035 36060 13544 36088
rect 13035 36057 13047 36060
rect 12989 36051 13047 36057
rect 13538 36048 13544 36060
rect 13596 36088 13602 36100
rect 15120 36088 15148 36119
rect 13596 36060 15148 36088
rect 15488 36088 15516 36196
rect 15580 36165 15608 36264
rect 15654 36252 15660 36264
rect 15712 36252 15718 36304
rect 21545 36295 21603 36301
rect 21545 36261 21557 36295
rect 21591 36261 21603 36295
rect 21545 36255 21603 36261
rect 15838 36184 15844 36236
rect 15896 36224 15902 36236
rect 17218 36224 17224 36236
rect 15896 36196 17224 36224
rect 15896 36184 15902 36196
rect 17218 36184 17224 36196
rect 17276 36184 17282 36236
rect 18782 36224 18788 36236
rect 18156 36196 18788 36224
rect 15565 36159 15623 36165
rect 15565 36125 15577 36159
rect 15611 36125 15623 36159
rect 15565 36119 15623 36125
rect 15657 36159 15715 36165
rect 15657 36125 15669 36159
rect 15703 36156 15715 36159
rect 15703 36128 16252 36156
rect 15703 36125 15715 36128
rect 15657 36119 15715 36125
rect 16114 36088 16120 36100
rect 15488 36060 16120 36088
rect 13596 36048 13602 36060
rect 16114 36048 16120 36060
rect 16172 36048 16178 36100
rect 13354 36020 13360 36032
rect 12912 35992 13360 36020
rect 12621 35983 12679 35989
rect 13354 35980 13360 35992
rect 13412 35980 13418 36032
rect 13722 35980 13728 36032
rect 13780 36020 13786 36032
rect 14093 36023 14151 36029
rect 14093 36020 14105 36023
rect 13780 35992 14105 36020
rect 13780 35980 13786 35992
rect 14093 35989 14105 35992
rect 14139 35989 14151 36023
rect 14093 35983 14151 35989
rect 14461 36023 14519 36029
rect 14461 35989 14473 36023
rect 14507 36020 14519 36023
rect 15470 36020 15476 36032
rect 14507 35992 15476 36020
rect 14507 35989 14519 35992
rect 14461 35983 14519 35989
rect 15470 35980 15476 35992
rect 15528 35980 15534 36032
rect 15838 35980 15844 36032
rect 15896 36020 15902 36032
rect 16224 36020 16252 36128
rect 16390 36116 16396 36168
rect 16448 36156 16454 36168
rect 18156 36165 18184 36196
rect 18782 36184 18788 36196
rect 18840 36184 18846 36236
rect 19242 36184 19248 36236
rect 19300 36224 19306 36236
rect 21560 36224 21588 36255
rect 19300 36196 21588 36224
rect 19300 36184 19306 36196
rect 18141 36159 18199 36165
rect 18141 36156 18153 36159
rect 16448 36128 18153 36156
rect 16448 36116 16454 36128
rect 18141 36125 18153 36128
rect 18187 36125 18199 36159
rect 18141 36119 18199 36125
rect 18230 36116 18236 36168
rect 18288 36156 18294 36168
rect 18325 36159 18383 36165
rect 18325 36156 18337 36159
rect 18288 36128 18337 36156
rect 18288 36116 18294 36128
rect 18325 36125 18337 36128
rect 18371 36125 18383 36159
rect 18325 36119 18383 36125
rect 19610 36116 19616 36168
rect 19668 36116 19674 36168
rect 16298 36048 16304 36100
rect 16356 36088 16362 36100
rect 16356 36060 18368 36088
rect 16356 36048 16362 36060
rect 17126 36020 17132 36032
rect 15896 35992 17132 36020
rect 15896 35980 15902 35992
rect 17126 35980 17132 35992
rect 17184 35980 17190 36032
rect 17954 35980 17960 36032
rect 18012 36020 18018 36032
rect 18233 36023 18291 36029
rect 18233 36020 18245 36023
rect 18012 35992 18245 36020
rect 18012 35980 18018 35992
rect 18233 35989 18245 35992
rect 18279 35989 18291 36023
rect 18340 36020 18368 36060
rect 19886 36048 19892 36100
rect 19944 36048 19950 36100
rect 20622 36048 20628 36100
rect 20680 36048 20686 36100
rect 21652 36088 21680 36332
rect 24136 36264 25268 36292
rect 24136 36233 24164 36264
rect 22005 36227 22063 36233
rect 22005 36193 22017 36227
rect 22051 36224 22063 36227
rect 22373 36227 22431 36233
rect 22373 36224 22385 36227
rect 22051 36196 22385 36224
rect 22051 36193 22063 36196
rect 22005 36187 22063 36193
rect 22373 36193 22385 36196
rect 22419 36193 22431 36227
rect 22373 36187 22431 36193
rect 24121 36227 24179 36233
rect 24121 36193 24133 36227
rect 24167 36193 24179 36227
rect 24121 36187 24179 36193
rect 24762 36184 24768 36236
rect 24820 36224 24826 36236
rect 25133 36227 25191 36233
rect 25133 36224 25145 36227
rect 24820 36196 25145 36224
rect 24820 36184 24826 36196
rect 25133 36193 25145 36196
rect 25179 36193 25191 36227
rect 25240 36224 25268 36264
rect 25774 36224 25780 36236
rect 25240 36196 25780 36224
rect 25133 36187 25191 36193
rect 25774 36184 25780 36196
rect 25832 36224 25838 36236
rect 25958 36224 25964 36236
rect 25832 36196 25964 36224
rect 25832 36184 25838 36196
rect 25958 36184 25964 36196
rect 26016 36184 26022 36236
rect 27154 36184 27160 36236
rect 27212 36224 27218 36236
rect 28350 36224 28356 36236
rect 27212 36196 28356 36224
rect 27212 36184 27218 36196
rect 28350 36184 28356 36196
rect 28408 36184 28414 36236
rect 21910 36116 21916 36168
rect 21968 36116 21974 36168
rect 22278 36116 22284 36168
rect 22336 36116 22342 36168
rect 22462 36116 22468 36168
rect 22520 36116 22526 36168
rect 23014 36116 23020 36168
rect 23072 36156 23078 36168
rect 23293 36159 23351 36165
rect 23293 36156 23305 36159
rect 23072 36128 23305 36156
rect 23072 36116 23078 36128
rect 23293 36125 23305 36128
rect 23339 36156 23351 36159
rect 24780 36156 24808 36184
rect 23339 36128 24808 36156
rect 23339 36125 23351 36128
rect 23293 36119 23351 36125
rect 23845 36091 23903 36097
rect 23845 36088 23857 36091
rect 21284 36060 21496 36088
rect 21652 36060 23857 36088
rect 21284 36020 21312 36060
rect 18340 35992 21312 36020
rect 18233 35983 18291 35989
rect 21358 35980 21364 36032
rect 21416 35980 21422 36032
rect 21468 36020 21496 36060
rect 23845 36057 23857 36060
rect 23891 36057 23903 36091
rect 23845 36051 23903 36057
rect 23937 36091 23995 36097
rect 23937 36057 23949 36091
rect 23983 36088 23995 36091
rect 25130 36088 25136 36100
rect 23983 36060 25136 36088
rect 23983 36057 23995 36060
rect 23937 36051 23995 36057
rect 25130 36048 25136 36060
rect 25188 36048 25194 36100
rect 25406 36048 25412 36100
rect 25464 36048 25470 36100
rect 30466 36088 30472 36100
rect 26634 36060 30472 36088
rect 30466 36048 30472 36060
rect 30524 36048 30530 36100
rect 22554 36020 22560 36032
rect 21468 35992 22560 36020
rect 22554 35980 22560 35992
rect 22612 35980 22618 36032
rect 23474 35980 23480 36032
rect 23532 35980 23538 36032
rect 1104 35930 40572 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 40572 35930
rect 1104 35856 40572 35878
rect 5626 35776 5632 35828
rect 5684 35816 5690 35828
rect 5994 35816 6000 35828
rect 5684 35788 6000 35816
rect 5684 35776 5690 35788
rect 5994 35776 6000 35788
rect 6052 35816 6058 35828
rect 6365 35819 6423 35825
rect 6365 35816 6377 35819
rect 6052 35788 6377 35816
rect 6052 35776 6058 35788
rect 6365 35785 6377 35788
rect 6411 35785 6423 35819
rect 6365 35779 6423 35785
rect 7558 35776 7564 35828
rect 7616 35776 7622 35828
rect 8846 35776 8852 35828
rect 8904 35776 8910 35828
rect 9030 35776 9036 35828
rect 9088 35776 9094 35828
rect 10781 35819 10839 35825
rect 10781 35785 10793 35819
rect 10827 35816 10839 35819
rect 10827 35788 10916 35816
rect 10827 35785 10839 35788
rect 10781 35779 10839 35785
rect 1302 35708 1308 35760
rect 1360 35748 1366 35760
rect 2317 35751 2375 35757
rect 2317 35748 2329 35751
rect 1360 35720 2329 35748
rect 1360 35708 1366 35720
rect 2317 35717 2329 35720
rect 2363 35717 2375 35751
rect 2317 35711 2375 35717
rect 2501 35751 2559 35757
rect 2501 35717 2513 35751
rect 2547 35748 2559 35751
rect 2958 35748 2964 35760
rect 2547 35720 2964 35748
rect 2547 35717 2559 35720
rect 2501 35711 2559 35717
rect 2958 35708 2964 35720
rect 3016 35708 3022 35760
rect 3786 35708 3792 35760
rect 3844 35708 3850 35760
rect 4246 35708 4252 35760
rect 4304 35708 4310 35760
rect 5442 35708 5448 35760
rect 5500 35748 5506 35760
rect 7101 35751 7159 35757
rect 7101 35748 7113 35751
rect 5500 35720 7113 35748
rect 5500 35708 5506 35720
rect 7101 35717 7113 35720
rect 7147 35748 7159 35751
rect 8018 35748 8024 35760
rect 7147 35720 8024 35748
rect 7147 35717 7159 35720
rect 7101 35711 7159 35717
rect 8018 35708 8024 35720
rect 8076 35748 8082 35760
rect 8076 35720 8524 35748
rect 8076 35708 8082 35720
rect 2133 35683 2191 35689
rect 2133 35649 2145 35683
rect 2179 35649 2191 35683
rect 2133 35643 2191 35649
rect 2148 35612 2176 35643
rect 2222 35640 2228 35692
rect 2280 35680 2286 35692
rect 2409 35683 2467 35689
rect 2409 35680 2421 35683
rect 2280 35652 2421 35680
rect 2280 35640 2286 35652
rect 2409 35649 2421 35652
rect 2455 35649 2467 35683
rect 2409 35643 2467 35649
rect 4525 35683 4583 35689
rect 4525 35649 4537 35683
rect 4571 35680 4583 35683
rect 5534 35680 5540 35692
rect 4571 35652 5540 35680
rect 4571 35649 4583 35652
rect 4525 35643 4583 35649
rect 5534 35640 5540 35652
rect 5592 35640 5598 35692
rect 5997 35683 6055 35689
rect 5997 35649 6009 35683
rect 6043 35649 6055 35683
rect 5997 35643 6055 35649
rect 5810 35612 5816 35624
rect 2148 35584 5816 35612
rect 5810 35572 5816 35584
rect 5868 35572 5874 35624
rect 1949 35479 2007 35485
rect 1949 35445 1961 35479
rect 1995 35476 2007 35479
rect 3142 35476 3148 35488
rect 1995 35448 3148 35476
rect 1995 35445 2007 35448
rect 1949 35439 2007 35445
rect 3142 35436 3148 35448
rect 3200 35436 3206 35488
rect 5810 35436 5816 35488
rect 5868 35476 5874 35488
rect 6012 35476 6040 35643
rect 6178 35640 6184 35692
rect 6236 35680 6242 35692
rect 6549 35683 6607 35689
rect 6549 35680 6561 35683
rect 6236 35652 6561 35680
rect 6236 35640 6242 35652
rect 6549 35649 6561 35652
rect 6595 35649 6607 35683
rect 6917 35683 6975 35689
rect 6917 35680 6929 35683
rect 6549 35643 6607 35649
rect 6656 35652 6929 35680
rect 6089 35547 6147 35553
rect 6089 35513 6101 35547
rect 6135 35544 6147 35547
rect 6546 35544 6552 35556
rect 6135 35516 6552 35544
rect 6135 35513 6147 35516
rect 6089 35507 6147 35513
rect 6546 35504 6552 35516
rect 6604 35504 6610 35556
rect 6656 35476 6684 35652
rect 6917 35649 6929 35652
rect 6963 35680 6975 35683
rect 7006 35680 7012 35692
rect 6963 35652 7012 35680
rect 6963 35649 6975 35652
rect 6917 35643 6975 35649
rect 7006 35640 7012 35652
rect 7064 35640 7070 35692
rect 7469 35683 7527 35689
rect 7469 35649 7481 35683
rect 7515 35680 7527 35683
rect 7558 35680 7564 35692
rect 7515 35652 7564 35680
rect 7515 35649 7527 35652
rect 7469 35643 7527 35649
rect 7558 35640 7564 35652
rect 7616 35640 7622 35692
rect 7653 35683 7711 35689
rect 7653 35649 7665 35683
rect 7699 35680 7711 35683
rect 7742 35680 7748 35692
rect 7699 35652 7748 35680
rect 7699 35649 7711 35652
rect 7653 35643 7711 35649
rect 7742 35640 7748 35652
rect 7800 35640 7806 35692
rect 8496 35689 8524 35720
rect 8570 35708 8576 35760
rect 8628 35748 8634 35760
rect 10594 35748 10600 35760
rect 8628 35720 10600 35748
rect 8628 35708 8634 35720
rect 10594 35708 10600 35720
rect 10652 35708 10658 35760
rect 10888 35748 10916 35788
rect 11054 35776 11060 35828
rect 11112 35816 11118 35828
rect 11882 35816 11888 35828
rect 11112 35788 11888 35816
rect 11112 35776 11118 35788
rect 11882 35776 11888 35788
rect 11940 35776 11946 35828
rect 12069 35819 12127 35825
rect 12069 35785 12081 35819
rect 12115 35816 12127 35819
rect 12526 35816 12532 35828
rect 12115 35788 12532 35816
rect 12115 35785 12127 35788
rect 12069 35779 12127 35785
rect 12526 35776 12532 35788
rect 12584 35816 12590 35828
rect 16298 35816 16304 35828
rect 12584 35788 15700 35816
rect 12584 35776 12590 35788
rect 11149 35751 11207 35757
rect 11149 35748 11161 35751
rect 10888 35720 11161 35748
rect 11149 35717 11161 35720
rect 11195 35717 11207 35751
rect 11149 35711 11207 35717
rect 11514 35708 11520 35760
rect 11572 35748 11578 35760
rect 11609 35751 11667 35757
rect 11609 35748 11621 35751
rect 11572 35720 11621 35748
rect 11572 35708 11578 35720
rect 11609 35717 11621 35720
rect 11655 35717 11667 35751
rect 11609 35711 11667 35717
rect 8481 35683 8539 35689
rect 8481 35649 8493 35683
rect 8527 35649 8539 35683
rect 8481 35643 8539 35649
rect 8665 35683 8723 35689
rect 8665 35649 8677 35683
rect 8711 35680 8723 35683
rect 9030 35680 9036 35692
rect 8711 35652 9036 35680
rect 8711 35649 8723 35652
rect 8665 35643 8723 35649
rect 6730 35572 6736 35624
rect 6788 35612 6794 35624
rect 6825 35615 6883 35621
rect 6825 35612 6837 35615
rect 6788 35584 6837 35612
rect 6788 35572 6794 35584
rect 6825 35581 6837 35584
rect 6871 35581 6883 35615
rect 6825 35575 6883 35581
rect 8386 35572 8392 35624
rect 8444 35612 8450 35624
rect 8680 35612 8708 35643
rect 9030 35640 9036 35652
rect 9088 35640 9094 35692
rect 9217 35683 9275 35689
rect 9217 35649 9229 35683
rect 9263 35649 9275 35683
rect 9217 35643 9275 35649
rect 8444 35584 8708 35612
rect 9232 35612 9260 35643
rect 9306 35640 9312 35692
rect 9364 35640 9370 35692
rect 9398 35640 9404 35692
rect 9456 35680 9462 35692
rect 9493 35683 9551 35689
rect 9493 35680 9505 35683
rect 9456 35652 9505 35680
rect 9456 35640 9462 35652
rect 9493 35649 9505 35652
rect 9539 35649 9551 35683
rect 9493 35643 9551 35649
rect 9674 35640 9680 35692
rect 9732 35680 9738 35692
rect 10502 35680 10508 35692
rect 9732 35652 10508 35680
rect 9732 35640 9738 35652
rect 10502 35640 10508 35652
rect 10560 35640 10566 35692
rect 10864 35683 10922 35689
rect 10864 35680 10876 35683
rect 10842 35678 10876 35680
rect 10704 35650 10876 35678
rect 9232 35584 9444 35612
rect 8444 35572 8450 35584
rect 7374 35544 7380 35556
rect 6748 35516 7380 35544
rect 6748 35485 6776 35516
rect 7374 35504 7380 35516
rect 7432 35504 7438 35556
rect 5868 35448 6684 35476
rect 6733 35479 6791 35485
rect 5868 35436 5874 35448
rect 6733 35445 6745 35479
rect 6779 35445 6791 35479
rect 6733 35439 6791 35445
rect 7190 35436 7196 35488
rect 7248 35476 7254 35488
rect 7285 35479 7343 35485
rect 7285 35476 7297 35479
rect 7248 35448 7297 35476
rect 7248 35436 7254 35448
rect 7285 35445 7297 35448
rect 7331 35445 7343 35479
rect 7285 35439 7343 35445
rect 9122 35436 9128 35488
rect 9180 35476 9186 35488
rect 9309 35479 9367 35485
rect 9309 35476 9321 35479
rect 9180 35448 9321 35476
rect 9180 35436 9186 35448
rect 9309 35445 9321 35448
rect 9355 35445 9367 35479
rect 9416 35476 9444 35584
rect 10410 35572 10416 35624
rect 10468 35612 10474 35624
rect 10597 35615 10655 35621
rect 10597 35612 10609 35615
rect 10468 35584 10609 35612
rect 10468 35572 10474 35584
rect 10597 35581 10609 35584
rect 10643 35612 10655 35615
rect 10704 35612 10732 35650
rect 10864 35649 10876 35650
rect 10910 35649 10922 35683
rect 10864 35643 10922 35649
rect 10962 35640 10968 35692
rect 11020 35640 11026 35692
rect 11698 35640 11704 35692
rect 11756 35640 11762 35692
rect 11900 35689 11928 35776
rect 13814 35748 13820 35760
rect 13464 35720 13820 35748
rect 11885 35683 11943 35689
rect 11885 35649 11897 35683
rect 11931 35649 11943 35683
rect 11885 35643 11943 35649
rect 12069 35683 12127 35689
rect 12069 35649 12081 35683
rect 12115 35680 12127 35683
rect 12434 35680 12440 35692
rect 12115 35652 12440 35680
rect 12115 35649 12127 35652
rect 12069 35643 12127 35649
rect 10643 35584 10732 35612
rect 10781 35615 10839 35621
rect 10643 35581 10655 35584
rect 10597 35575 10655 35581
rect 10781 35581 10793 35615
rect 10827 35581 10839 35615
rect 10980 35612 11008 35640
rect 12084 35612 12112 35643
rect 12434 35640 12440 35652
rect 12492 35680 12498 35692
rect 12802 35680 12808 35692
rect 12492 35652 12808 35680
rect 12492 35640 12498 35652
rect 12802 35640 12808 35652
rect 12860 35640 12866 35692
rect 13464 35689 13492 35720
rect 13814 35708 13820 35720
rect 13872 35708 13878 35760
rect 15010 35748 15016 35760
rect 14950 35720 15016 35748
rect 15010 35708 15016 35720
rect 15068 35708 15074 35760
rect 13449 35683 13507 35689
rect 13449 35649 13461 35683
rect 13495 35649 13507 35683
rect 13449 35643 13507 35649
rect 15102 35640 15108 35692
rect 15160 35680 15166 35692
rect 15672 35689 15700 35788
rect 15764 35788 16304 35816
rect 15764 35689 15792 35788
rect 16298 35776 16304 35788
rect 16356 35776 16362 35828
rect 17310 35776 17316 35828
rect 17368 35816 17374 35828
rect 17368 35788 18460 35816
rect 17368 35776 17374 35788
rect 17221 35751 17279 35757
rect 17221 35717 17233 35751
rect 17267 35748 17279 35751
rect 17954 35748 17960 35760
rect 17267 35720 17960 35748
rect 17267 35717 17279 35720
rect 17221 35711 17279 35717
rect 17954 35708 17960 35720
rect 18012 35708 18018 35760
rect 15657 35683 15715 35689
rect 15160 35652 15608 35680
rect 15160 35640 15166 35652
rect 10980 35584 12112 35612
rect 10781 35575 10839 35581
rect 10134 35476 10140 35488
rect 9416 35448 10140 35476
rect 9309 35439 9367 35445
rect 10134 35436 10140 35448
rect 10192 35436 10198 35488
rect 10594 35436 10600 35488
rect 10652 35476 10658 35488
rect 10796 35476 10824 35575
rect 13722 35572 13728 35624
rect 13780 35572 13786 35624
rect 15470 35572 15476 35624
rect 15528 35572 15534 35624
rect 15580 35612 15608 35652
rect 15657 35649 15669 35683
rect 15703 35649 15715 35683
rect 15657 35643 15715 35649
rect 15749 35683 15807 35689
rect 15749 35649 15761 35683
rect 15795 35649 15807 35683
rect 15749 35643 15807 35649
rect 15764 35612 15792 35643
rect 15838 35640 15844 35692
rect 15896 35640 15902 35692
rect 15933 35683 15991 35689
rect 15933 35649 15945 35683
rect 15979 35680 15991 35683
rect 16022 35680 16028 35692
rect 15979 35652 16028 35680
rect 15979 35649 15991 35652
rect 15933 35643 15991 35649
rect 16022 35640 16028 35652
rect 16080 35640 16086 35692
rect 17129 35683 17187 35689
rect 17129 35649 17141 35683
rect 17175 35649 17187 35683
rect 17129 35643 17187 35649
rect 17405 35683 17463 35689
rect 17405 35649 17417 35683
rect 17451 35680 17463 35683
rect 17494 35680 17500 35692
rect 17451 35652 17500 35680
rect 17451 35649 17463 35652
rect 17405 35643 17463 35649
rect 15580 35584 15792 35612
rect 16114 35572 16120 35624
rect 16172 35572 16178 35624
rect 16666 35572 16672 35624
rect 16724 35612 16730 35624
rect 17144 35612 17172 35643
rect 17494 35640 17500 35652
rect 17552 35640 17558 35692
rect 17589 35683 17647 35689
rect 17589 35649 17601 35683
rect 17635 35680 17647 35683
rect 18325 35683 18383 35689
rect 18325 35680 18337 35683
rect 17635 35652 18337 35680
rect 17635 35649 17647 35652
rect 17589 35643 17647 35649
rect 18325 35649 18337 35652
rect 18371 35649 18383 35683
rect 18432 35680 18460 35788
rect 18506 35776 18512 35828
rect 18564 35816 18570 35828
rect 19058 35816 19064 35828
rect 18564 35788 19064 35816
rect 18564 35776 18570 35788
rect 19058 35776 19064 35788
rect 19116 35816 19122 35828
rect 19426 35816 19432 35828
rect 19116 35788 19432 35816
rect 19116 35776 19122 35788
rect 19426 35776 19432 35788
rect 19484 35776 19490 35828
rect 19797 35819 19855 35825
rect 19797 35785 19809 35819
rect 19843 35816 19855 35819
rect 19886 35816 19892 35828
rect 19843 35788 19892 35816
rect 19843 35785 19855 35788
rect 19797 35779 19855 35785
rect 19886 35776 19892 35788
rect 19944 35776 19950 35828
rect 21177 35819 21235 35825
rect 21177 35785 21189 35819
rect 21223 35816 21235 35819
rect 22462 35816 22468 35828
rect 21223 35788 22468 35816
rect 21223 35785 21235 35788
rect 21177 35779 21235 35785
rect 21358 35748 21364 35760
rect 19628 35720 21364 35748
rect 18506 35680 18512 35692
rect 18432 35652 18512 35680
rect 18325 35643 18383 35649
rect 18506 35640 18512 35652
rect 18564 35640 18570 35692
rect 19061 35683 19119 35689
rect 19061 35649 19073 35683
rect 19107 35649 19119 35683
rect 19061 35643 19119 35649
rect 17865 35615 17923 35621
rect 17865 35612 17877 35615
rect 16724 35584 17877 35612
rect 16724 35572 16730 35584
rect 17865 35581 17877 35584
rect 17911 35581 17923 35615
rect 17865 35575 17923 35581
rect 17954 35572 17960 35624
rect 18012 35572 18018 35624
rect 18046 35572 18052 35624
rect 18104 35572 18110 35624
rect 18141 35615 18199 35621
rect 18141 35581 18153 35615
rect 18187 35612 18199 35615
rect 18417 35615 18475 35621
rect 18417 35612 18429 35615
rect 18187 35584 18429 35612
rect 18187 35581 18199 35584
rect 18141 35575 18199 35581
rect 18417 35581 18429 35584
rect 18463 35581 18475 35615
rect 18417 35575 18475 35581
rect 11146 35504 11152 35556
rect 11204 35504 11210 35556
rect 15488 35544 15516 35572
rect 16206 35544 16212 35556
rect 15488 35516 16212 35544
rect 16206 35504 16212 35516
rect 16264 35504 16270 35556
rect 16298 35504 16304 35556
rect 16356 35544 16362 35556
rect 17402 35544 17408 35556
rect 16356 35516 17408 35544
rect 16356 35504 16362 35516
rect 17402 35504 17408 35516
rect 17460 35504 17466 35556
rect 17681 35547 17739 35553
rect 17681 35513 17693 35547
rect 17727 35544 17739 35547
rect 19076 35544 19104 35643
rect 19242 35640 19248 35692
rect 19300 35640 19306 35692
rect 19426 35640 19432 35692
rect 19484 35640 19490 35692
rect 19518 35640 19524 35692
rect 19576 35680 19582 35692
rect 19628 35689 19656 35720
rect 19613 35683 19671 35689
rect 19613 35680 19625 35683
rect 19576 35652 19625 35680
rect 19576 35640 19582 35652
rect 19613 35649 19625 35652
rect 19659 35649 19671 35683
rect 19613 35643 19671 35649
rect 19794 35640 19800 35692
rect 19852 35680 19858 35692
rect 21192 35689 21220 35720
rect 21358 35708 21364 35720
rect 21416 35708 21422 35760
rect 21560 35689 21588 35788
rect 22462 35776 22468 35788
rect 22520 35776 22526 35828
rect 23474 35816 23480 35828
rect 23308 35788 23480 35816
rect 21910 35748 21916 35760
rect 21652 35720 21916 35748
rect 21652 35689 21680 35720
rect 21910 35708 21916 35720
rect 21968 35708 21974 35760
rect 23308 35757 23336 35788
rect 23474 35776 23480 35788
rect 23532 35776 23538 35828
rect 25317 35819 25375 35825
rect 25317 35785 25329 35819
rect 25363 35816 25375 35819
rect 25406 35816 25412 35828
rect 25363 35788 25412 35816
rect 25363 35785 25375 35788
rect 25317 35779 25375 35785
rect 25406 35776 25412 35788
rect 25464 35776 25470 35828
rect 25777 35819 25835 35825
rect 25777 35785 25789 35819
rect 25823 35816 25835 35819
rect 27154 35816 27160 35828
rect 25823 35788 27160 35816
rect 25823 35785 25835 35788
rect 25777 35779 25835 35785
rect 27154 35776 27160 35788
rect 27212 35776 27218 35828
rect 23293 35751 23351 35757
rect 23293 35717 23305 35751
rect 23339 35717 23351 35751
rect 24946 35748 24952 35760
rect 24518 35720 24952 35748
rect 23293 35711 23351 35717
rect 24946 35708 24952 35720
rect 25004 35708 25010 35760
rect 25041 35751 25099 35757
rect 25041 35717 25053 35751
rect 25087 35748 25099 35751
rect 25130 35748 25136 35760
rect 25087 35720 25136 35748
rect 25087 35717 25099 35720
rect 25041 35711 25099 35717
rect 25130 35708 25136 35720
rect 25188 35708 25194 35760
rect 20993 35683 21051 35689
rect 20993 35680 21005 35683
rect 19852 35652 21005 35680
rect 19852 35640 19858 35652
rect 20993 35649 21005 35652
rect 21039 35649 21051 35683
rect 20993 35643 21051 35649
rect 21177 35683 21235 35689
rect 21177 35649 21189 35683
rect 21223 35649 21235 35683
rect 21177 35643 21235 35649
rect 21544 35683 21602 35689
rect 21544 35649 21556 35683
rect 21590 35649 21602 35683
rect 21544 35643 21602 35649
rect 21637 35683 21695 35689
rect 21637 35649 21649 35683
rect 21683 35649 21695 35683
rect 21637 35643 21695 35649
rect 21821 35683 21879 35689
rect 21821 35649 21833 35683
rect 21867 35680 21879 35683
rect 22002 35680 22008 35692
rect 21867 35652 22008 35680
rect 21867 35649 21879 35652
rect 21821 35643 21879 35649
rect 19150 35572 19156 35624
rect 19208 35612 19214 35624
rect 19337 35615 19395 35621
rect 19337 35612 19349 35615
rect 19208 35584 19349 35612
rect 19208 35572 19214 35584
rect 19337 35581 19349 35584
rect 19383 35581 19395 35615
rect 21008 35612 21036 35643
rect 22002 35640 22008 35652
rect 22060 35640 22066 35692
rect 23014 35640 23020 35692
rect 23072 35640 23078 35692
rect 25685 35683 25743 35689
rect 25685 35649 25697 35683
rect 25731 35649 25743 35683
rect 25685 35643 25743 35649
rect 21266 35612 21272 35624
rect 21008 35584 21272 35612
rect 19337 35575 19395 35581
rect 21266 35572 21272 35584
rect 21324 35572 21330 35624
rect 22557 35615 22615 35621
rect 22557 35612 22569 35615
rect 22066 35584 22569 35612
rect 17727 35516 19104 35544
rect 21376 35516 21588 35544
rect 17727 35513 17739 35516
rect 17681 35507 17739 35513
rect 11238 35476 11244 35488
rect 10652 35448 11244 35476
rect 10652 35436 10658 35448
rect 11238 35436 11244 35448
rect 11296 35436 11302 35488
rect 13538 35436 13544 35488
rect 13596 35476 13602 35488
rect 14734 35476 14740 35488
rect 13596 35448 14740 35476
rect 13596 35436 13602 35448
rect 14734 35436 14740 35448
rect 14792 35476 14798 35488
rect 15838 35476 15844 35488
rect 14792 35448 15844 35476
rect 14792 35436 14798 35448
rect 15838 35436 15844 35448
rect 15896 35436 15902 35488
rect 18230 35436 18236 35488
rect 18288 35476 18294 35488
rect 21376 35476 21404 35516
rect 18288 35448 21404 35476
rect 18288 35436 18294 35448
rect 21450 35436 21456 35488
rect 21508 35436 21514 35488
rect 21560 35476 21588 35516
rect 21634 35504 21640 35556
rect 21692 35544 21698 35556
rect 22066 35544 22094 35584
rect 22557 35581 22569 35584
rect 22603 35581 22615 35615
rect 22557 35575 22615 35581
rect 21692 35516 22094 35544
rect 21692 35504 21698 35516
rect 25700 35476 25728 35643
rect 25866 35572 25872 35624
rect 25924 35572 25930 35624
rect 21560 35448 25728 35476
rect 1104 35386 40572 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 40572 35386
rect 1104 35312 40572 35334
rect 4157 35275 4215 35281
rect 4157 35241 4169 35275
rect 4203 35272 4215 35275
rect 5442 35272 5448 35284
rect 4203 35244 5448 35272
rect 4203 35241 4215 35244
rect 4157 35235 4215 35241
rect 5442 35232 5448 35244
rect 5500 35232 5506 35284
rect 6730 35232 6736 35284
rect 6788 35272 6794 35284
rect 7377 35275 7435 35281
rect 7377 35272 7389 35275
rect 6788 35244 7389 35272
rect 6788 35232 6794 35244
rect 7377 35241 7389 35244
rect 7423 35241 7435 35275
rect 7377 35235 7435 35241
rect 7742 35232 7748 35284
rect 7800 35232 7806 35284
rect 8205 35275 8263 35281
rect 8205 35241 8217 35275
rect 8251 35272 8263 35275
rect 9306 35272 9312 35284
rect 8251 35244 9312 35272
rect 8251 35241 8263 35244
rect 8205 35235 8263 35241
rect 9306 35232 9312 35244
rect 9364 35232 9370 35284
rect 16114 35232 16120 35284
rect 16172 35272 16178 35284
rect 16209 35275 16267 35281
rect 16209 35272 16221 35275
rect 16172 35244 16221 35272
rect 16172 35232 16178 35244
rect 16209 35241 16221 35244
rect 16255 35241 16267 35275
rect 16209 35235 16267 35241
rect 16666 35232 16672 35284
rect 16724 35232 16730 35284
rect 16776 35244 18460 35272
rect 7009 35207 7067 35213
rect 7009 35173 7021 35207
rect 7055 35204 7067 35207
rect 8941 35207 8999 35213
rect 8941 35204 8953 35207
rect 7055 35176 8953 35204
rect 7055 35173 7067 35176
rect 7009 35167 7067 35173
rect 8941 35173 8953 35176
rect 8987 35173 8999 35207
rect 8941 35167 8999 35173
rect 9030 35164 9036 35216
rect 9088 35204 9094 35216
rect 9088 35176 9352 35204
rect 9088 35164 9094 35176
rect 3142 35096 3148 35148
rect 3200 35096 3206 35148
rect 3421 35139 3479 35145
rect 3421 35105 3433 35139
rect 3467 35136 3479 35139
rect 5534 35136 5540 35148
rect 3467 35108 5540 35136
rect 3467 35105 3479 35108
rect 3421 35099 3479 35105
rect 5534 35096 5540 35108
rect 5592 35136 5598 35148
rect 5905 35139 5963 35145
rect 5905 35136 5917 35139
rect 5592 35108 5917 35136
rect 5592 35096 5598 35108
rect 5905 35105 5917 35108
rect 5951 35105 5963 35139
rect 5905 35099 5963 35105
rect 5994 35096 6000 35148
rect 6052 35096 6058 35148
rect 6454 35096 6460 35148
rect 6512 35096 6518 35148
rect 6546 35096 6552 35148
rect 6604 35136 6610 35148
rect 8297 35139 8355 35145
rect 6604 35108 6776 35136
rect 6604 35096 6610 35108
rect 6365 35071 6423 35077
rect 6365 35037 6377 35071
rect 6411 35068 6423 35071
rect 6638 35068 6644 35080
rect 6411 35040 6644 35068
rect 6411 35037 6423 35040
rect 6365 35031 6423 35037
rect 6638 35028 6644 35040
rect 6696 35028 6702 35080
rect 6748 35068 6776 35108
rect 8297 35105 8309 35139
rect 8343 35136 8355 35139
rect 8386 35136 8392 35148
rect 8343 35108 8392 35136
rect 8343 35105 8355 35108
rect 8297 35099 8355 35105
rect 8386 35096 8392 35108
rect 8444 35096 8450 35148
rect 8754 35096 8760 35148
rect 8812 35136 8818 35148
rect 9324 35145 9352 35176
rect 11238 35164 11244 35216
rect 11296 35204 11302 35216
rect 16776 35204 16804 35244
rect 11296 35176 16804 35204
rect 11296 35164 11302 35176
rect 17034 35164 17040 35216
rect 17092 35164 17098 35216
rect 17221 35207 17279 35213
rect 17221 35173 17233 35207
rect 17267 35204 17279 35207
rect 17402 35204 17408 35216
rect 17267 35176 17408 35204
rect 17267 35173 17279 35176
rect 17221 35167 17279 35173
rect 17402 35164 17408 35176
rect 17460 35204 17466 35216
rect 17460 35176 18368 35204
rect 17460 35164 17466 35176
rect 9217 35139 9275 35145
rect 9217 35136 9229 35139
rect 8812 35108 9229 35136
rect 8812 35096 8818 35108
rect 9217 35105 9229 35108
rect 9263 35105 9275 35139
rect 9217 35099 9275 35105
rect 9309 35139 9367 35145
rect 9309 35105 9321 35139
rect 9355 35105 9367 35139
rect 9309 35099 9367 35105
rect 12529 35139 12587 35145
rect 12529 35105 12541 35139
rect 12575 35136 12587 35139
rect 13078 35136 13084 35148
rect 12575 35108 13084 35136
rect 12575 35105 12587 35108
rect 12529 35099 12587 35105
rect 13078 35096 13084 35108
rect 13136 35096 13142 35148
rect 13446 35096 13452 35148
rect 13504 35136 13510 35148
rect 16298 35136 16304 35148
rect 13504 35108 16304 35136
rect 13504 35096 13510 35108
rect 16298 35096 16304 35108
rect 16356 35096 16362 35148
rect 17052 35136 17080 35164
rect 17494 35136 17500 35148
rect 17052 35108 17500 35136
rect 17494 35096 17500 35108
rect 17552 35096 17558 35148
rect 17589 35139 17647 35145
rect 17589 35105 17601 35139
rect 17635 35136 17647 35139
rect 17635 35108 18000 35136
rect 17635 35105 17647 35108
rect 17589 35099 17647 35105
rect 17972 35080 18000 35108
rect 6917 35071 6975 35077
rect 6917 35068 6929 35071
rect 6748 35040 6929 35068
rect 6917 35037 6929 35040
rect 6963 35037 6975 35071
rect 6917 35031 6975 35037
rect 1302 34960 1308 35012
rect 1360 35000 1366 35012
rect 1397 35003 1455 35009
rect 1397 35000 1409 35003
rect 1360 34972 1409 35000
rect 1360 34960 1366 34972
rect 1397 34969 1409 34972
rect 1443 34969 1455 35003
rect 1397 34963 1455 34969
rect 2682 34960 2688 35012
rect 2740 34960 2746 35012
rect 5629 35003 5687 35009
rect 5198 34972 5304 35000
rect 5276 34932 5304 34972
rect 5629 34969 5641 35003
rect 5675 35000 5687 35003
rect 6733 35003 6791 35009
rect 6733 35000 6745 35003
rect 5675 34972 6745 35000
rect 5675 34969 5687 34972
rect 5629 34963 5687 34969
rect 6733 34969 6745 34972
rect 6779 34969 6791 35003
rect 6733 34963 6791 34969
rect 5902 34932 5908 34944
rect 5276 34904 5908 34932
rect 5902 34892 5908 34904
rect 5960 34892 5966 34944
rect 6546 34892 6552 34944
rect 6604 34932 6610 34944
rect 6641 34935 6699 34941
rect 6641 34932 6653 34935
rect 6604 34904 6653 34932
rect 6604 34892 6610 34904
rect 6641 34901 6653 34904
rect 6687 34901 6699 34935
rect 6932 34932 6960 35031
rect 7098 35028 7104 35080
rect 7156 35028 7162 35080
rect 7190 35028 7196 35080
rect 7248 35028 7254 35080
rect 7374 35028 7380 35080
rect 7432 35028 7438 35080
rect 7466 35028 7472 35080
rect 7524 35068 7530 35080
rect 7561 35071 7619 35077
rect 7561 35068 7573 35071
rect 7524 35040 7573 35068
rect 7524 35028 7530 35040
rect 7561 35037 7573 35040
rect 7607 35037 7619 35071
rect 7561 35031 7619 35037
rect 7576 35000 7604 35031
rect 8018 35028 8024 35080
rect 8076 35028 8082 35080
rect 8202 35028 8208 35080
rect 8260 35028 8266 35080
rect 8481 35071 8539 35077
rect 8481 35037 8493 35071
rect 8527 35037 8539 35071
rect 8481 35031 8539 35037
rect 8665 35071 8723 35077
rect 8665 35037 8677 35071
rect 8711 35068 8723 35071
rect 9030 35068 9036 35080
rect 8711 35040 9036 35068
rect 8711 35037 8723 35040
rect 8665 35031 8723 35037
rect 8110 35000 8116 35012
rect 7576 34972 8116 35000
rect 8110 34960 8116 34972
rect 8168 34960 8174 35012
rect 8496 35000 8524 35031
rect 9030 35028 9036 35040
rect 9088 35028 9094 35080
rect 9122 35028 9128 35080
rect 9180 35028 9186 35080
rect 9398 35028 9404 35080
rect 9456 35028 9462 35080
rect 12250 35028 12256 35080
rect 12308 35028 12314 35080
rect 12434 35028 12440 35080
rect 12492 35028 12498 35080
rect 12894 35028 12900 35080
rect 12952 35028 12958 35080
rect 16485 35071 16543 35077
rect 16485 35037 16497 35071
rect 16531 35068 16543 35071
rect 16850 35068 16856 35080
rect 16531 35040 16856 35068
rect 16531 35037 16543 35040
rect 16485 35031 16543 35037
rect 16850 35028 16856 35040
rect 16908 35028 16914 35080
rect 17678 35028 17684 35080
rect 17736 35068 17742 35080
rect 17865 35071 17923 35077
rect 17865 35068 17877 35071
rect 17736 35040 17877 35068
rect 17736 35028 17742 35040
rect 17865 35037 17877 35040
rect 17911 35037 17923 35071
rect 17865 35031 17923 35037
rect 17954 35028 17960 35080
rect 18012 35068 18018 35080
rect 18340 35077 18368 35176
rect 18432 35136 18460 35244
rect 19242 35232 19248 35284
rect 19300 35272 19306 35284
rect 20806 35272 20812 35284
rect 19300 35244 20812 35272
rect 19300 35232 19306 35244
rect 20806 35232 20812 35244
rect 20864 35232 20870 35284
rect 22278 35272 22284 35284
rect 21008 35244 22284 35272
rect 18506 35164 18512 35216
rect 18564 35204 18570 35216
rect 18874 35204 18880 35216
rect 18564 35176 18880 35204
rect 18564 35164 18570 35176
rect 18874 35164 18880 35176
rect 18932 35204 18938 35216
rect 19337 35207 19395 35213
rect 19337 35204 19349 35207
rect 18932 35176 19349 35204
rect 18932 35164 18938 35176
rect 19337 35173 19349 35176
rect 19383 35173 19395 35207
rect 19702 35204 19708 35216
rect 19337 35167 19395 35173
rect 19536 35176 19708 35204
rect 18432 35108 19334 35136
rect 18049 35071 18107 35077
rect 18049 35068 18061 35071
rect 18012 35040 18061 35068
rect 18012 35028 18018 35040
rect 18049 35037 18061 35040
rect 18095 35037 18107 35071
rect 18049 35031 18107 35037
rect 18325 35071 18383 35077
rect 18325 35037 18337 35071
rect 18371 35037 18383 35071
rect 19306 35068 19334 35108
rect 19536 35077 19564 35176
rect 19702 35164 19708 35176
rect 19760 35164 19766 35216
rect 21008 35136 21036 35244
rect 22278 35232 22284 35244
rect 22336 35232 22342 35284
rect 21634 35164 21640 35216
rect 21692 35204 21698 35216
rect 21692 35176 21956 35204
rect 21692 35164 21698 35176
rect 20916 35108 21036 35136
rect 19521 35071 19579 35077
rect 19521 35068 19533 35071
rect 19306 35040 19533 35068
rect 18325 35031 18383 35037
rect 19521 35037 19533 35040
rect 19567 35037 19579 35071
rect 19521 35031 19579 35037
rect 19886 35028 19892 35080
rect 19944 35028 19950 35080
rect 20530 35028 20536 35080
rect 20588 35068 20594 35080
rect 20916 35077 20944 35108
rect 21266 35096 21272 35148
rect 21324 35096 21330 35148
rect 21545 35139 21603 35145
rect 21545 35105 21557 35139
rect 21591 35136 21603 35139
rect 21726 35136 21732 35148
rect 21591 35108 21732 35136
rect 21591 35105 21603 35108
rect 21545 35099 21603 35105
rect 21726 35096 21732 35108
rect 21784 35096 21790 35148
rect 20717 35071 20775 35077
rect 20717 35068 20729 35071
rect 20588 35040 20729 35068
rect 20588 35028 20594 35040
rect 20717 35037 20729 35040
rect 20763 35037 20775 35071
rect 20717 35031 20775 35037
rect 20901 35071 20959 35077
rect 20901 35037 20913 35071
rect 20947 35037 20959 35071
rect 20901 35031 20959 35037
rect 20990 35028 20996 35080
rect 21048 35068 21054 35080
rect 21177 35071 21235 35077
rect 21177 35068 21189 35071
rect 21048 35040 21189 35068
rect 21048 35028 21054 35040
rect 21177 35037 21189 35040
rect 21223 35037 21235 35071
rect 21284 35068 21312 35096
rect 21928 35077 21956 35176
rect 21913 35071 21971 35077
rect 21284 35040 21772 35068
rect 21177 35031 21235 35037
rect 9140 35000 9168 35028
rect 8496 34972 9168 35000
rect 11882 34960 11888 35012
rect 11940 35000 11946 35012
rect 15654 35000 15660 35012
rect 11940 34972 15660 35000
rect 11940 34960 11946 34972
rect 15654 34960 15660 34972
rect 15712 34960 15718 35012
rect 15838 34960 15844 35012
rect 15896 35000 15902 35012
rect 16209 35003 16267 35009
rect 16209 35000 16221 35003
rect 15896 34972 16221 35000
rect 15896 34960 15902 34972
rect 16209 34969 16221 34972
rect 16255 35000 16267 35003
rect 16390 35000 16396 35012
rect 16255 34972 16396 35000
rect 16255 34969 16267 34972
rect 16209 34963 16267 34969
rect 16390 34960 16396 34972
rect 16448 34960 16454 35012
rect 16666 34960 16672 35012
rect 16724 35000 16730 35012
rect 16761 35003 16819 35009
rect 16761 35000 16773 35003
rect 16724 34972 16773 35000
rect 16724 34960 16730 34972
rect 16761 34969 16773 34972
rect 16807 34969 16819 35003
rect 16761 34963 16819 34969
rect 10778 34932 10784 34944
rect 6932 34904 10784 34932
rect 6641 34895 6699 34901
rect 10778 34892 10784 34904
rect 10836 34892 10842 34944
rect 11330 34892 11336 34944
rect 11388 34932 11394 34944
rect 12069 34935 12127 34941
rect 12069 34932 12081 34935
rect 11388 34904 12081 34932
rect 11388 34892 11394 34904
rect 12069 34901 12081 34904
rect 12115 34901 12127 34935
rect 12069 34895 12127 34901
rect 12342 34892 12348 34944
rect 12400 34932 12406 34944
rect 12713 34935 12771 34941
rect 12713 34932 12725 34935
rect 12400 34904 12725 34932
rect 12400 34892 12406 34904
rect 12713 34901 12725 34904
rect 12759 34901 12771 34935
rect 16868 34932 16896 35028
rect 17310 34960 17316 35012
rect 17368 34960 17374 35012
rect 17770 34960 17776 35012
rect 17828 34960 17834 35012
rect 18690 34960 18696 35012
rect 18748 35000 18754 35012
rect 21744 35000 21772 35040
rect 21913 35037 21925 35071
rect 21959 35037 21971 35071
rect 21913 35031 21971 35037
rect 22462 35028 22468 35080
rect 22520 35028 22526 35080
rect 22554 35000 22560 35012
rect 18748 34972 21680 35000
rect 21744 34972 22560 35000
rect 18748 34960 18754 34972
rect 21192 34944 21220 34972
rect 17405 34935 17463 34941
rect 17405 34932 17417 34935
rect 16868 34904 17417 34932
rect 12713 34895 12771 34901
rect 17405 34901 17417 34904
rect 17451 34932 17463 34935
rect 17494 34932 17500 34944
rect 17451 34904 17500 34932
rect 17451 34901 17463 34904
rect 17405 34895 17463 34901
rect 17494 34892 17500 34904
rect 17552 34892 17558 34944
rect 18506 34892 18512 34944
rect 18564 34892 18570 34944
rect 18782 34892 18788 34944
rect 18840 34932 18846 34944
rect 19702 34932 19708 34944
rect 18840 34904 19708 34932
rect 18840 34892 18846 34904
rect 19702 34892 19708 34904
rect 19760 34892 19766 34944
rect 20898 34892 20904 34944
rect 20956 34892 20962 34944
rect 21174 34892 21180 34944
rect 21232 34892 21238 34944
rect 21652 34932 21680 34972
rect 22554 34960 22560 34972
rect 22612 35000 22618 35012
rect 22649 35003 22707 35009
rect 22649 35000 22661 35003
rect 22612 34972 22661 35000
rect 22612 34960 22618 34972
rect 22649 34969 22661 34972
rect 22695 34969 22707 35003
rect 22649 34963 22707 34969
rect 22922 34960 22928 35012
rect 22980 34960 22986 35012
rect 22830 34932 22836 34944
rect 21652 34904 22836 34932
rect 22830 34892 22836 34904
rect 22888 34892 22894 34944
rect 1104 34842 40572 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 40572 34842
rect 1104 34768 40572 34790
rect 2682 34688 2688 34740
rect 2740 34728 2746 34740
rect 7009 34731 7067 34737
rect 2740 34700 3740 34728
rect 2740 34688 2746 34700
rect 3712 34660 3740 34700
rect 7009 34697 7021 34731
rect 7055 34728 7067 34731
rect 7098 34728 7104 34740
rect 7055 34700 7104 34728
rect 7055 34697 7067 34700
rect 7009 34691 7067 34697
rect 7098 34688 7104 34700
rect 7156 34688 7162 34740
rect 8757 34731 8815 34737
rect 8757 34697 8769 34731
rect 8803 34728 8815 34731
rect 9398 34728 9404 34740
rect 8803 34700 9404 34728
rect 8803 34697 8815 34700
rect 8757 34691 8815 34697
rect 9398 34688 9404 34700
rect 9456 34688 9462 34740
rect 13814 34728 13820 34740
rect 11992 34700 13820 34728
rect 5902 34660 5908 34672
rect 3634 34632 5908 34660
rect 5902 34620 5908 34632
rect 5960 34620 5966 34672
rect 6178 34620 6184 34672
rect 6236 34660 6242 34672
rect 8202 34660 8208 34672
rect 6236 34632 8208 34660
rect 6236 34620 6242 34632
rect 4341 34595 4399 34601
rect 4341 34561 4353 34595
rect 4387 34592 4399 34595
rect 5534 34592 5540 34604
rect 4387 34564 5540 34592
rect 4387 34561 4399 34564
rect 4341 34555 4399 34561
rect 5534 34552 5540 34564
rect 5592 34552 5598 34604
rect 6086 34552 6092 34604
rect 6144 34592 6150 34604
rect 6365 34595 6423 34601
rect 6365 34592 6377 34595
rect 6144 34564 6377 34592
rect 6144 34552 6150 34564
rect 6365 34561 6377 34564
rect 6411 34561 6423 34595
rect 6365 34555 6423 34561
rect 6546 34552 6552 34604
rect 6604 34552 6610 34604
rect 6638 34552 6644 34604
rect 6696 34552 6702 34604
rect 6748 34601 6776 34632
rect 8202 34620 8208 34632
rect 8260 34620 8266 34672
rect 8478 34620 8484 34672
rect 8536 34660 8542 34672
rect 10965 34663 11023 34669
rect 8536 34632 8892 34660
rect 8536 34620 8542 34632
rect 6733 34595 6791 34601
rect 6733 34561 6745 34595
rect 6779 34561 6791 34595
rect 8570 34592 8576 34604
rect 6733 34555 6791 34561
rect 7576 34564 8576 34592
rect 2314 34484 2320 34536
rect 2372 34484 2378 34536
rect 4062 34484 4068 34536
rect 4120 34484 4126 34536
rect 5552 34524 5580 34552
rect 6822 34524 6828 34536
rect 5552 34496 6828 34524
rect 6822 34484 6828 34496
rect 6880 34484 6886 34536
rect 6086 34416 6092 34468
rect 6144 34456 6150 34468
rect 7098 34456 7104 34468
rect 6144 34428 7104 34456
rect 6144 34416 6150 34428
rect 7098 34416 7104 34428
rect 7156 34456 7162 34468
rect 7576 34456 7604 34564
rect 8570 34552 8576 34564
rect 8628 34592 8634 34604
rect 8864 34601 8892 34632
rect 10965 34629 10977 34663
rect 11011 34660 11023 34663
rect 11422 34660 11428 34672
rect 11011 34632 11428 34660
rect 11011 34629 11023 34632
rect 10965 34623 11023 34629
rect 11422 34620 11428 34632
rect 11480 34620 11486 34672
rect 8665 34595 8723 34601
rect 8665 34592 8677 34595
rect 8628 34564 8677 34592
rect 8628 34552 8634 34564
rect 8665 34561 8677 34564
rect 8711 34561 8723 34595
rect 8665 34555 8723 34561
rect 8849 34595 8907 34601
rect 8849 34561 8861 34595
rect 8895 34561 8907 34595
rect 8849 34555 8907 34561
rect 8938 34552 8944 34604
rect 8996 34592 9002 34604
rect 9217 34595 9275 34601
rect 9217 34592 9229 34595
rect 8996 34564 9229 34592
rect 8996 34552 9002 34564
rect 9217 34561 9229 34564
rect 9263 34561 9275 34595
rect 9217 34555 9275 34561
rect 9401 34595 9459 34601
rect 9401 34561 9413 34595
rect 9447 34561 9459 34595
rect 9401 34555 9459 34561
rect 8478 34484 8484 34536
rect 8536 34524 8542 34536
rect 9416 34524 9444 34555
rect 9582 34552 9588 34604
rect 9640 34592 9646 34604
rect 9953 34595 10011 34601
rect 9953 34592 9965 34595
rect 9640 34564 9965 34592
rect 9640 34552 9646 34564
rect 9953 34561 9965 34564
rect 9999 34561 10011 34595
rect 9953 34555 10011 34561
rect 10134 34552 10140 34604
rect 10192 34552 10198 34604
rect 10594 34552 10600 34604
rect 10652 34552 10658 34604
rect 10778 34552 10784 34604
rect 10836 34601 10842 34604
rect 10836 34595 10885 34601
rect 10836 34561 10839 34595
rect 10873 34561 10885 34595
rect 10836 34555 10885 34561
rect 10836 34552 10842 34555
rect 11054 34552 11060 34604
rect 11112 34552 11118 34604
rect 11238 34592 11244 34604
rect 11199 34564 11244 34592
rect 11238 34552 11244 34564
rect 11296 34552 11302 34604
rect 11330 34552 11336 34604
rect 11388 34552 11394 34604
rect 11882 34552 11888 34604
rect 11940 34552 11946 34604
rect 8536 34496 9444 34524
rect 8536 34484 8542 34496
rect 10318 34484 10324 34536
rect 10376 34484 10382 34536
rect 10686 34484 10692 34536
rect 10744 34524 10750 34536
rect 11992 34533 12020 34700
rect 13814 34688 13820 34700
rect 13872 34688 13878 34740
rect 17402 34688 17408 34740
rect 17460 34688 17466 34740
rect 17494 34688 17500 34740
rect 17552 34728 17558 34740
rect 18325 34731 18383 34737
rect 17552 34700 18276 34728
rect 17552 34688 17558 34700
rect 15010 34660 15016 34672
rect 13478 34632 15016 34660
rect 15010 34620 15016 34632
rect 15068 34620 15074 34672
rect 17589 34663 17647 34669
rect 17589 34629 17601 34663
rect 17635 34660 17647 34663
rect 17770 34660 17776 34672
rect 17635 34632 17776 34660
rect 17635 34629 17647 34632
rect 17589 34623 17647 34629
rect 17770 34620 17776 34632
rect 17828 34620 17834 34672
rect 18248 34660 18276 34700
rect 18325 34697 18337 34731
rect 18371 34728 18383 34731
rect 18506 34728 18512 34740
rect 18371 34700 18512 34728
rect 18371 34697 18383 34700
rect 18325 34691 18383 34697
rect 18506 34688 18512 34700
rect 18564 34688 18570 34740
rect 18782 34688 18788 34740
rect 18840 34688 18846 34740
rect 21542 34728 21548 34740
rect 18984 34700 21548 34728
rect 18800 34660 18828 34688
rect 18248 34632 18828 34660
rect 14369 34595 14427 34601
rect 14369 34561 14381 34595
rect 14415 34592 14427 34595
rect 15286 34592 15292 34604
rect 14415 34564 15292 34592
rect 14415 34561 14427 34564
rect 14369 34555 14427 34561
rect 15286 34552 15292 34564
rect 15344 34552 15350 34604
rect 16022 34552 16028 34604
rect 16080 34592 16086 34604
rect 17310 34592 17316 34604
rect 16080 34564 17316 34592
rect 16080 34552 16086 34564
rect 17310 34552 17316 34564
rect 17368 34592 17374 34604
rect 18230 34592 18236 34604
rect 17368 34564 18236 34592
rect 17368 34552 17374 34564
rect 18230 34552 18236 34564
rect 18288 34552 18294 34604
rect 18509 34595 18567 34601
rect 18509 34561 18521 34595
rect 18555 34592 18567 34595
rect 18598 34592 18604 34604
rect 18555 34564 18604 34592
rect 18555 34561 18567 34564
rect 18509 34555 18567 34561
rect 18598 34552 18604 34564
rect 18656 34552 18662 34604
rect 18984 34601 19012 34700
rect 21542 34688 21548 34700
rect 21600 34688 21606 34740
rect 23750 34688 23756 34740
rect 23808 34728 23814 34740
rect 31110 34728 31116 34740
rect 23808 34700 31116 34728
rect 23808 34688 23814 34700
rect 31110 34688 31116 34700
rect 31168 34688 31174 34740
rect 19058 34620 19064 34672
rect 19116 34660 19122 34672
rect 19521 34663 19579 34669
rect 19116 34632 19196 34660
rect 19116 34620 19122 34632
rect 19168 34601 19196 34632
rect 19521 34629 19533 34663
rect 19567 34660 19579 34663
rect 19889 34663 19947 34669
rect 19889 34660 19901 34663
rect 19567 34632 19901 34660
rect 19567 34629 19579 34632
rect 19521 34623 19579 34629
rect 19889 34629 19901 34632
rect 19935 34629 19947 34663
rect 19889 34623 19947 34629
rect 21174 34620 21180 34672
rect 21232 34660 21238 34672
rect 21634 34660 21640 34672
rect 21232 34632 21640 34660
rect 21232 34620 21238 34632
rect 21634 34620 21640 34632
rect 21692 34660 21698 34672
rect 25593 34663 25651 34669
rect 21692 34632 23612 34660
rect 21692 34620 21698 34632
rect 18693 34595 18751 34601
rect 18693 34561 18705 34595
rect 18739 34592 18751 34595
rect 18785 34595 18843 34601
rect 18785 34592 18797 34595
rect 18739 34564 18797 34592
rect 18739 34561 18751 34564
rect 18693 34555 18751 34561
rect 18785 34561 18797 34564
rect 18831 34561 18843 34595
rect 18785 34555 18843 34561
rect 18969 34595 19027 34601
rect 18969 34561 18981 34595
rect 19015 34561 19027 34595
rect 18969 34555 19027 34561
rect 19153 34595 19211 34601
rect 19153 34561 19165 34595
rect 19199 34561 19211 34595
rect 19153 34555 19211 34561
rect 19242 34552 19248 34604
rect 19300 34592 19306 34604
rect 19337 34595 19395 34601
rect 19337 34592 19349 34595
rect 19300 34564 19349 34592
rect 19300 34552 19306 34564
rect 19337 34561 19349 34564
rect 19383 34561 19395 34595
rect 19337 34555 19395 34561
rect 11977 34527 12035 34533
rect 11977 34524 11989 34527
rect 10744 34496 11989 34524
rect 10744 34484 10750 34496
rect 11977 34493 11989 34496
rect 12023 34493 12035 34527
rect 12253 34527 12311 34533
rect 12253 34524 12265 34527
rect 11977 34487 12035 34493
rect 12084 34496 12265 34524
rect 7156 34428 7604 34456
rect 7156 34416 7162 34428
rect 8386 34416 8392 34468
rect 8444 34456 8450 34468
rect 9766 34456 9772 34468
rect 8444 34428 9772 34456
rect 8444 34416 8450 34428
rect 9766 34416 9772 34428
rect 9824 34416 9830 34468
rect 10505 34459 10563 34465
rect 10505 34425 10517 34459
rect 10551 34456 10563 34459
rect 10962 34456 10968 34468
rect 10551 34428 10968 34456
rect 10551 34425 10563 34428
rect 10505 34419 10563 34425
rect 10962 34416 10968 34428
rect 11020 34416 11026 34468
rect 12084 34456 12112 34496
rect 12253 34493 12265 34496
rect 12299 34493 12311 34527
rect 13725 34527 13783 34533
rect 13725 34524 13737 34527
rect 12253 34487 12311 34493
rect 13280 34496 13737 34524
rect 11532 34428 12112 34456
rect 9122 34348 9128 34400
rect 9180 34388 9186 34400
rect 9217 34391 9275 34397
rect 9217 34388 9229 34391
rect 9180 34360 9229 34388
rect 9180 34348 9186 34360
rect 9217 34357 9229 34360
rect 9263 34357 9275 34391
rect 9217 34351 9275 34357
rect 10134 34348 10140 34400
rect 10192 34348 10198 34400
rect 10226 34348 10232 34400
rect 10284 34388 10290 34400
rect 10413 34391 10471 34397
rect 10413 34388 10425 34391
rect 10284 34360 10425 34388
rect 10284 34348 10290 34360
rect 10413 34357 10425 34360
rect 10459 34357 10471 34391
rect 10413 34351 10471 34357
rect 10689 34391 10747 34397
rect 10689 34357 10701 34391
rect 10735 34388 10747 34391
rect 11532 34388 11560 34428
rect 10735 34360 11560 34388
rect 10735 34357 10747 34360
rect 10689 34351 10747 34357
rect 11698 34348 11704 34400
rect 11756 34348 11762 34400
rect 12066 34348 12072 34400
rect 12124 34388 12130 34400
rect 13280 34388 13308 34496
rect 13725 34493 13737 34496
rect 13771 34493 13783 34527
rect 13725 34487 13783 34493
rect 14274 34484 14280 34536
rect 14332 34484 14338 34536
rect 15654 34484 15660 34536
rect 15712 34524 15718 34536
rect 19061 34527 19119 34533
rect 19061 34524 19073 34527
rect 15712 34496 19073 34524
rect 15712 34484 15718 34496
rect 19061 34493 19073 34496
rect 19107 34493 19119 34527
rect 19610 34524 19616 34536
rect 19061 34487 19119 34493
rect 19168 34496 19616 34524
rect 17678 34416 17684 34468
rect 17736 34456 17742 34468
rect 19168 34456 19196 34496
rect 19610 34484 19616 34496
rect 19668 34484 19674 34536
rect 21008 34524 21036 34578
rect 21450 34552 21456 34604
rect 21508 34592 21514 34604
rect 22005 34595 22063 34601
rect 22005 34592 22017 34595
rect 21508 34564 22017 34592
rect 21508 34552 21514 34564
rect 22005 34561 22017 34564
rect 22051 34561 22063 34595
rect 22005 34555 22063 34561
rect 22097 34595 22155 34601
rect 22097 34561 22109 34595
rect 22143 34561 22155 34595
rect 22097 34555 22155 34561
rect 19720 34496 21036 34524
rect 17736 34428 19196 34456
rect 17736 34416 17742 34428
rect 19242 34416 19248 34468
rect 19300 34456 19306 34468
rect 19720 34456 19748 34496
rect 21082 34484 21088 34536
rect 21140 34524 21146 34536
rect 21637 34527 21695 34533
rect 21637 34524 21649 34527
rect 21140 34496 21649 34524
rect 21140 34484 21146 34496
rect 21637 34493 21649 34496
rect 21683 34524 21695 34527
rect 21683 34496 21772 34524
rect 21683 34493 21695 34496
rect 21637 34487 21695 34493
rect 19300 34428 19748 34456
rect 21744 34456 21772 34496
rect 21818 34484 21824 34536
rect 21876 34524 21882 34536
rect 22112 34524 22140 34555
rect 22186 34552 22192 34604
rect 22244 34552 22250 34604
rect 22327 34595 22385 34601
rect 22327 34561 22339 34595
rect 22373 34592 22385 34595
rect 22554 34592 22560 34604
rect 22373 34564 22560 34592
rect 22373 34561 22385 34564
rect 22327 34555 22385 34561
rect 22554 34552 22560 34564
rect 22612 34552 22618 34604
rect 22830 34552 22836 34604
rect 22888 34592 22894 34604
rect 23584 34601 23612 34632
rect 25593 34629 25605 34663
rect 25639 34660 25651 34663
rect 25682 34660 25688 34672
rect 25639 34632 25688 34660
rect 25639 34629 25651 34632
rect 25593 34623 25651 34629
rect 25682 34620 25688 34632
rect 25740 34620 25746 34672
rect 22925 34595 22983 34601
rect 22925 34592 22937 34595
rect 22888 34564 22937 34592
rect 22888 34552 22894 34564
rect 22925 34561 22937 34564
rect 22971 34561 22983 34595
rect 22925 34555 22983 34561
rect 23569 34595 23627 34601
rect 23569 34561 23581 34595
rect 23615 34561 23627 34595
rect 23569 34555 23627 34561
rect 24946 34552 24952 34604
rect 25004 34592 25010 34604
rect 28258 34592 28264 34604
rect 25004 34564 28264 34592
rect 25004 34552 25010 34564
rect 28258 34552 28264 34564
rect 28316 34552 28322 34604
rect 28902 34552 28908 34604
rect 28960 34592 28966 34604
rect 30377 34595 30435 34601
rect 30377 34592 30389 34595
rect 28960 34564 30389 34592
rect 28960 34552 28966 34564
rect 30377 34561 30389 34564
rect 30423 34561 30435 34595
rect 30377 34555 30435 34561
rect 22465 34527 22523 34533
rect 22465 34524 22477 34527
rect 21876 34496 22140 34524
rect 22204 34496 22477 34524
rect 21876 34484 21882 34496
rect 22204 34456 22232 34496
rect 22465 34493 22477 34496
rect 22511 34493 22523 34527
rect 22465 34487 22523 34493
rect 23842 34484 23848 34536
rect 23900 34484 23906 34536
rect 28350 34484 28356 34536
rect 28408 34484 28414 34536
rect 21744 34428 22232 34456
rect 19300 34416 19306 34428
rect 12124 34360 13308 34388
rect 14645 34391 14703 34397
rect 12124 34348 12130 34360
rect 14645 34357 14657 34391
rect 14691 34388 14703 34391
rect 14734 34388 14740 34400
rect 14691 34360 14740 34388
rect 14691 34357 14703 34360
rect 14645 34351 14703 34357
rect 14734 34348 14740 34360
rect 14792 34348 14798 34400
rect 17402 34348 17408 34400
rect 17460 34388 17466 34400
rect 17589 34391 17647 34397
rect 17589 34388 17601 34391
rect 17460 34360 17601 34388
rect 17460 34348 17466 34360
rect 17589 34357 17601 34360
rect 17635 34357 17647 34391
rect 17589 34351 17647 34357
rect 18138 34348 18144 34400
rect 18196 34388 18202 34400
rect 19058 34388 19064 34400
rect 18196 34360 19064 34388
rect 18196 34348 18202 34360
rect 19058 34348 19064 34360
rect 19116 34348 19122 34400
rect 21818 34348 21824 34400
rect 21876 34348 21882 34400
rect 28994 34348 29000 34400
rect 29052 34348 29058 34400
rect 1104 34298 40572 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 40572 34298
rect 1104 34224 40572 34246
rect 3053 34187 3111 34193
rect 3053 34153 3065 34187
rect 3099 34184 3111 34187
rect 4062 34184 4068 34196
rect 3099 34156 4068 34184
rect 3099 34153 3111 34156
rect 3053 34147 3111 34153
rect 4062 34144 4068 34156
rect 4120 34144 4126 34196
rect 6546 34144 6552 34196
rect 6604 34184 6610 34196
rect 7282 34184 7288 34196
rect 6604 34156 7288 34184
rect 6604 34144 6610 34156
rect 7282 34144 7288 34156
rect 7340 34144 7346 34196
rect 8754 34144 8760 34196
rect 8812 34144 8818 34196
rect 9030 34144 9036 34196
rect 9088 34184 9094 34196
rect 9217 34187 9275 34193
rect 9217 34184 9229 34187
rect 9088 34156 9229 34184
rect 9088 34144 9094 34156
rect 9217 34153 9229 34156
rect 9263 34153 9275 34187
rect 9217 34147 9275 34153
rect 9674 34144 9680 34196
rect 9732 34184 9738 34196
rect 9953 34187 10011 34193
rect 9953 34184 9965 34187
rect 9732 34156 9965 34184
rect 9732 34144 9738 34156
rect 9953 34153 9965 34156
rect 9999 34153 10011 34187
rect 9953 34147 10011 34153
rect 10594 34144 10600 34196
rect 10652 34184 10658 34196
rect 10781 34187 10839 34193
rect 10781 34184 10793 34187
rect 10652 34156 10793 34184
rect 10652 34144 10658 34156
rect 10781 34153 10793 34156
rect 10827 34153 10839 34187
rect 10781 34147 10839 34153
rect 8938 34116 8944 34128
rect 8588 34088 8944 34116
rect 6730 34048 6736 34060
rect 3252 34020 6736 34048
rect 3252 33989 3280 34020
rect 6730 34008 6736 34020
rect 6788 34008 6794 34060
rect 8202 34008 8208 34060
rect 8260 34048 8266 34060
rect 8588 34048 8616 34088
rect 8938 34076 8944 34088
rect 8996 34076 9002 34128
rect 9585 34119 9643 34125
rect 9585 34085 9597 34119
rect 9631 34116 9643 34119
rect 9631 34088 10180 34116
rect 9631 34085 9643 34088
rect 9585 34079 9643 34085
rect 8260 34020 8616 34048
rect 8260 34008 8266 34020
rect 3237 33983 3295 33989
rect 3237 33949 3249 33983
rect 3283 33949 3295 33983
rect 3237 33943 3295 33949
rect 3513 33983 3571 33989
rect 3513 33949 3525 33983
rect 3559 33980 3571 33983
rect 4154 33980 4160 33992
rect 3559 33952 4160 33980
rect 3559 33949 3571 33952
rect 3513 33943 3571 33949
rect 4154 33940 4160 33952
rect 4212 33980 4218 33992
rect 4614 33980 4620 33992
rect 4212 33952 4620 33980
rect 4212 33940 4218 33952
rect 4614 33940 4620 33952
rect 4672 33940 4678 33992
rect 5626 33940 5632 33992
rect 5684 33980 5690 33992
rect 8478 33980 8484 33992
rect 5684 33952 8484 33980
rect 5684 33940 5690 33952
rect 8478 33940 8484 33952
rect 8536 33940 8542 33992
rect 8588 33989 8616 34020
rect 9033 34051 9091 34057
rect 9033 34017 9045 34051
rect 9079 34048 9091 34051
rect 10045 34051 10103 34057
rect 10045 34048 10057 34051
rect 9079 34020 10057 34048
rect 9079 34017 9091 34020
rect 9033 34011 9091 34017
rect 8573 33983 8631 33989
rect 8573 33949 8585 33983
rect 8619 33949 8631 33983
rect 8573 33943 8631 33949
rect 8754 33940 8760 33992
rect 8812 33980 8818 33992
rect 8941 33983 8999 33989
rect 8941 33980 8953 33983
rect 8812 33952 8953 33980
rect 8812 33940 8818 33952
rect 8941 33949 8953 33952
rect 8987 33949 8999 33983
rect 8941 33943 8999 33949
rect 9122 33940 9128 33992
rect 9180 33940 9186 33992
rect 9416 33989 9444 34020
rect 10045 34017 10057 34020
rect 10091 34017 10103 34051
rect 10045 34011 10103 34017
rect 10152 34048 10180 34088
rect 10413 34051 10471 34057
rect 10413 34048 10425 34051
rect 10152 34020 10425 34048
rect 9401 33983 9459 33989
rect 9401 33949 9413 33983
rect 9447 33949 9459 33983
rect 9401 33943 9459 33949
rect 9674 33940 9680 33992
rect 9732 33940 9738 33992
rect 10152 33989 10180 34020
rect 10413 34017 10425 34020
rect 10459 34017 10471 34051
rect 10413 34011 10471 34017
rect 10137 33983 10195 33989
rect 10137 33949 10149 33983
rect 10183 33949 10195 33983
rect 10137 33943 10195 33949
rect 1670 33872 1676 33924
rect 1728 33912 1734 33924
rect 2314 33912 2320 33924
rect 1728 33884 2320 33912
rect 1728 33872 1734 33884
rect 2314 33872 2320 33884
rect 2372 33912 2378 33924
rect 3421 33915 3479 33921
rect 3421 33912 3433 33915
rect 2372 33884 3433 33912
rect 2372 33872 2378 33884
rect 3421 33881 3433 33884
rect 3467 33881 3479 33915
rect 3421 33875 3479 33881
rect 8662 33872 8668 33924
rect 8720 33912 8726 33924
rect 8720 33884 9996 33912
rect 8720 33872 8726 33884
rect 9766 33804 9772 33856
rect 9824 33804 9830 33856
rect 9968 33844 9996 33884
rect 10042 33872 10048 33924
rect 10100 33912 10106 33924
rect 10152 33912 10180 33943
rect 10318 33940 10324 33992
rect 10376 33980 10382 33992
rect 10597 33983 10655 33989
rect 10597 33980 10609 33983
rect 10376 33952 10609 33980
rect 10376 33940 10382 33952
rect 10597 33949 10609 33952
rect 10643 33949 10655 33983
rect 10597 33943 10655 33949
rect 10100 33884 10180 33912
rect 10796 33912 10824 34147
rect 10962 34144 10968 34196
rect 11020 34144 11026 34196
rect 11977 34187 12035 34193
rect 11977 34153 11989 34187
rect 12023 34184 12035 34187
rect 12250 34184 12256 34196
rect 12023 34156 12256 34184
rect 12023 34153 12035 34156
rect 11977 34147 12035 34153
rect 12250 34144 12256 34156
rect 12308 34144 12314 34196
rect 12434 34144 12440 34196
rect 12492 34184 12498 34196
rect 12621 34187 12679 34193
rect 12621 34184 12633 34187
rect 12492 34156 12633 34184
rect 12492 34144 12498 34156
rect 12621 34153 12633 34156
rect 12667 34153 12679 34187
rect 12621 34147 12679 34153
rect 10873 34051 10931 34057
rect 10873 34017 10885 34051
rect 10919 34048 10931 34051
rect 10980 34048 11008 34144
rect 10919 34020 11008 34048
rect 11164 34088 12388 34116
rect 10919 34017 10931 34020
rect 10873 34011 10931 34017
rect 11164 33992 11192 34088
rect 12360 34060 12388 34088
rect 12066 34048 12072 34060
rect 11348 34020 12072 34048
rect 11348 33992 11376 34020
rect 12066 34008 12072 34020
rect 12124 34048 12130 34060
rect 12124 34020 12296 34048
rect 12124 34008 12130 34020
rect 11146 33940 11152 33992
rect 11204 33940 11210 33992
rect 11330 33940 11336 33992
rect 11388 33940 11394 33992
rect 11698 33940 11704 33992
rect 11756 33980 11762 33992
rect 12268 33989 12296 34020
rect 12342 34008 12348 34060
rect 12400 34008 12406 34060
rect 11793 33983 11851 33989
rect 11793 33980 11805 33983
rect 11756 33952 11805 33980
rect 11756 33940 11762 33952
rect 11793 33949 11805 33952
rect 11839 33949 11851 33983
rect 11793 33943 11851 33949
rect 11977 33983 12035 33989
rect 11977 33949 11989 33983
rect 12023 33949 12035 33983
rect 11977 33943 12035 33949
rect 12253 33983 12311 33989
rect 12253 33949 12265 33983
rect 12299 33949 12311 33983
rect 12636 33980 12664 34147
rect 18322 34144 18328 34196
rect 18380 34184 18386 34196
rect 18417 34187 18475 34193
rect 18417 34184 18429 34187
rect 18380 34156 18429 34184
rect 18380 34144 18386 34156
rect 18417 34153 18429 34156
rect 18463 34153 18475 34187
rect 18417 34147 18475 34153
rect 18598 34144 18604 34196
rect 18656 34184 18662 34196
rect 18785 34187 18843 34193
rect 18785 34184 18797 34187
rect 18656 34156 18797 34184
rect 18656 34144 18662 34156
rect 18785 34153 18797 34156
rect 18831 34153 18843 34187
rect 18785 34147 18843 34153
rect 23842 34144 23848 34196
rect 23900 34184 23906 34196
rect 24397 34187 24455 34193
rect 24397 34184 24409 34187
rect 23900 34156 24409 34184
rect 23900 34144 23906 34156
rect 24397 34153 24409 34156
rect 24443 34153 24455 34187
rect 24397 34147 24455 34153
rect 27433 34187 27491 34193
rect 27433 34153 27445 34187
rect 27479 34184 27491 34187
rect 28350 34184 28356 34196
rect 27479 34156 28356 34184
rect 27479 34153 27491 34156
rect 27433 34147 27491 34153
rect 28350 34144 28356 34156
rect 28408 34144 28414 34196
rect 16574 34076 16580 34128
rect 16632 34116 16638 34128
rect 16632 34088 17816 34116
rect 16632 34076 16638 34088
rect 13814 34008 13820 34060
rect 13872 34048 13878 34060
rect 14461 34051 14519 34057
rect 14461 34048 14473 34051
rect 13872 34020 14473 34048
rect 13872 34008 13878 34020
rect 14461 34017 14473 34020
rect 14507 34017 14519 34051
rect 14461 34011 14519 34017
rect 14734 34008 14740 34060
rect 14792 34008 14798 34060
rect 17037 34051 17095 34057
rect 17037 34017 17049 34051
rect 17083 34048 17095 34051
rect 17126 34048 17132 34060
rect 17083 34020 17132 34048
rect 17083 34017 17095 34020
rect 17037 34011 17095 34017
rect 17126 34008 17132 34020
rect 17184 34008 17190 34060
rect 17788 34057 17816 34088
rect 18230 34076 18236 34128
rect 18288 34116 18294 34128
rect 18693 34119 18751 34125
rect 18693 34116 18705 34119
rect 18288 34088 18705 34116
rect 18288 34076 18294 34088
rect 18693 34085 18705 34088
rect 18739 34085 18751 34119
rect 18693 34079 18751 34085
rect 21542 34076 21548 34128
rect 21600 34116 21606 34128
rect 21637 34119 21695 34125
rect 21637 34116 21649 34119
rect 21600 34088 21649 34116
rect 21600 34076 21606 34088
rect 21637 34085 21649 34088
rect 21683 34085 21695 34119
rect 21637 34079 21695 34085
rect 17221 34051 17279 34057
rect 17221 34017 17233 34051
rect 17267 34048 17279 34051
rect 17589 34051 17647 34057
rect 17589 34048 17601 34051
rect 17267 34020 17601 34048
rect 17267 34017 17279 34020
rect 17221 34011 17279 34017
rect 17589 34017 17601 34020
rect 17635 34017 17647 34051
rect 17589 34011 17647 34017
rect 17773 34051 17831 34057
rect 17773 34017 17785 34051
rect 17819 34048 17831 34051
rect 17819 34020 18460 34048
rect 17819 34017 17831 34020
rect 17773 34011 17831 34017
rect 12897 33983 12955 33989
rect 12897 33980 12909 33983
rect 12636 33952 12909 33980
rect 12253 33943 12311 33949
rect 12897 33949 12909 33952
rect 12943 33949 12955 33983
rect 12897 33943 12955 33949
rect 11992 33912 12020 33943
rect 13078 33940 13084 33992
rect 13136 33940 13142 33992
rect 17402 33940 17408 33992
rect 17460 33940 17466 33992
rect 17497 33983 17555 33989
rect 17497 33949 17509 33983
rect 17543 33980 17555 33983
rect 17788 33980 17816 34011
rect 17543 33952 17816 33980
rect 17865 33983 17923 33989
rect 17543 33949 17555 33952
rect 17497 33943 17555 33949
rect 17865 33949 17877 33983
rect 17911 33949 17923 33983
rect 17865 33943 17923 33949
rect 12713 33915 12771 33921
rect 12713 33912 12725 33915
rect 10796 33884 12725 33912
rect 10100 33872 10106 33884
rect 12713 33881 12725 33884
rect 12759 33881 12771 33915
rect 12713 33875 12771 33881
rect 15010 33872 15016 33924
rect 15068 33912 15074 33924
rect 17420 33912 17448 33940
rect 17880 33912 17908 33943
rect 18138 33940 18144 33992
rect 18196 33940 18202 33992
rect 15068 33884 15226 33912
rect 17420 33884 17908 33912
rect 18432 33912 18460 34020
rect 18874 34008 18880 34060
rect 18932 34008 18938 34060
rect 20162 34008 20168 34060
rect 20220 34048 20226 34060
rect 20349 34051 20407 34057
rect 20349 34048 20361 34051
rect 20220 34020 20361 34048
rect 20220 34008 20226 34020
rect 20349 34017 20361 34020
rect 20395 34017 20407 34051
rect 20349 34011 20407 34017
rect 20898 34008 20904 34060
rect 20956 34048 20962 34060
rect 21913 34051 21971 34057
rect 21913 34048 21925 34051
rect 20956 34020 21925 34048
rect 20956 34008 20962 34020
rect 21913 34017 21925 34020
rect 21959 34017 21971 34051
rect 21913 34011 21971 34017
rect 25041 34051 25099 34057
rect 25041 34017 25053 34051
rect 25087 34048 25099 34051
rect 25130 34048 25136 34060
rect 25087 34020 25136 34048
rect 25087 34017 25099 34020
rect 25041 34011 25099 34017
rect 25130 34008 25136 34020
rect 25188 34048 25194 34060
rect 25866 34048 25872 34060
rect 25188 34020 25872 34048
rect 25188 34008 25194 34020
rect 25866 34008 25872 34020
rect 25924 34008 25930 34060
rect 28902 34008 28908 34060
rect 28960 34048 28966 34060
rect 29181 34051 29239 34057
rect 29181 34048 29193 34051
rect 28960 34020 29193 34048
rect 28960 34008 28966 34020
rect 29181 34017 29193 34020
rect 29227 34048 29239 34051
rect 29733 34051 29791 34057
rect 29733 34048 29745 34051
rect 29227 34020 29745 34048
rect 29227 34017 29239 34020
rect 29181 34011 29239 34017
rect 29733 34017 29745 34020
rect 29779 34048 29791 34051
rect 29914 34048 29920 34060
rect 29779 34020 29920 34048
rect 29779 34017 29791 34020
rect 29733 34011 29791 34017
rect 29914 34008 29920 34020
rect 29972 34008 29978 34060
rect 18506 33940 18512 33992
rect 18564 33980 18570 33992
rect 18601 33983 18659 33989
rect 18601 33980 18613 33983
rect 18564 33952 18613 33980
rect 18564 33940 18570 33952
rect 18601 33949 18613 33952
rect 18647 33949 18659 33983
rect 18601 33943 18659 33949
rect 20441 33983 20499 33989
rect 20441 33949 20453 33983
rect 20487 33980 20499 33983
rect 21818 33980 21824 33992
rect 20487 33952 21824 33980
rect 20487 33949 20499 33952
rect 20441 33943 20499 33949
rect 21818 33940 21824 33952
rect 21876 33940 21882 33992
rect 22005 33983 22063 33989
rect 22005 33949 22017 33983
rect 22051 33949 22063 33983
rect 22005 33943 22063 33949
rect 24857 33983 24915 33989
rect 24857 33949 24869 33983
rect 24903 33980 24915 33983
rect 25682 33980 25688 33992
rect 24903 33952 25688 33980
rect 24903 33949 24915 33952
rect 24857 33943 24915 33949
rect 18432 33884 20208 33912
rect 15068 33872 15074 33884
rect 11698 33844 11704 33856
rect 9968 33816 11704 33844
rect 11698 33804 11704 33816
rect 11756 33804 11762 33856
rect 16209 33847 16267 33853
rect 16209 33813 16221 33847
rect 16255 33844 16267 33847
rect 16298 33844 16304 33856
rect 16255 33816 16304 33844
rect 16255 33813 16267 33816
rect 16209 33807 16267 33813
rect 16298 33804 16304 33816
rect 16356 33804 16362 33856
rect 17586 33804 17592 33856
rect 17644 33804 17650 33856
rect 18322 33804 18328 33856
rect 18380 33844 18386 33856
rect 20073 33847 20131 33853
rect 20073 33844 20085 33847
rect 18380 33816 20085 33844
rect 18380 33804 18386 33816
rect 20073 33813 20085 33816
rect 20119 33813 20131 33847
rect 20180 33844 20208 33884
rect 21726 33872 21732 33924
rect 21784 33912 21790 33924
rect 22020 33912 22048 33943
rect 25682 33940 25688 33952
rect 25740 33940 25746 33992
rect 30101 33983 30159 33989
rect 30101 33949 30113 33983
rect 30147 33980 30159 33983
rect 30190 33980 30196 33992
rect 30147 33952 30196 33980
rect 30147 33949 30159 33952
rect 30101 33943 30159 33949
rect 30190 33940 30196 33952
rect 30248 33940 30254 33992
rect 32030 33940 32036 33992
rect 32088 33980 32094 33992
rect 32125 33983 32183 33989
rect 32125 33980 32137 33983
rect 32088 33952 32137 33980
rect 32088 33940 32094 33952
rect 32125 33949 32137 33952
rect 32171 33949 32183 33983
rect 32125 33943 32183 33949
rect 21784 33884 22048 33912
rect 21784 33872 21790 33884
rect 28350 33872 28356 33924
rect 28408 33872 28414 33924
rect 28905 33915 28963 33921
rect 28905 33881 28917 33915
rect 28951 33912 28963 33915
rect 29730 33912 29736 33924
rect 28951 33884 29736 33912
rect 28951 33881 28963 33884
rect 28905 33875 28963 33881
rect 29730 33872 29736 33884
rect 29788 33872 29794 33924
rect 30466 33872 30472 33924
rect 30524 33872 30530 33924
rect 32401 33915 32459 33921
rect 32401 33881 32413 33915
rect 32447 33912 32459 33915
rect 32674 33912 32680 33924
rect 32447 33884 32680 33912
rect 32447 33881 32459 33884
rect 32401 33875 32459 33881
rect 32674 33872 32680 33884
rect 32732 33872 32738 33924
rect 32784 33884 32890 33912
rect 24765 33847 24823 33853
rect 24765 33844 24777 33847
rect 20180 33816 24777 33844
rect 20073 33807 20131 33813
rect 24765 33813 24777 33816
rect 24811 33813 24823 33847
rect 24765 33807 24823 33813
rect 31386 33804 31392 33856
rect 31444 33844 31450 33856
rect 31527 33847 31585 33853
rect 31527 33844 31539 33847
rect 31444 33816 31539 33844
rect 31444 33804 31450 33816
rect 31527 33813 31539 33816
rect 31573 33813 31585 33847
rect 31527 33807 31585 33813
rect 32490 33804 32496 33856
rect 32548 33844 32554 33856
rect 32784 33844 32812 33884
rect 32548 33816 32812 33844
rect 33873 33847 33931 33853
rect 32548 33804 32554 33816
rect 33873 33813 33885 33847
rect 33919 33844 33931 33847
rect 34054 33844 34060 33856
rect 33919 33816 34060 33844
rect 33919 33813 33931 33816
rect 33873 33807 33931 33813
rect 34054 33804 34060 33816
rect 34112 33804 34118 33856
rect 1104 33754 40572 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 40572 33754
rect 1104 33680 40572 33702
rect 2222 33600 2228 33652
rect 2280 33640 2286 33652
rect 4154 33640 4160 33652
rect 2280 33612 4160 33640
rect 2280 33600 2286 33612
rect 4154 33600 4160 33612
rect 4212 33600 4218 33652
rect 5534 33600 5540 33652
rect 5592 33600 5598 33652
rect 5629 33643 5687 33649
rect 5629 33609 5641 33643
rect 5675 33640 5687 33643
rect 6365 33643 6423 33649
rect 6365 33640 6377 33643
rect 5675 33612 6377 33640
rect 5675 33609 5687 33612
rect 5629 33603 5687 33609
rect 6365 33609 6377 33612
rect 6411 33609 6423 33643
rect 6365 33603 6423 33609
rect 6733 33643 6791 33649
rect 6733 33609 6745 33643
rect 6779 33640 6791 33643
rect 8941 33643 8999 33649
rect 8941 33640 8953 33643
rect 6779 33612 8953 33640
rect 6779 33609 6791 33612
rect 6733 33603 6791 33609
rect 8941 33609 8953 33612
rect 8987 33609 8999 33643
rect 8941 33603 8999 33609
rect 9674 33600 9680 33652
rect 9732 33640 9738 33652
rect 9861 33643 9919 33649
rect 9861 33640 9873 33643
rect 9732 33612 9873 33640
rect 9732 33600 9738 33612
rect 9861 33609 9873 33612
rect 9907 33640 9919 33643
rect 9907 33612 10272 33640
rect 9907 33609 9919 33612
rect 9861 33603 9919 33609
rect 1486 33532 1492 33584
rect 1544 33572 1550 33584
rect 2317 33575 2375 33581
rect 2317 33572 2329 33575
rect 1544 33544 2329 33572
rect 1544 33532 1550 33544
rect 2317 33541 2329 33544
rect 2363 33541 2375 33575
rect 5552 33572 5580 33600
rect 2317 33535 2375 33541
rect 2746 33544 5580 33572
rect 6089 33575 6147 33581
rect 2222 33464 2228 33516
rect 2280 33464 2286 33516
rect 2501 33507 2559 33513
rect 2501 33473 2513 33507
rect 2547 33504 2559 33507
rect 2746 33504 2774 33544
rect 6089 33541 6101 33575
rect 6135 33572 6147 33575
rect 6638 33572 6644 33584
rect 6135 33544 6644 33572
rect 6135 33541 6147 33544
rect 6089 33535 6147 33541
rect 6638 33532 6644 33544
rect 6696 33532 6702 33584
rect 10137 33575 10195 33581
rect 10137 33572 10149 33575
rect 8036 33544 10149 33572
rect 2547 33476 2774 33504
rect 3145 33507 3203 33513
rect 2547 33473 2559 33476
rect 2501 33467 2559 33473
rect 3145 33473 3157 33507
rect 3191 33504 3203 33507
rect 5537 33507 5595 33513
rect 3191 33476 3372 33504
rect 3191 33473 3203 33476
rect 3145 33467 3203 33473
rect 1670 33396 1676 33448
rect 1728 33436 1734 33448
rect 3237 33439 3295 33445
rect 3237 33436 3249 33439
rect 1728 33408 3249 33436
rect 1728 33396 1734 33408
rect 3237 33405 3249 33408
rect 3283 33405 3295 33439
rect 3237 33399 3295 33405
rect 2685 33371 2743 33377
rect 2685 33337 2697 33371
rect 2731 33368 2743 33371
rect 2866 33368 2872 33380
rect 2731 33340 2872 33368
rect 2731 33337 2743 33340
rect 2685 33331 2743 33337
rect 2866 33328 2872 33340
rect 2924 33328 2930 33380
rect 3344 33368 3372 33476
rect 5537 33473 5549 33507
rect 5583 33504 5595 33507
rect 5626 33504 5632 33516
rect 5583 33476 5632 33504
rect 5583 33473 5595 33476
rect 5537 33467 5595 33473
rect 5626 33464 5632 33476
rect 5684 33464 5690 33516
rect 5994 33464 6000 33516
rect 6052 33464 6058 33516
rect 6181 33507 6239 33513
rect 6181 33473 6193 33507
rect 6227 33504 6239 33507
rect 6362 33504 6368 33516
rect 6227 33476 6368 33504
rect 6227 33473 6239 33476
rect 6181 33467 6239 33473
rect 6362 33464 6368 33476
rect 6420 33464 6426 33516
rect 7190 33464 7196 33516
rect 7248 33464 7254 33516
rect 7282 33464 7288 33516
rect 7340 33504 7346 33516
rect 7377 33507 7435 33513
rect 7377 33504 7389 33507
rect 7340 33476 7389 33504
rect 7340 33464 7346 33476
rect 7377 33473 7389 33476
rect 7423 33473 7435 33507
rect 7377 33467 7435 33473
rect 7834 33464 7840 33516
rect 7892 33464 7898 33516
rect 8036 33513 8064 33544
rect 10137 33541 10149 33544
rect 10183 33541 10195 33575
rect 10244 33572 10272 33612
rect 10318 33600 10324 33652
rect 10376 33640 10382 33652
rect 10413 33643 10471 33649
rect 10413 33640 10425 33643
rect 10376 33612 10425 33640
rect 10376 33600 10382 33612
rect 10413 33609 10425 33612
rect 10459 33609 10471 33643
rect 10413 33603 10471 33609
rect 14185 33643 14243 33649
rect 14185 33609 14197 33643
rect 14231 33640 14243 33643
rect 14274 33640 14280 33652
rect 14231 33612 14280 33640
rect 14231 33609 14243 33612
rect 14185 33603 14243 33609
rect 14274 33600 14280 33612
rect 14332 33600 14338 33652
rect 14734 33600 14740 33652
rect 14792 33640 14798 33652
rect 14792 33612 15516 33640
rect 14792 33600 14798 33612
rect 10244 33544 10364 33572
rect 10137 33535 10195 33541
rect 8021 33507 8079 33513
rect 8021 33473 8033 33507
rect 8067 33473 8079 33507
rect 8021 33467 8079 33473
rect 8297 33507 8355 33513
rect 8297 33473 8309 33507
rect 8343 33504 8355 33507
rect 8386 33504 8392 33516
rect 8343 33476 8392 33504
rect 8343 33473 8355 33476
rect 8297 33467 8355 33473
rect 8386 33464 8392 33476
rect 8444 33464 8450 33516
rect 8478 33464 8484 33516
rect 8536 33464 8542 33516
rect 9030 33464 9036 33516
rect 9088 33504 9094 33516
rect 9401 33507 9459 33513
rect 9401 33504 9413 33507
rect 9088 33476 9413 33504
rect 9088 33464 9094 33476
rect 9401 33473 9413 33476
rect 9447 33473 9459 33507
rect 9401 33467 9459 33473
rect 9582 33464 9588 33516
rect 9640 33464 9646 33516
rect 9677 33507 9735 33513
rect 9677 33473 9689 33507
rect 9723 33504 9735 33507
rect 9723 33476 9757 33504
rect 9723 33473 9735 33476
rect 9677 33467 9735 33473
rect 3421 33439 3479 33445
rect 3421 33405 3433 33439
rect 3467 33436 3479 33439
rect 4154 33436 4160 33448
rect 3467 33408 4160 33436
rect 3467 33405 3479 33408
rect 3421 33399 3479 33405
rect 4154 33396 4160 33408
rect 4212 33396 4218 33448
rect 5810 33396 5816 33448
rect 5868 33436 5874 33448
rect 5868 33408 6776 33436
rect 5868 33396 5874 33408
rect 6086 33368 6092 33380
rect 3344 33340 6092 33368
rect 6086 33328 6092 33340
rect 6144 33328 6150 33380
rect 6748 33368 6776 33408
rect 6822 33396 6828 33448
rect 6880 33396 6886 33448
rect 6917 33439 6975 33445
rect 6917 33405 6929 33439
rect 6963 33436 6975 33439
rect 7098 33436 7104 33448
rect 6963 33408 7104 33436
rect 6963 33405 6975 33408
rect 6917 33399 6975 33405
rect 7098 33396 7104 33408
rect 7156 33436 7162 33448
rect 7466 33436 7472 33448
rect 7156 33408 7472 33436
rect 7156 33396 7162 33408
rect 7466 33396 7472 33408
rect 7524 33396 7530 33448
rect 8113 33439 8171 33445
rect 8113 33405 8125 33439
rect 8159 33436 8171 33439
rect 8662 33436 8668 33448
rect 8159 33408 8668 33436
rect 8159 33405 8171 33408
rect 8113 33399 8171 33405
rect 8662 33396 8668 33408
rect 8720 33396 8726 33448
rect 8938 33396 8944 33448
rect 8996 33436 9002 33448
rect 9692 33436 9720 33467
rect 10042 33464 10048 33516
rect 10100 33464 10106 33516
rect 10226 33464 10232 33516
rect 10284 33464 10290 33516
rect 10336 33513 10364 33544
rect 15286 33532 15292 33584
rect 15344 33532 15350 33584
rect 15488 33581 15516 33612
rect 15654 33600 15660 33652
rect 15712 33640 15718 33652
rect 16390 33640 16396 33652
rect 15712 33612 16396 33640
rect 15712 33600 15718 33612
rect 16390 33600 16396 33612
rect 16448 33600 16454 33652
rect 16666 33600 16672 33652
rect 16724 33640 16730 33652
rect 18138 33640 18144 33652
rect 16724 33612 18144 33640
rect 16724 33600 16730 33612
rect 18138 33600 18144 33612
rect 18196 33600 18202 33652
rect 18230 33600 18236 33652
rect 18288 33640 18294 33652
rect 18598 33640 18604 33652
rect 18288 33612 18604 33640
rect 18288 33600 18294 33612
rect 18598 33600 18604 33612
rect 18656 33600 18662 33652
rect 20162 33600 20168 33652
rect 20220 33600 20226 33652
rect 29730 33600 29736 33652
rect 29788 33640 29794 33652
rect 30101 33643 30159 33649
rect 30101 33640 30113 33643
rect 29788 33612 30113 33640
rect 29788 33600 29794 33612
rect 30101 33609 30113 33612
rect 30147 33609 30159 33643
rect 30101 33603 30159 33609
rect 30190 33600 30196 33652
rect 30248 33600 30254 33652
rect 32674 33600 32680 33652
rect 32732 33600 32738 33652
rect 15473 33575 15531 33581
rect 15473 33541 15485 33575
rect 15519 33572 15531 33575
rect 16114 33572 16120 33584
rect 15519 33544 16120 33572
rect 15519 33541 15531 33544
rect 15473 33535 15531 33541
rect 16114 33532 16120 33544
rect 16172 33572 16178 33584
rect 17126 33572 17132 33584
rect 16172 33544 17132 33572
rect 16172 33532 16178 33544
rect 17126 33532 17132 33544
rect 17184 33532 17190 33584
rect 19242 33572 19248 33584
rect 19182 33558 19248 33572
rect 19168 33544 19248 33558
rect 10321 33507 10379 33513
rect 10321 33473 10333 33507
rect 10367 33473 10379 33507
rect 10321 33467 10379 33473
rect 10505 33507 10563 33513
rect 10505 33473 10517 33507
rect 10551 33473 10563 33507
rect 10505 33467 10563 33473
rect 8996 33408 9904 33436
rect 8996 33396 9002 33408
rect 7006 33368 7012 33380
rect 6748 33340 7012 33368
rect 7006 33328 7012 33340
rect 7064 33328 7070 33380
rect 7285 33371 7343 33377
rect 7285 33337 7297 33371
rect 7331 33368 7343 33371
rect 7374 33368 7380 33380
rect 7331 33340 7380 33368
rect 7331 33337 7343 33340
rect 7285 33331 7343 33337
rect 7374 33328 7380 33340
rect 7432 33328 7438 33380
rect 9125 33371 9183 33377
rect 9125 33337 9137 33371
rect 9171 33368 9183 33371
rect 9766 33368 9772 33380
rect 9171 33340 9772 33368
rect 9171 33337 9183 33340
rect 9125 33331 9183 33337
rect 9766 33328 9772 33340
rect 9824 33328 9830 33380
rect 9876 33368 9904 33408
rect 10134 33396 10140 33448
rect 10192 33436 10198 33448
rect 10520 33436 10548 33467
rect 13078 33464 13084 33516
rect 13136 33504 13142 33516
rect 14553 33507 14611 33513
rect 14553 33504 14565 33507
rect 13136 33476 14565 33504
rect 13136 33464 13142 33476
rect 14553 33473 14565 33476
rect 14599 33504 14611 33507
rect 14599 33476 14872 33504
rect 14599 33473 14611 33476
rect 14553 33467 14611 33473
rect 14645 33439 14703 33445
rect 14645 33436 14657 33439
rect 10192 33408 10548 33436
rect 12406 33408 14657 33436
rect 10192 33396 10198 33408
rect 11146 33368 11152 33380
rect 9876 33340 11152 33368
rect 11146 33328 11152 33340
rect 11204 33328 11210 33380
rect 2777 33303 2835 33309
rect 2777 33269 2789 33303
rect 2823 33300 2835 33303
rect 3602 33300 3608 33312
rect 2823 33272 3608 33300
rect 2823 33269 2835 33272
rect 2777 33263 2835 33269
rect 3602 33260 3608 33272
rect 3660 33260 3666 33312
rect 5166 33260 5172 33312
rect 5224 33260 5230 33312
rect 7650 33260 7656 33312
rect 7708 33260 7714 33312
rect 9030 33260 9036 33312
rect 9088 33300 9094 33312
rect 12406 33300 12434 33408
rect 14645 33405 14657 33408
rect 14691 33405 14703 33439
rect 14645 33399 14703 33405
rect 14734 33396 14740 33448
rect 14792 33396 14798 33448
rect 14844 33436 14872 33476
rect 16298 33436 16304 33448
rect 14844 33408 16304 33436
rect 16298 33396 16304 33408
rect 16356 33396 16362 33448
rect 17218 33396 17224 33448
rect 17276 33436 17282 33448
rect 17678 33436 17684 33448
rect 17276 33408 17684 33436
rect 17276 33396 17282 33408
rect 17678 33396 17684 33408
rect 17736 33396 17742 33448
rect 17954 33396 17960 33448
rect 18012 33396 18018 33448
rect 18506 33396 18512 33448
rect 18564 33436 18570 33448
rect 19168 33436 19196 33544
rect 19242 33532 19248 33544
rect 19300 33532 19306 33584
rect 28350 33572 28356 33584
rect 28014 33544 28356 33572
rect 28350 33532 28356 33544
rect 28408 33532 28414 33584
rect 28994 33532 29000 33584
rect 29052 33572 29058 33584
rect 29825 33575 29883 33581
rect 29825 33572 29837 33575
rect 29052 33544 29837 33572
rect 29052 33532 29058 33544
rect 29825 33541 29837 33544
rect 29871 33541 29883 33575
rect 29825 33535 29883 33541
rect 33045 33575 33103 33581
rect 33045 33541 33057 33575
rect 33091 33572 33103 33575
rect 33505 33575 33563 33581
rect 33505 33572 33517 33575
rect 33091 33544 33517 33572
rect 33091 33541 33103 33544
rect 33045 33535 33103 33541
rect 33505 33541 33517 33544
rect 33551 33541 33563 33575
rect 34425 33575 34483 33581
rect 34425 33572 34437 33575
rect 33505 33535 33563 33541
rect 34072 33544 34437 33572
rect 34072 33516 34100 33544
rect 34425 33541 34437 33544
rect 34471 33541 34483 33575
rect 34425 33535 34483 33541
rect 19797 33507 19855 33513
rect 19797 33504 19809 33507
rect 18564 33408 19196 33436
rect 19444 33476 19809 33504
rect 18564 33396 18570 33408
rect 9088 33272 12434 33300
rect 9088 33260 9094 33272
rect 18138 33260 18144 33312
rect 18196 33300 18202 33312
rect 19444 33309 19472 33476
rect 19797 33473 19809 33476
rect 19843 33473 19855 33507
rect 19797 33467 19855 33473
rect 28721 33507 28779 33513
rect 28721 33473 28733 33507
rect 28767 33504 28779 33507
rect 28902 33504 28908 33516
rect 28767 33476 28908 33504
rect 28767 33473 28779 33476
rect 28721 33467 28779 33473
rect 28902 33464 28908 33476
rect 28960 33464 28966 33516
rect 29546 33464 29552 33516
rect 29604 33464 29610 33516
rect 29638 33464 29644 33516
rect 29696 33504 29702 33516
rect 29733 33507 29791 33513
rect 29733 33504 29745 33507
rect 29696 33476 29745 33504
rect 29696 33464 29702 33476
rect 29733 33473 29745 33476
rect 29779 33473 29791 33507
rect 29733 33467 29791 33473
rect 29917 33507 29975 33513
rect 29917 33473 29929 33507
rect 29963 33504 29975 33507
rect 30469 33507 30527 33513
rect 29963 33476 30420 33504
rect 29963 33473 29975 33476
rect 29917 33467 29975 33473
rect 19702 33396 19708 33448
rect 19760 33396 19766 33448
rect 28442 33396 28448 33448
rect 28500 33396 28506 33448
rect 28813 33439 28871 33445
rect 28813 33436 28825 33439
rect 28644 33408 28825 33436
rect 19429 33303 19487 33309
rect 19429 33300 19441 33303
rect 18196 33272 19441 33300
rect 18196 33260 18202 33272
rect 19429 33269 19441 33272
rect 19475 33269 19487 33303
rect 19429 33263 19487 33269
rect 19886 33260 19892 33312
rect 19944 33300 19950 33312
rect 24394 33300 24400 33312
rect 19944 33272 24400 33300
rect 19944 33260 19950 33272
rect 24394 33260 24400 33272
rect 24452 33260 24458 33312
rect 26973 33303 27031 33309
rect 26973 33269 26985 33303
rect 27019 33300 27031 33303
rect 28074 33300 28080 33312
rect 27019 33272 28080 33300
rect 27019 33269 27031 33272
rect 26973 33263 27031 33269
rect 28074 33260 28080 33272
rect 28132 33300 28138 33312
rect 28644 33300 28672 33408
rect 28813 33405 28825 33408
rect 28859 33405 28871 33439
rect 28813 33399 28871 33405
rect 28994 33396 29000 33448
rect 29052 33436 29058 33448
rect 29656 33436 29684 33464
rect 29052 33408 29684 33436
rect 29052 33396 29058 33408
rect 29086 33328 29092 33380
rect 29144 33368 29150 33380
rect 29932 33368 29960 33467
rect 30098 33396 30104 33448
rect 30156 33436 30162 33448
rect 30193 33439 30251 33445
rect 30193 33436 30205 33439
rect 30156 33408 30205 33436
rect 30156 33396 30162 33408
rect 30193 33405 30205 33408
rect 30239 33405 30251 33439
rect 30193 33399 30251 33405
rect 29144 33340 29960 33368
rect 29144 33328 29150 33340
rect 28132 33272 28672 33300
rect 28132 33260 28138 33272
rect 29454 33260 29460 33312
rect 29512 33260 29518 33312
rect 30392 33309 30420 33476
rect 30469 33473 30481 33507
rect 30515 33504 30527 33507
rect 30745 33507 30803 33513
rect 30745 33504 30757 33507
rect 30515 33476 30757 33504
rect 30515 33473 30527 33476
rect 30469 33467 30527 33473
rect 30745 33473 30757 33476
rect 30791 33473 30803 33507
rect 30745 33467 30803 33473
rect 31386 33464 31392 33516
rect 31444 33464 31450 33516
rect 31938 33464 31944 33516
rect 31996 33464 32002 33516
rect 32861 33507 32919 33513
rect 32861 33473 32873 33507
rect 32907 33473 32919 33507
rect 32861 33467 32919 33473
rect 31665 33439 31723 33445
rect 31665 33405 31677 33439
rect 31711 33405 31723 33439
rect 32876 33436 32904 33467
rect 32950 33464 32956 33516
rect 33008 33504 33014 33516
rect 33137 33507 33195 33513
rect 33137 33504 33149 33507
rect 33008 33476 33149 33504
rect 33008 33464 33014 33476
rect 33137 33473 33149 33476
rect 33183 33473 33195 33507
rect 33137 33467 33195 33473
rect 34054 33464 34060 33516
rect 34112 33464 34118 33516
rect 34238 33464 34244 33516
rect 34296 33464 34302 33516
rect 38746 33436 38752 33448
rect 32876 33408 38752 33436
rect 31665 33399 31723 33405
rect 30742 33328 30748 33380
rect 30800 33368 30806 33380
rect 31680 33368 31708 33399
rect 38746 33396 38752 33408
rect 38804 33396 38810 33448
rect 30800 33340 31708 33368
rect 30800 33328 30806 33340
rect 30377 33303 30435 33309
rect 30377 33269 30389 33303
rect 30423 33300 30435 33303
rect 31018 33300 31024 33312
rect 30423 33272 31024 33300
rect 30423 33269 30435 33272
rect 30377 33263 30435 33269
rect 31018 33260 31024 33272
rect 31076 33260 31082 33312
rect 33134 33260 33140 33312
rect 33192 33300 33198 33312
rect 34609 33303 34667 33309
rect 34609 33300 34621 33303
rect 33192 33272 34621 33300
rect 33192 33260 33198 33272
rect 34609 33269 34621 33272
rect 34655 33269 34667 33303
rect 34609 33263 34667 33269
rect 1104 33210 40572 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 40572 33210
rect 1104 33136 40572 33158
rect 3786 33056 3792 33108
rect 3844 33096 3850 33108
rect 3844 33068 5212 33096
rect 3844 33056 3850 33068
rect 5184 33028 5212 33068
rect 5626 33056 5632 33108
rect 5684 33056 5690 33108
rect 8386 33096 8392 33108
rect 5736 33068 8392 33096
rect 5736 33028 5764 33068
rect 8386 33056 8392 33068
rect 8444 33056 8450 33108
rect 8665 33099 8723 33105
rect 8665 33065 8677 33099
rect 8711 33096 8723 33099
rect 9214 33096 9220 33108
rect 8711 33068 9220 33096
rect 8711 33065 8723 33068
rect 8665 33059 8723 33065
rect 9214 33056 9220 33068
rect 9272 33096 9278 33108
rect 9582 33096 9588 33108
rect 9272 33068 9588 33096
rect 9272 33056 9278 33068
rect 9582 33056 9588 33068
rect 9640 33056 9646 33108
rect 15286 33056 15292 33108
rect 15344 33096 15350 33108
rect 15565 33099 15623 33105
rect 15565 33096 15577 33099
rect 15344 33068 15577 33096
rect 15344 33056 15350 33068
rect 15565 33065 15577 33068
rect 15611 33065 15623 33099
rect 16393 33099 16451 33105
rect 16393 33096 16405 33099
rect 15565 33059 15623 33065
rect 16040 33068 16405 33096
rect 5184 33000 5764 33028
rect 12434 32988 12440 33040
rect 12492 33028 12498 33040
rect 15838 33028 15844 33040
rect 12492 33000 15844 33028
rect 12492 32988 12498 33000
rect 15838 32988 15844 33000
rect 15896 32988 15902 33040
rect 2866 32920 2872 32972
rect 2924 32960 2930 32972
rect 3237 32963 3295 32969
rect 3237 32960 3249 32963
rect 2924 32932 3249 32960
rect 2924 32920 2930 32932
rect 3237 32929 3249 32932
rect 3283 32929 3295 32963
rect 3237 32923 3295 32929
rect 4157 32963 4215 32969
rect 4157 32929 4169 32963
rect 4203 32960 4215 32963
rect 5166 32960 5172 32972
rect 4203 32932 5172 32960
rect 4203 32929 4215 32932
rect 4157 32923 4215 32929
rect 5166 32920 5172 32932
rect 5224 32920 5230 32972
rect 6546 32920 6552 32972
rect 6604 32960 6610 32972
rect 6641 32963 6699 32969
rect 6641 32960 6653 32963
rect 6604 32932 6653 32960
rect 6604 32920 6610 32932
rect 6641 32929 6653 32932
rect 6687 32929 6699 32963
rect 6641 32923 6699 32929
rect 6914 32920 6920 32972
rect 6972 32920 6978 32972
rect 7193 32963 7251 32969
rect 7193 32929 7205 32963
rect 7239 32960 7251 32963
rect 7650 32960 7656 32972
rect 7239 32932 7656 32960
rect 7239 32929 7251 32932
rect 7193 32923 7251 32929
rect 7650 32920 7656 32932
rect 7708 32920 7714 32972
rect 8386 32920 8392 32972
rect 8444 32920 8450 32972
rect 8662 32920 8668 32972
rect 8720 32960 8726 32972
rect 8720 32932 15608 32960
rect 8720 32920 8726 32932
rect 3513 32895 3571 32901
rect 3513 32861 3525 32895
rect 3559 32892 3571 32895
rect 3878 32892 3884 32904
rect 3559 32864 3884 32892
rect 3559 32861 3571 32864
rect 3513 32855 3571 32861
rect 3878 32852 3884 32864
rect 3936 32852 3942 32904
rect 8404 32892 8432 32920
rect 15580 32904 15608 32932
rect 8326 32864 8432 32892
rect 10594 32852 10600 32904
rect 10652 32892 10658 32904
rect 11609 32895 11667 32901
rect 11609 32892 11621 32895
rect 10652 32864 11621 32892
rect 10652 32852 10658 32864
rect 11609 32861 11621 32864
rect 11655 32861 11667 32895
rect 11609 32855 11667 32861
rect 11701 32895 11759 32901
rect 11701 32861 11713 32895
rect 11747 32892 11759 32895
rect 12526 32892 12532 32904
rect 11747 32864 12532 32892
rect 11747 32861 11759 32864
rect 11701 32855 11759 32861
rect 12526 32852 12532 32864
rect 12584 32852 12590 32904
rect 15562 32852 15568 32904
rect 15620 32852 15626 32904
rect 15749 32895 15807 32901
rect 15749 32861 15761 32895
rect 15795 32892 15807 32895
rect 16040 32892 16068 33068
rect 16393 33065 16405 33068
rect 16439 33065 16451 33099
rect 16393 33059 16451 33065
rect 16408 33028 16436 33059
rect 17954 33056 17960 33108
rect 18012 33096 18018 33108
rect 18325 33099 18383 33105
rect 18325 33096 18337 33099
rect 18012 33068 18337 33096
rect 18012 33056 18018 33068
rect 18325 33065 18337 33068
rect 18371 33065 18383 33099
rect 18325 33059 18383 33065
rect 28442 33056 28448 33108
rect 28500 33096 28506 33108
rect 28537 33099 28595 33105
rect 28537 33096 28549 33099
rect 28500 33068 28549 33096
rect 28500 33056 28506 33068
rect 28537 33065 28549 33068
rect 28583 33065 28595 33099
rect 28537 33059 28595 33065
rect 29546 33056 29552 33108
rect 29604 33096 29610 33108
rect 29641 33099 29699 33105
rect 29641 33096 29653 33099
rect 29604 33068 29653 33096
rect 29604 33056 29610 33068
rect 29641 33065 29653 33068
rect 29687 33065 29699 33099
rect 29641 33059 29699 33065
rect 29730 33056 29736 33108
rect 29788 33096 29794 33108
rect 29788 33068 33180 33096
rect 29788 33056 29794 33068
rect 22554 33028 22560 33040
rect 16408 33000 22560 33028
rect 22554 32988 22560 33000
rect 22612 32988 22618 33040
rect 33152 33028 33180 33068
rect 33226 33056 33232 33108
rect 33284 33096 33290 33108
rect 33551 33099 33609 33105
rect 33551 33096 33563 33099
rect 33284 33068 33563 33096
rect 33284 33056 33290 33068
rect 33551 33065 33563 33068
rect 33597 33096 33609 33099
rect 34238 33096 34244 33108
rect 33597 33068 34244 33096
rect 33597 33065 33609 33068
rect 33551 33059 33609 33065
rect 34238 33056 34244 33068
rect 34296 33056 34302 33108
rect 34330 33028 34336 33040
rect 33152 33000 34336 33028
rect 34330 32988 34336 33000
rect 34388 33028 34394 33040
rect 34388 33000 34744 33028
rect 34388 32988 34394 33000
rect 18322 32960 18328 32972
rect 17788 32932 18328 32960
rect 15795 32864 16068 32892
rect 15795 32861 15807 32864
rect 15749 32855 15807 32861
rect 16114 32852 16120 32904
rect 16172 32892 16178 32904
rect 16301 32895 16359 32901
rect 16301 32892 16313 32895
rect 16172 32864 16313 32892
rect 16172 32852 16178 32864
rect 16301 32861 16313 32864
rect 16347 32861 16359 32895
rect 16301 32855 16359 32861
rect 16482 32852 16488 32904
rect 16540 32852 16546 32904
rect 17586 32852 17592 32904
rect 17644 32852 17650 32904
rect 17788 32901 17816 32932
rect 18322 32920 18328 32932
rect 18380 32920 18386 32972
rect 26786 32960 26792 32972
rect 25700 32932 26792 32960
rect 17773 32895 17831 32901
rect 17773 32861 17785 32895
rect 17819 32861 17831 32895
rect 17773 32855 17831 32861
rect 17865 32895 17923 32901
rect 17865 32861 17877 32895
rect 17911 32861 17923 32895
rect 17865 32855 17923 32861
rect 17957 32895 18015 32901
rect 17957 32861 17969 32895
rect 18003 32861 18015 32895
rect 17957 32855 18015 32861
rect 1486 32784 1492 32836
rect 1544 32784 1550 32836
rect 2774 32784 2780 32836
rect 2832 32824 2838 32836
rect 2832 32796 3188 32824
rect 2832 32784 2838 32796
rect 3160 32756 3188 32796
rect 3344 32796 4646 32824
rect 3344 32756 3372 32796
rect 5534 32784 5540 32836
rect 5592 32824 5598 32836
rect 6270 32824 6276 32836
rect 5592 32796 6276 32824
rect 5592 32784 5598 32796
rect 6270 32784 6276 32796
rect 6328 32784 6334 32836
rect 6457 32827 6515 32833
rect 6457 32793 6469 32827
rect 6503 32824 6515 32827
rect 7282 32824 7288 32836
rect 6503 32796 7288 32824
rect 6503 32793 6515 32796
rect 6457 32787 6515 32793
rect 7282 32784 7288 32796
rect 7340 32784 7346 32836
rect 16666 32824 16672 32836
rect 16132 32796 16672 32824
rect 3160 32728 3372 32756
rect 5810 32716 5816 32768
rect 5868 32756 5874 32768
rect 6089 32759 6147 32765
rect 6089 32756 6101 32759
rect 5868 32728 6101 32756
rect 5868 32716 5874 32728
rect 6089 32725 6101 32728
rect 6135 32725 6147 32759
rect 6089 32719 6147 32725
rect 6546 32716 6552 32768
rect 6604 32716 6610 32768
rect 11054 32716 11060 32768
rect 11112 32756 11118 32768
rect 11241 32759 11299 32765
rect 11241 32756 11253 32759
rect 11112 32728 11253 32756
rect 11112 32716 11118 32728
rect 11241 32725 11253 32728
rect 11287 32725 11299 32759
rect 11241 32719 11299 32725
rect 11885 32759 11943 32765
rect 11885 32725 11897 32759
rect 11931 32756 11943 32759
rect 16022 32756 16028 32768
rect 11931 32728 16028 32756
rect 11931 32725 11943 32728
rect 11885 32719 11943 32725
rect 16022 32716 16028 32728
rect 16080 32716 16086 32768
rect 16132 32765 16160 32796
rect 16666 32784 16672 32796
rect 16724 32784 16730 32836
rect 16117 32759 16175 32765
rect 16117 32725 16129 32759
rect 16163 32725 16175 32759
rect 16117 32719 16175 32725
rect 16390 32716 16396 32768
rect 16448 32756 16454 32768
rect 17880 32756 17908 32855
rect 17972 32824 18000 32855
rect 18138 32852 18144 32904
rect 18196 32852 18202 32904
rect 18230 32852 18236 32904
rect 18288 32892 18294 32904
rect 23937 32895 23995 32901
rect 18288 32864 23888 32892
rect 18288 32852 18294 32864
rect 18598 32824 18604 32836
rect 17972 32796 18604 32824
rect 18598 32784 18604 32796
rect 18656 32784 18662 32836
rect 23658 32784 23664 32836
rect 23716 32784 23722 32836
rect 23860 32824 23888 32864
rect 23937 32861 23949 32895
rect 23983 32892 23995 32895
rect 24118 32892 24124 32904
rect 23983 32864 24124 32892
rect 23983 32861 23995 32864
rect 23937 32855 23995 32861
rect 24118 32852 24124 32864
rect 24176 32892 24182 32904
rect 24670 32892 24676 32904
rect 24176 32864 24676 32892
rect 24176 32852 24182 32864
rect 24670 32852 24676 32864
rect 24728 32852 24734 32904
rect 25700 32901 25728 32932
rect 26786 32920 26792 32932
rect 26844 32920 26850 32972
rect 28902 32960 28908 32972
rect 28644 32932 28908 32960
rect 25685 32895 25743 32901
rect 25685 32861 25697 32895
rect 25731 32861 25743 32895
rect 25685 32855 25743 32861
rect 25774 32852 25780 32904
rect 25832 32892 25838 32904
rect 26142 32901 26148 32904
rect 25961 32895 26019 32901
rect 25961 32892 25973 32895
rect 25832 32864 25973 32892
rect 25832 32852 25838 32864
rect 25961 32861 25973 32864
rect 26007 32861 26019 32895
rect 25961 32855 26019 32861
rect 26115 32895 26148 32901
rect 26115 32861 26127 32895
rect 26115 32855 26148 32861
rect 26142 32852 26148 32855
rect 26200 32852 26206 32904
rect 28644 32892 28672 32932
rect 28902 32920 28908 32932
rect 28960 32920 28966 32972
rect 29181 32963 29239 32969
rect 29181 32929 29193 32963
rect 29227 32960 29239 32963
rect 29454 32960 29460 32972
rect 29227 32932 29460 32960
rect 29227 32929 29239 32932
rect 29181 32923 29239 32929
rect 29454 32920 29460 32932
rect 29512 32920 29518 32972
rect 29914 32920 29920 32972
rect 29972 32960 29978 32972
rect 30190 32960 30196 32972
rect 29972 32932 30196 32960
rect 29972 32920 29978 32932
rect 30190 32920 30196 32932
rect 30248 32920 30254 32972
rect 31757 32963 31815 32969
rect 31757 32929 31769 32963
rect 31803 32960 31815 32963
rect 32030 32960 32036 32972
rect 31803 32932 32036 32960
rect 31803 32929 31815 32932
rect 31757 32923 31815 32929
rect 32030 32920 32036 32932
rect 32088 32960 32094 32972
rect 32088 32932 34652 32960
rect 32088 32920 32094 32932
rect 33704 32904 33732 32932
rect 28721 32895 28779 32901
rect 28721 32892 28733 32895
rect 28644 32864 28733 32892
rect 28721 32861 28733 32864
rect 28767 32861 28779 32895
rect 28721 32855 28779 32861
rect 28810 32852 28816 32904
rect 28868 32852 28874 32904
rect 29086 32901 29092 32904
rect 29043 32895 29092 32901
rect 29043 32861 29055 32895
rect 29089 32861 29092 32895
rect 29043 32855 29092 32861
rect 29086 32852 29092 32855
rect 29144 32852 29150 32904
rect 29546 32852 29552 32904
rect 29604 32852 29610 32904
rect 29733 32895 29791 32901
rect 29733 32861 29745 32895
rect 29779 32861 29791 32895
rect 29733 32855 29791 32861
rect 32125 32895 32183 32901
rect 32125 32861 32137 32895
rect 32171 32892 32183 32895
rect 32214 32892 32220 32904
rect 32171 32864 32220 32892
rect 32171 32861 32183 32864
rect 32125 32855 32183 32861
rect 28905 32827 28963 32833
rect 28905 32824 28917 32827
rect 23860 32796 28917 32824
rect 28905 32793 28917 32796
rect 28951 32824 28963 32827
rect 29564 32824 29592 32852
rect 28951 32796 29592 32824
rect 28951 32793 28963 32796
rect 28905 32787 28963 32793
rect 16448 32728 17908 32756
rect 16448 32716 16454 32728
rect 23750 32716 23756 32768
rect 23808 32765 23814 32768
rect 23808 32719 23817 32765
rect 23845 32759 23903 32765
rect 23845 32725 23857 32759
rect 23891 32756 23903 32759
rect 25038 32756 25044 32768
rect 23891 32728 25044 32756
rect 23891 32725 23903 32728
rect 23845 32719 23903 32725
rect 23808 32716 23814 32719
rect 25038 32716 25044 32728
rect 25096 32716 25102 32768
rect 25501 32759 25559 32765
rect 25501 32725 25513 32759
rect 25547 32756 25559 32759
rect 25590 32756 25596 32768
rect 25547 32728 25596 32756
rect 25547 32725 25559 32728
rect 25501 32719 25559 32725
rect 25590 32716 25596 32728
rect 25648 32716 25654 32768
rect 26329 32759 26387 32765
rect 26329 32725 26341 32759
rect 26375 32756 26387 32759
rect 26418 32756 26424 32768
rect 26375 32728 26424 32756
rect 26375 32725 26387 32728
rect 26329 32719 26387 32725
rect 26418 32716 26424 32728
rect 26476 32716 26482 32768
rect 28810 32716 28816 32768
rect 28868 32756 28874 32768
rect 29748 32756 29776 32855
rect 32214 32852 32220 32864
rect 32272 32852 32278 32904
rect 33686 32852 33692 32904
rect 33744 32852 33750 32904
rect 30193 32827 30251 32833
rect 30193 32793 30205 32827
rect 30239 32824 30251 32827
rect 30466 32824 30472 32836
rect 30239 32796 30472 32824
rect 30239 32793 30251 32796
rect 30193 32787 30251 32793
rect 30466 32784 30472 32796
rect 30524 32784 30530 32836
rect 30926 32784 30932 32836
rect 30984 32784 30990 32836
rect 32490 32784 32496 32836
rect 32548 32784 32554 32836
rect 34333 32827 34391 32833
rect 34333 32793 34345 32827
rect 34379 32793 34391 32827
rect 34624 32824 34652 32932
rect 34716 32901 34744 33000
rect 34900 32932 36768 32960
rect 34701 32895 34759 32901
rect 34701 32861 34713 32895
rect 34747 32861 34759 32895
rect 34701 32855 34759 32861
rect 34900 32824 34928 32932
rect 36740 32901 36768 32932
rect 36725 32895 36783 32901
rect 36725 32861 36737 32895
rect 36771 32892 36783 32895
rect 37274 32892 37280 32904
rect 36771 32864 37280 32892
rect 36771 32861 36783 32864
rect 36725 32855 36783 32861
rect 37274 32852 37280 32864
rect 37332 32852 37338 32904
rect 34624 32796 34928 32824
rect 34333 32787 34391 32793
rect 30282 32756 30288 32768
rect 28868 32728 30288 32756
rect 28868 32716 28874 32728
rect 30282 32716 30288 32728
rect 30340 32716 30346 32768
rect 31662 32716 31668 32768
rect 31720 32716 31726 32768
rect 32398 32716 32404 32768
rect 32456 32756 32462 32768
rect 34348 32756 34376 32787
rect 35986 32784 35992 32836
rect 36044 32824 36050 32836
rect 36044 32796 36216 32824
rect 36044 32784 36050 32796
rect 32456 32728 34376 32756
rect 32456 32716 32462 32728
rect 34422 32716 34428 32768
rect 34480 32716 34486 32768
rect 36188 32756 36216 32796
rect 36446 32784 36452 32836
rect 36504 32784 36510 32836
rect 39666 32756 39672 32768
rect 36188 32728 39672 32756
rect 39666 32716 39672 32728
rect 39724 32716 39730 32768
rect 1104 32666 40572 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 40572 32666
rect 1104 32592 40572 32614
rect 5353 32555 5411 32561
rect 5353 32521 5365 32555
rect 5399 32552 5411 32555
rect 5534 32552 5540 32564
rect 5399 32524 5540 32552
rect 5399 32521 5411 32524
rect 5353 32515 5411 32521
rect 5534 32512 5540 32524
rect 5592 32512 5598 32564
rect 6089 32555 6147 32561
rect 6089 32521 6101 32555
rect 6135 32552 6147 32555
rect 6822 32552 6828 32564
rect 6135 32524 6828 32552
rect 6135 32521 6147 32524
rect 6089 32515 6147 32521
rect 6822 32512 6828 32524
rect 6880 32512 6886 32564
rect 7374 32512 7380 32564
rect 7432 32512 7438 32564
rect 7561 32555 7619 32561
rect 7561 32521 7573 32555
rect 7607 32552 7619 32555
rect 7834 32552 7840 32564
rect 7607 32524 7840 32552
rect 7607 32521 7619 32524
rect 7561 32515 7619 32521
rect 7834 32512 7840 32524
rect 7892 32512 7898 32564
rect 12526 32512 12532 32564
rect 12584 32552 12590 32564
rect 12897 32555 12955 32561
rect 12897 32552 12909 32555
rect 12584 32524 12909 32552
rect 12584 32512 12590 32524
rect 12897 32521 12909 32524
rect 12943 32521 12955 32555
rect 12897 32515 12955 32521
rect 15838 32512 15844 32564
rect 15896 32552 15902 32564
rect 18138 32552 18144 32564
rect 15896 32524 18144 32552
rect 15896 32512 15902 32524
rect 18138 32512 18144 32524
rect 18196 32512 18202 32564
rect 24029 32555 24087 32561
rect 24029 32521 24041 32555
rect 24075 32521 24087 32555
rect 25494 32555 25552 32561
rect 25494 32552 25506 32555
rect 24029 32515 24087 32521
rect 24504 32524 25506 32552
rect 1670 32444 1676 32496
rect 1728 32484 1734 32496
rect 1857 32487 1915 32493
rect 1857 32484 1869 32487
rect 1728 32456 1869 32484
rect 1728 32444 1734 32456
rect 1857 32453 1869 32456
rect 1903 32453 1915 32487
rect 1857 32447 1915 32453
rect 2590 32444 2596 32496
rect 2648 32444 2654 32496
rect 3602 32444 3608 32496
rect 3660 32444 3666 32496
rect 6546 32493 6552 32496
rect 6517 32487 6552 32493
rect 6517 32484 6529 32487
rect 5644 32456 6529 32484
rect 5644 32428 5672 32456
rect 6517 32453 6529 32456
rect 6517 32447 6552 32453
rect 6546 32444 6552 32447
rect 6604 32444 6610 32496
rect 6638 32444 6644 32496
rect 6696 32484 6702 32496
rect 6733 32487 6791 32493
rect 6733 32484 6745 32487
rect 6696 32456 6745 32484
rect 6696 32444 6702 32456
rect 6733 32453 6745 32456
rect 6779 32453 6791 32487
rect 6733 32447 6791 32453
rect 6914 32444 6920 32496
rect 6972 32484 6978 32496
rect 7745 32487 7803 32493
rect 7745 32484 7757 32487
rect 6972 32456 7757 32484
rect 6972 32444 6978 32456
rect 7745 32453 7757 32456
rect 7791 32484 7803 32487
rect 8757 32487 8815 32493
rect 8757 32484 8769 32487
rect 7791 32456 8769 32484
rect 7791 32453 7803 32456
rect 7745 32447 7803 32453
rect 8757 32453 8769 32456
rect 8803 32453 8815 32487
rect 8757 32447 8815 32453
rect 8846 32444 8852 32496
rect 8904 32484 8910 32496
rect 8904 32456 13768 32484
rect 8904 32444 8910 32456
rect 5169 32419 5227 32425
rect 5169 32385 5181 32419
rect 5215 32385 5227 32419
rect 5169 32379 5227 32385
rect 5445 32419 5503 32425
rect 5445 32385 5457 32419
rect 5491 32416 5503 32419
rect 5626 32416 5632 32428
rect 5491 32388 5632 32416
rect 5491 32385 5503 32388
rect 5445 32379 5503 32385
rect 3878 32308 3884 32360
rect 3936 32308 3942 32360
rect 5184 32348 5212 32379
rect 5626 32376 5632 32388
rect 5684 32376 5690 32428
rect 5721 32419 5779 32425
rect 5721 32385 5733 32419
rect 5767 32416 5779 32419
rect 6178 32416 6184 32428
rect 5767 32388 6184 32416
rect 5767 32385 5779 32388
rect 5721 32379 5779 32385
rect 6178 32376 6184 32388
rect 6236 32416 6242 32428
rect 7190 32416 7196 32428
rect 6236 32388 7196 32416
rect 6236 32376 6242 32388
rect 7190 32376 7196 32388
rect 7248 32376 7254 32428
rect 7466 32425 7472 32428
rect 7436 32419 7472 32425
rect 7436 32385 7448 32419
rect 7436 32379 7472 32385
rect 7466 32376 7472 32379
rect 7524 32376 7530 32428
rect 8570 32376 8576 32428
rect 8628 32376 8634 32428
rect 11606 32376 11612 32428
rect 11664 32416 11670 32428
rect 12253 32419 12311 32425
rect 12253 32416 12265 32419
rect 11664 32388 12265 32416
rect 11664 32376 11670 32388
rect 12253 32385 12265 32388
rect 12299 32385 12311 32419
rect 13078 32416 13084 32428
rect 12253 32379 12311 32385
rect 12452 32388 13084 32416
rect 5534 32348 5540 32360
rect 5184 32320 5540 32348
rect 5534 32308 5540 32320
rect 5592 32308 5598 32360
rect 5810 32308 5816 32360
rect 5868 32308 5874 32360
rect 6914 32308 6920 32360
rect 6972 32308 6978 32360
rect 7009 32351 7067 32357
rect 7009 32317 7021 32351
rect 7055 32348 7067 32351
rect 9214 32348 9220 32360
rect 7055 32320 9220 32348
rect 7055 32317 7067 32320
rect 7009 32311 7067 32317
rect 9214 32308 9220 32320
rect 9272 32308 9278 32360
rect 10962 32308 10968 32360
rect 11020 32348 11026 32360
rect 11517 32351 11575 32357
rect 11517 32348 11529 32351
rect 11020 32320 11529 32348
rect 11020 32308 11026 32320
rect 11517 32317 11529 32320
rect 11563 32317 11575 32351
rect 11517 32311 11575 32317
rect 11882 32308 11888 32360
rect 11940 32348 11946 32360
rect 12452 32348 12480 32388
rect 13078 32376 13084 32388
rect 13136 32376 13142 32428
rect 13740 32416 13768 32456
rect 14568 32456 16068 32484
rect 13906 32416 13912 32428
rect 13740 32388 13912 32416
rect 13906 32376 13912 32388
rect 13964 32376 13970 32428
rect 14182 32376 14188 32428
rect 14240 32376 14246 32428
rect 11940 32320 12480 32348
rect 11940 32308 11946 32320
rect 12526 32308 12532 32360
rect 12584 32308 12590 32360
rect 12618 32308 12624 32360
rect 12676 32348 12682 32360
rect 13265 32351 13323 32357
rect 13265 32348 13277 32351
rect 12676 32320 13277 32348
rect 12676 32308 12682 32320
rect 13265 32317 13277 32320
rect 13311 32317 13323 32351
rect 13265 32311 13323 32317
rect 13814 32308 13820 32360
rect 13872 32348 13878 32360
rect 14461 32351 14519 32357
rect 14461 32348 14473 32351
rect 13872 32320 14473 32348
rect 13872 32308 13878 32320
rect 14461 32317 14473 32320
rect 14507 32317 14519 32351
rect 14461 32311 14519 32317
rect 3896 32280 3924 32308
rect 5902 32280 5908 32292
rect 3896 32252 5908 32280
rect 5902 32240 5908 32252
rect 5960 32240 5966 32292
rect 6362 32240 6368 32292
rect 6420 32240 6426 32292
rect 11977 32283 12035 32289
rect 11977 32249 11989 32283
rect 12023 32249 12035 32283
rect 11977 32243 12035 32249
rect 5169 32215 5227 32221
rect 5169 32181 5181 32215
rect 5215 32212 5227 32215
rect 5994 32212 6000 32224
rect 5215 32184 6000 32212
rect 5215 32181 5227 32184
rect 5169 32175 5227 32181
rect 5994 32172 6000 32184
rect 6052 32172 6058 32224
rect 6270 32172 6276 32224
rect 6328 32212 6334 32224
rect 6546 32212 6552 32224
rect 6328 32184 6552 32212
rect 6328 32172 6334 32184
rect 6546 32172 6552 32184
rect 6604 32172 6610 32224
rect 11992 32212 12020 32243
rect 12066 32240 12072 32292
rect 12124 32280 12130 32292
rect 12124 32252 12572 32280
rect 12124 32240 12130 32252
rect 12434 32212 12440 32224
rect 11992 32184 12440 32212
rect 12434 32172 12440 32184
rect 12492 32172 12498 32224
rect 12544 32212 12572 32252
rect 12986 32240 12992 32292
rect 13044 32280 13050 32292
rect 14568 32280 14596 32456
rect 14642 32376 14648 32428
rect 14700 32416 14706 32428
rect 14829 32419 14887 32425
rect 14829 32416 14841 32419
rect 14700 32388 14841 32416
rect 14700 32376 14706 32388
rect 14829 32385 14841 32388
rect 14875 32385 14887 32419
rect 16040 32416 16068 32456
rect 16114 32444 16120 32496
rect 16172 32484 16178 32496
rect 18230 32484 18236 32496
rect 16172 32456 18236 32484
rect 16172 32444 16178 32456
rect 18230 32444 18236 32456
rect 18288 32444 18294 32496
rect 20346 32444 20352 32496
rect 20404 32484 20410 32496
rect 21450 32484 21456 32496
rect 20404 32456 21456 32484
rect 20404 32444 20410 32456
rect 21450 32444 21456 32456
rect 21508 32484 21514 32496
rect 24044 32484 24072 32515
rect 21508 32456 22324 32484
rect 21508 32444 21514 32456
rect 17034 32416 17040 32428
rect 16040 32388 17040 32416
rect 14829 32379 14887 32385
rect 17034 32376 17040 32388
rect 17092 32376 17098 32428
rect 20257 32419 20315 32425
rect 20257 32385 20269 32419
rect 20303 32416 20315 32419
rect 20898 32416 20904 32428
rect 20303 32388 20904 32416
rect 20303 32385 20315 32388
rect 20257 32379 20315 32385
rect 20898 32376 20904 32388
rect 20956 32376 20962 32428
rect 22005 32419 22063 32425
rect 22005 32385 22017 32419
rect 22051 32416 22063 32419
rect 22186 32416 22192 32428
rect 22051 32388 22192 32416
rect 22051 32385 22063 32388
rect 22005 32379 22063 32385
rect 22186 32376 22192 32388
rect 22244 32376 22250 32428
rect 22296 32425 22324 32456
rect 22480 32456 24072 32484
rect 22480 32425 22508 32456
rect 22281 32419 22339 32425
rect 22281 32385 22293 32419
rect 22327 32385 22339 32419
rect 22281 32379 22339 32385
rect 22465 32419 22523 32425
rect 22465 32385 22477 32419
rect 22511 32385 22523 32419
rect 22465 32379 22523 32385
rect 14734 32308 14740 32360
rect 14792 32308 14798 32360
rect 15378 32308 15384 32360
rect 15436 32348 15442 32360
rect 16206 32348 16212 32360
rect 15436 32320 16212 32348
rect 15436 32308 15442 32320
rect 16206 32308 16212 32320
rect 16264 32308 16270 32360
rect 19426 32308 19432 32360
rect 19484 32348 19490 32360
rect 20165 32351 20223 32357
rect 20165 32348 20177 32351
rect 19484 32320 20177 32348
rect 19484 32308 19490 32320
rect 20165 32317 20177 32320
rect 20211 32317 20223 32351
rect 20165 32311 20223 32317
rect 20346 32308 20352 32360
rect 20404 32308 20410 32360
rect 20441 32351 20499 32357
rect 20441 32317 20453 32351
rect 20487 32348 20499 32351
rect 22097 32351 22155 32357
rect 22097 32348 22109 32351
rect 20487 32320 22109 32348
rect 20487 32317 20499 32320
rect 20441 32311 20499 32317
rect 13044 32252 14596 32280
rect 14645 32283 14703 32289
rect 13044 32240 13050 32252
rect 14645 32249 14657 32283
rect 14691 32280 14703 32283
rect 15194 32280 15200 32292
rect 14691 32252 15200 32280
rect 14691 32249 14703 32252
rect 14645 32243 14703 32249
rect 15194 32240 15200 32252
rect 15252 32240 15258 32292
rect 14550 32212 14556 32224
rect 12544 32184 14556 32212
rect 14550 32172 14556 32184
rect 14608 32172 14614 32224
rect 20346 32172 20352 32224
rect 20404 32212 20410 32224
rect 20625 32215 20683 32221
rect 20625 32212 20637 32215
rect 20404 32184 20637 32212
rect 20404 32172 20410 32184
rect 20625 32181 20637 32184
rect 20671 32181 20683 32215
rect 20625 32175 20683 32181
rect 21818 32172 21824 32224
rect 21876 32172 21882 32224
rect 22020 32212 22048 32320
rect 22097 32317 22109 32320
rect 22143 32317 22155 32351
rect 22296 32348 22324 32379
rect 22738 32376 22744 32428
rect 22796 32376 22802 32428
rect 22833 32419 22891 32425
rect 22833 32385 22845 32419
rect 22879 32385 22891 32419
rect 22833 32379 22891 32385
rect 22925 32419 22983 32425
rect 22925 32385 22937 32419
rect 22971 32416 22983 32419
rect 23014 32416 23020 32428
rect 22971 32388 23020 32416
rect 22971 32385 22983 32388
rect 22925 32379 22983 32385
rect 22646 32348 22652 32360
rect 22296 32320 22652 32348
rect 22097 32311 22155 32317
rect 22646 32308 22652 32320
rect 22704 32308 22710 32360
rect 22848 32348 22876 32379
rect 23014 32376 23020 32388
rect 23072 32376 23078 32428
rect 23109 32419 23167 32425
rect 23109 32385 23121 32419
rect 23155 32416 23167 32419
rect 23290 32416 23296 32428
rect 23155 32388 23296 32416
rect 23155 32385 23167 32388
rect 23109 32379 23167 32385
rect 23290 32376 23296 32388
rect 23348 32376 23354 32428
rect 23382 32376 23388 32428
rect 23440 32376 23446 32428
rect 23750 32376 23756 32428
rect 23808 32416 23814 32428
rect 24213 32419 24271 32425
rect 24213 32416 24225 32419
rect 23808 32388 24225 32416
rect 23808 32376 23814 32388
rect 24213 32385 24225 32388
rect 24259 32385 24271 32419
rect 24213 32379 24271 32385
rect 24397 32419 24455 32425
rect 24397 32385 24409 32419
rect 24443 32416 24455 32419
rect 24504 32416 24532 32524
rect 25494 32521 25506 32524
rect 25540 32552 25552 32555
rect 25682 32552 25688 32564
rect 25540 32524 25688 32552
rect 25540 32521 25552 32524
rect 25494 32515 25552 32521
rect 25682 32512 25688 32524
rect 25740 32512 25746 32564
rect 25774 32512 25780 32564
rect 25832 32552 25838 32564
rect 28902 32552 28908 32564
rect 25832 32524 26648 32552
rect 25832 32512 25838 32524
rect 24670 32444 24676 32496
rect 24728 32444 24734 32496
rect 25130 32444 25136 32496
rect 25188 32484 25194 32496
rect 25188 32456 25820 32484
rect 25188 32444 25194 32456
rect 24443 32388 24532 32416
rect 24443 32385 24455 32388
rect 24397 32379 24455 32385
rect 24854 32376 24860 32428
rect 24912 32376 24918 32428
rect 24946 32376 24952 32428
rect 25004 32376 25010 32428
rect 25038 32376 25044 32428
rect 25096 32425 25102 32428
rect 25096 32416 25104 32425
rect 25096 32388 25141 32416
rect 25096 32379 25104 32388
rect 25096 32376 25102 32379
rect 25314 32376 25320 32428
rect 25372 32376 25378 32428
rect 25406 32376 25412 32428
rect 25464 32376 25470 32428
rect 25590 32376 25596 32428
rect 25648 32376 25654 32428
rect 25792 32425 25820 32456
rect 26418 32444 26424 32496
rect 26476 32444 26482 32496
rect 26620 32493 26648 32524
rect 28184 32524 28908 32552
rect 26605 32487 26663 32493
rect 26605 32453 26617 32487
rect 26651 32453 26663 32487
rect 26605 32447 26663 32453
rect 28074 32444 28080 32496
rect 28132 32484 28138 32496
rect 28184 32493 28212 32524
rect 28902 32512 28908 32524
rect 28960 32512 28966 32564
rect 28994 32512 29000 32564
rect 29052 32552 29058 32564
rect 29730 32552 29736 32564
rect 29052 32524 29736 32552
rect 29052 32512 29058 32524
rect 29730 32512 29736 32524
rect 29788 32512 29794 32564
rect 29914 32512 29920 32564
rect 29972 32512 29978 32564
rect 31849 32555 31907 32561
rect 31849 32521 31861 32555
rect 31895 32552 31907 32555
rect 31938 32552 31944 32564
rect 31895 32524 31944 32552
rect 31895 32521 31907 32524
rect 31849 32515 31907 32521
rect 31938 32512 31944 32524
rect 31996 32512 32002 32564
rect 34330 32552 34336 32564
rect 34256 32524 34336 32552
rect 28169 32487 28227 32493
rect 28169 32484 28181 32487
rect 28132 32456 28181 32484
rect 28132 32444 28138 32456
rect 28169 32453 28181 32456
rect 28215 32453 28227 32487
rect 28169 32447 28227 32453
rect 28353 32487 28411 32493
rect 28353 32453 28365 32487
rect 28399 32484 28411 32487
rect 28399 32456 29040 32484
rect 28399 32453 28411 32456
rect 28353 32447 28411 32453
rect 25777 32419 25835 32425
rect 25777 32385 25789 32419
rect 25823 32385 25835 32419
rect 25777 32379 25835 32385
rect 25961 32419 26019 32425
rect 25961 32385 25973 32419
rect 26007 32385 26019 32419
rect 25961 32379 26019 32385
rect 23400 32348 23428 32376
rect 22848 32320 23428 32348
rect 23661 32351 23719 32357
rect 23661 32317 23673 32351
rect 23707 32348 23719 32351
rect 23842 32348 23848 32360
rect 23707 32320 23848 32348
rect 23707 32317 23719 32320
rect 23661 32311 23719 32317
rect 22189 32283 22247 32289
rect 22189 32249 22201 32283
rect 22235 32280 22247 32283
rect 23201 32283 23259 32289
rect 23201 32280 23213 32283
rect 22235 32252 23213 32280
rect 22235 32249 22247 32252
rect 22189 32243 22247 32249
rect 23201 32249 23213 32252
rect 23247 32249 23259 32283
rect 23676 32280 23704 32311
rect 23842 32308 23848 32320
rect 23900 32308 23906 32360
rect 24305 32351 24363 32357
rect 24305 32317 24317 32351
rect 24351 32317 24363 32351
rect 24305 32311 24363 32317
rect 23201 32243 23259 32249
rect 23308 32252 23704 32280
rect 24320 32280 24348 32311
rect 24486 32308 24492 32360
rect 24544 32308 24550 32360
rect 24765 32351 24823 32357
rect 24765 32317 24777 32351
rect 24811 32348 24823 32351
rect 25976 32348 26004 32379
rect 26050 32376 26056 32428
rect 26108 32376 26114 32428
rect 26237 32419 26295 32425
rect 26237 32385 26249 32419
rect 26283 32385 26295 32419
rect 26237 32379 26295 32385
rect 24811 32320 26004 32348
rect 26252 32348 26280 32379
rect 26326 32376 26332 32428
rect 26384 32376 26390 32428
rect 27890 32376 27896 32428
rect 27948 32416 27954 32428
rect 27948 32388 28764 32416
rect 27948 32376 27954 32388
rect 26694 32348 26700 32360
rect 26252 32320 26700 32348
rect 24811 32317 24823 32320
rect 24765 32311 24823 32317
rect 26694 32308 26700 32320
rect 26752 32308 26758 32360
rect 28442 32308 28448 32360
rect 28500 32308 28506 32360
rect 28736 32348 28764 32388
rect 28810 32376 28816 32428
rect 28868 32376 28874 32428
rect 29012 32425 29040 32456
rect 30190 32444 30196 32496
rect 30248 32484 30254 32496
rect 30285 32487 30343 32493
rect 30285 32484 30297 32487
rect 30248 32456 30297 32484
rect 30248 32444 30254 32456
rect 30285 32453 30297 32456
rect 30331 32453 30343 32487
rect 30285 32447 30343 32453
rect 31110 32444 31116 32496
rect 31168 32484 31174 32496
rect 32861 32487 32919 32493
rect 32861 32484 32873 32487
rect 31168 32456 32873 32484
rect 31168 32444 31174 32456
rect 32861 32453 32873 32456
rect 32907 32453 32919 32487
rect 32861 32447 32919 32453
rect 33042 32444 33048 32496
rect 33100 32484 33106 32496
rect 33686 32484 33692 32496
rect 33100 32456 33692 32484
rect 33100 32444 33106 32456
rect 33686 32444 33692 32456
rect 33744 32444 33750 32496
rect 34256 32493 34284 32524
rect 34330 32512 34336 32524
rect 34388 32512 34394 32564
rect 34517 32555 34575 32561
rect 34517 32521 34529 32555
rect 34563 32552 34575 32555
rect 36446 32552 36452 32564
rect 34563 32524 36452 32552
rect 34563 32521 34575 32524
rect 34517 32515 34575 32521
rect 36446 32512 36452 32524
rect 36504 32512 36510 32564
rect 34241 32487 34299 32493
rect 34241 32453 34253 32487
rect 34287 32453 34299 32487
rect 34241 32447 34299 32453
rect 34606 32444 34612 32496
rect 34664 32484 34670 32496
rect 34664 32456 34914 32484
rect 34664 32444 34670 32456
rect 28997 32419 29055 32425
rect 28997 32385 29009 32419
rect 29043 32416 29055 32419
rect 29086 32416 29092 32428
rect 29043 32388 29092 32416
rect 29043 32385 29055 32388
rect 28997 32379 29055 32385
rect 29086 32376 29092 32388
rect 29144 32376 29150 32428
rect 29976 32419 30034 32425
rect 29976 32385 29988 32419
rect 30022 32416 30034 32419
rect 31205 32419 31263 32425
rect 31205 32416 31217 32419
rect 30022 32388 31217 32416
rect 30022 32385 30034 32388
rect 29976 32379 30034 32385
rect 31205 32385 31217 32388
rect 31251 32416 31263 32419
rect 31386 32416 31392 32428
rect 31251 32388 31392 32416
rect 31251 32385 31263 32388
rect 31205 32379 31263 32385
rect 31386 32376 31392 32388
rect 31444 32376 31450 32428
rect 31478 32376 31484 32428
rect 31536 32416 31542 32428
rect 31665 32419 31723 32425
rect 31665 32416 31677 32419
rect 31536 32388 31677 32416
rect 31536 32376 31542 32388
rect 31665 32385 31677 32388
rect 31711 32385 31723 32419
rect 32398 32416 32404 32428
rect 31665 32379 31723 32385
rect 31772 32388 32404 32416
rect 29362 32348 29368 32360
rect 28736 32320 29368 32348
rect 29362 32308 29368 32320
rect 29420 32308 29426 32360
rect 29457 32351 29515 32357
rect 29457 32317 29469 32351
rect 29503 32348 29515 32351
rect 29730 32348 29736 32360
rect 29503 32320 29736 32348
rect 29503 32317 29515 32320
rect 29457 32311 29515 32317
rect 29730 32308 29736 32320
rect 29788 32308 29794 32360
rect 31573 32351 31631 32357
rect 31573 32317 31585 32351
rect 31619 32348 31631 32351
rect 31772 32348 31800 32388
rect 32398 32376 32404 32388
rect 32456 32376 32462 32428
rect 33962 32376 33968 32428
rect 34020 32376 34026 32428
rect 34146 32376 34152 32428
rect 34204 32376 34210 32428
rect 34333 32419 34391 32425
rect 34333 32385 34345 32419
rect 34379 32385 34391 32419
rect 34333 32379 34391 32385
rect 36357 32419 36415 32425
rect 36357 32385 36369 32419
rect 36403 32416 36415 32419
rect 37274 32416 37280 32428
rect 36403 32388 37280 32416
rect 36403 32385 36415 32388
rect 36357 32379 36415 32385
rect 31619 32320 31800 32348
rect 32677 32351 32735 32357
rect 31619 32317 31631 32320
rect 31573 32311 31631 32317
rect 32677 32317 32689 32351
rect 32723 32317 32735 32351
rect 34348 32348 34376 32379
rect 37274 32376 37280 32388
rect 37332 32416 37338 32428
rect 38194 32416 38200 32428
rect 37332 32388 38200 32416
rect 37332 32376 37338 32388
rect 38194 32376 38200 32388
rect 38252 32376 38258 32428
rect 34422 32348 34428 32360
rect 34348 32320 34428 32348
rect 32677 32311 32735 32317
rect 26789 32283 26847 32289
rect 26789 32280 26801 32283
rect 24320 32252 26801 32280
rect 22557 32215 22615 32221
rect 22557 32212 22569 32215
rect 22020 32184 22569 32212
rect 22557 32181 22569 32184
rect 22603 32181 22615 32215
rect 22557 32175 22615 32181
rect 22738 32172 22744 32224
rect 22796 32212 22802 32224
rect 23308 32212 23336 32252
rect 26789 32249 26801 32252
rect 26835 32249 26847 32283
rect 26789 32243 26847 32249
rect 28534 32240 28540 32292
rect 28592 32280 28598 32292
rect 29549 32283 29607 32289
rect 29549 32280 29561 32283
rect 28592 32252 29561 32280
rect 28592 32240 28598 32252
rect 29549 32249 29561 32252
rect 29595 32280 29607 32283
rect 30006 32280 30012 32292
rect 29595 32252 30012 32280
rect 29595 32249 29607 32252
rect 29549 32243 29607 32249
rect 30006 32240 30012 32252
rect 30064 32240 30070 32292
rect 30098 32240 30104 32292
rect 30156 32240 30162 32292
rect 31662 32280 31668 32292
rect 31588 32252 31668 32280
rect 22796 32184 23336 32212
rect 23569 32215 23627 32221
rect 22796 32172 22802 32184
rect 23569 32181 23581 32215
rect 23615 32212 23627 32215
rect 24210 32212 24216 32224
rect 23615 32184 24216 32212
rect 23615 32181 23627 32184
rect 23569 32175 23627 32181
rect 24210 32172 24216 32184
rect 24268 32172 24274 32224
rect 25314 32172 25320 32224
rect 25372 32212 25378 32224
rect 26142 32212 26148 32224
rect 25372 32184 26148 32212
rect 25372 32172 25378 32184
rect 26142 32172 26148 32184
rect 26200 32172 26206 32224
rect 27985 32215 28043 32221
rect 27985 32181 27997 32215
rect 28031 32212 28043 32215
rect 28074 32212 28080 32224
rect 28031 32184 28080 32212
rect 28031 32181 28043 32184
rect 27985 32175 28043 32181
rect 28074 32172 28080 32184
rect 28132 32172 28138 32224
rect 31588 32221 31616 32252
rect 31662 32240 31668 32252
rect 31720 32280 31726 32292
rect 32692 32280 32720 32311
rect 34422 32308 34428 32320
rect 34480 32348 34486 32360
rect 35986 32348 35992 32360
rect 34480 32320 35992 32348
rect 34480 32308 34486 32320
rect 35986 32308 35992 32320
rect 36044 32308 36050 32360
rect 36078 32308 36084 32360
rect 36136 32308 36142 32360
rect 37458 32308 37464 32360
rect 37516 32308 37522 32360
rect 37550 32308 37556 32360
rect 37608 32308 37614 32360
rect 37645 32351 37703 32357
rect 37645 32317 37657 32351
rect 37691 32317 37703 32351
rect 37645 32311 37703 32317
rect 37737 32351 37795 32357
rect 37737 32317 37749 32351
rect 37783 32348 37795 32351
rect 37826 32348 37832 32360
rect 37783 32320 37832 32348
rect 37783 32317 37795 32320
rect 37737 32311 37795 32317
rect 31720 32252 32720 32280
rect 31720 32240 31726 32252
rect 37366 32240 37372 32292
rect 37424 32280 37430 32292
rect 37660 32280 37688 32311
rect 37826 32308 37832 32320
rect 37884 32308 37890 32360
rect 37424 32252 37688 32280
rect 37424 32240 37430 32252
rect 31573 32215 31631 32221
rect 31573 32181 31585 32215
rect 31619 32181 31631 32215
rect 31573 32175 31631 32181
rect 31846 32172 31852 32224
rect 31904 32212 31910 32224
rect 32125 32215 32183 32221
rect 32125 32212 32137 32215
rect 31904 32184 32137 32212
rect 31904 32172 31910 32184
rect 32125 32181 32137 32184
rect 32171 32181 32183 32215
rect 32125 32175 32183 32181
rect 34609 32215 34667 32221
rect 34609 32181 34621 32215
rect 34655 32212 34667 32215
rect 34790 32212 34796 32224
rect 34655 32184 34796 32212
rect 34655 32181 34667 32184
rect 34609 32175 34667 32181
rect 34790 32172 34796 32184
rect 34848 32172 34854 32224
rect 37277 32215 37335 32221
rect 37277 32181 37289 32215
rect 37323 32212 37335 32215
rect 38010 32212 38016 32224
rect 37323 32184 38016 32212
rect 37323 32181 37335 32184
rect 37277 32175 37335 32181
rect 38010 32172 38016 32184
rect 38068 32172 38074 32224
rect 1104 32122 40572 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 40572 32122
rect 1104 32048 40572 32070
rect 2590 31968 2596 32020
rect 2648 32008 2654 32020
rect 4525 32011 4583 32017
rect 4525 32008 4537 32011
rect 2648 31980 4537 32008
rect 2648 31968 2654 31980
rect 4525 31977 4537 31980
rect 4571 31977 4583 32011
rect 4525 31971 4583 31977
rect 5718 31968 5724 32020
rect 5776 32008 5782 32020
rect 6270 32008 6276 32020
rect 5776 31980 6276 32008
rect 5776 31968 5782 31980
rect 6270 31968 6276 31980
rect 6328 31968 6334 32020
rect 7374 31968 7380 32020
rect 7432 32008 7438 32020
rect 7837 32011 7895 32017
rect 7837 32008 7849 32011
rect 7432 31980 7849 32008
rect 7432 31968 7438 31980
rect 7837 31977 7849 31980
rect 7883 31977 7895 32011
rect 7837 31971 7895 31977
rect 8573 32011 8631 32017
rect 8573 31977 8585 32011
rect 8619 32008 8631 32011
rect 8662 32008 8668 32020
rect 8619 31980 8668 32008
rect 8619 31977 8631 31980
rect 8573 31971 8631 31977
rect 8662 31968 8668 31980
rect 8720 31968 8726 32020
rect 9030 31968 9036 32020
rect 9088 31968 9094 32020
rect 10962 31968 10968 32020
rect 11020 31968 11026 32020
rect 11054 31968 11060 32020
rect 11112 31968 11118 32020
rect 11698 31968 11704 32020
rect 11756 32008 11762 32020
rect 11756 31980 14261 32008
rect 11756 31968 11762 31980
rect 5534 31900 5540 31952
rect 5592 31940 5598 31952
rect 6638 31940 6644 31952
rect 5592 31912 6644 31940
rect 5592 31900 5598 31912
rect 6638 31900 6644 31912
rect 6696 31900 6702 31952
rect 9048 31940 9076 31968
rect 12526 31940 12532 31952
rect 6748 31912 9076 31940
rect 12176 31912 12532 31940
rect 5810 31832 5816 31884
rect 5868 31872 5874 31884
rect 6086 31872 6092 31884
rect 5868 31844 6092 31872
rect 5868 31832 5874 31844
rect 6086 31832 6092 31844
rect 6144 31872 6150 31884
rect 6748 31872 6776 31912
rect 6144 31844 6776 31872
rect 6144 31832 6150 31844
rect 8018 31832 8024 31884
rect 8076 31832 8082 31884
rect 10413 31875 10471 31881
rect 8772 31844 9168 31872
rect 3786 31764 3792 31816
rect 3844 31804 3850 31816
rect 4801 31807 4859 31813
rect 4801 31804 4813 31807
rect 3844 31776 4813 31804
rect 3844 31764 3850 31776
rect 4801 31773 4813 31776
rect 4847 31773 4859 31807
rect 4801 31767 4859 31773
rect 5721 31807 5779 31813
rect 5721 31773 5733 31807
rect 5767 31804 5779 31807
rect 5902 31804 5908 31816
rect 5767 31776 5908 31804
rect 5767 31773 5779 31776
rect 5721 31767 5779 31773
rect 5902 31764 5908 31776
rect 5960 31764 5966 31816
rect 8113 31807 8171 31813
rect 8113 31773 8125 31807
rect 8159 31773 8171 31807
rect 8113 31767 8171 31773
rect 5258 31696 5264 31748
rect 5316 31736 5322 31748
rect 7834 31736 7840 31748
rect 5316 31708 7840 31736
rect 5316 31696 5322 31708
rect 7834 31696 7840 31708
rect 7892 31736 7898 31748
rect 8128 31736 8156 31767
rect 8772 31748 8800 31844
rect 9140 31813 9168 31844
rect 10413 31841 10425 31875
rect 10459 31872 10471 31875
rect 11609 31875 11667 31881
rect 11609 31872 11621 31875
rect 10459 31844 11621 31872
rect 10459 31841 10471 31844
rect 10413 31835 10471 31841
rect 11609 31841 11621 31844
rect 11655 31872 11667 31875
rect 11882 31872 11888 31884
rect 11655 31844 11888 31872
rect 11655 31841 11667 31844
rect 11609 31835 11667 31841
rect 11882 31832 11888 31844
rect 11940 31832 11946 31884
rect 12069 31875 12127 31881
rect 12069 31841 12081 31875
rect 12115 31872 12127 31875
rect 12176 31872 12204 31912
rect 12526 31900 12532 31912
rect 12584 31900 12590 31952
rect 14093 31943 14151 31949
rect 14093 31940 14105 31943
rect 13648 31912 14105 31940
rect 12115 31844 12204 31872
rect 12115 31841 12127 31844
rect 12069 31835 12127 31841
rect 12250 31832 12256 31884
rect 12308 31872 12314 31884
rect 12897 31875 12955 31881
rect 12897 31872 12909 31875
rect 12308 31844 12909 31872
rect 12308 31832 12314 31844
rect 12897 31841 12909 31844
rect 12943 31841 12955 31875
rect 12897 31835 12955 31841
rect 9125 31807 9183 31813
rect 9125 31773 9137 31807
rect 9171 31773 9183 31807
rect 9125 31767 9183 31773
rect 11238 31764 11244 31816
rect 11296 31804 11302 31816
rect 11517 31807 11575 31813
rect 11517 31804 11529 31807
rect 11296 31776 11529 31804
rect 11296 31764 11302 31776
rect 11517 31773 11529 31776
rect 11563 31773 11575 31807
rect 11517 31767 11575 31773
rect 12158 31764 12164 31816
rect 12216 31764 12222 31816
rect 12528 31807 12586 31813
rect 12528 31773 12540 31807
rect 12574 31804 12586 31807
rect 12710 31804 12716 31816
rect 12574 31776 12716 31804
rect 12574 31773 12586 31776
rect 12528 31767 12586 31773
rect 12710 31764 12716 31776
rect 12768 31764 12774 31816
rect 13357 31807 13415 31813
rect 13357 31773 13369 31807
rect 13403 31804 13415 31807
rect 13648 31804 13676 31912
rect 14093 31909 14105 31912
rect 14139 31909 14151 31943
rect 14093 31903 14151 31909
rect 13832 31844 14044 31872
rect 13403 31776 13676 31804
rect 13403 31773 13415 31776
rect 13357 31767 13415 31773
rect 13722 31764 13728 31816
rect 13780 31764 13786 31816
rect 7892 31708 8156 31736
rect 7892 31696 7898 31708
rect 8202 31696 8208 31748
rect 8260 31736 8266 31748
rect 8260 31708 8600 31736
rect 8260 31696 8266 31708
rect 8294 31628 8300 31680
rect 8352 31668 8358 31680
rect 8572 31677 8600 31708
rect 8754 31696 8760 31748
rect 8812 31696 8818 31748
rect 8938 31696 8944 31748
rect 8996 31736 9002 31748
rect 11146 31736 11152 31748
rect 8996 31708 11152 31736
rect 8996 31696 9002 31708
rect 11146 31696 11152 31708
rect 11204 31696 11210 31748
rect 11422 31696 11428 31748
rect 11480 31736 11486 31748
rect 13832 31736 13860 31844
rect 13906 31764 13912 31816
rect 13964 31764 13970 31816
rect 11480 31708 13860 31736
rect 14016 31736 14044 31844
rect 14233 31813 14261 31980
rect 14550 31968 14556 32020
rect 14608 32008 14614 32020
rect 14645 32011 14703 32017
rect 14645 32008 14657 32011
rect 14608 31980 14657 32008
rect 14608 31968 14614 31980
rect 14645 31977 14657 31980
rect 14691 32008 14703 32011
rect 14918 32008 14924 32020
rect 14691 31980 14924 32008
rect 14691 31977 14703 31980
rect 14645 31971 14703 31977
rect 14918 31968 14924 31980
rect 14976 31968 14982 32020
rect 17218 31968 17224 32020
rect 17276 32008 17282 32020
rect 21082 32008 21088 32020
rect 17276 31980 21088 32008
rect 17276 31968 17282 31980
rect 14734 31832 14740 31884
rect 14792 31872 14798 31884
rect 15197 31875 15255 31881
rect 15197 31872 15209 31875
rect 14792 31844 15209 31872
rect 14792 31832 14798 31844
rect 15197 31841 15209 31844
rect 15243 31841 15255 31875
rect 15197 31835 15255 31841
rect 16114 31832 16120 31884
rect 16172 31832 16178 31884
rect 17218 31832 17224 31884
rect 17276 31832 17282 31884
rect 17497 31875 17555 31881
rect 17497 31841 17509 31875
rect 17543 31872 17555 31875
rect 18046 31872 18052 31884
rect 17543 31844 18052 31872
rect 17543 31841 17555 31844
rect 17497 31835 17555 31841
rect 18046 31832 18052 31844
rect 18104 31832 18110 31884
rect 19352 31881 19380 31980
rect 21082 31968 21088 31980
rect 21140 31968 21146 32020
rect 22554 31968 22560 32020
rect 22612 31968 22618 32020
rect 23014 31968 23020 32020
rect 23072 32008 23078 32020
rect 25314 32008 25320 32020
rect 23072 31980 25320 32008
rect 23072 31968 23078 31980
rect 25314 31968 25320 31980
rect 25372 31968 25378 32020
rect 26602 32008 26608 32020
rect 25884 31980 26608 32008
rect 25593 31943 25651 31949
rect 22388 31912 22968 31940
rect 19337 31875 19395 31881
rect 19337 31841 19349 31875
rect 19383 31841 19395 31875
rect 19337 31835 19395 31841
rect 20622 31832 20628 31884
rect 20680 31872 20686 31884
rect 21085 31875 21143 31881
rect 20680 31844 20944 31872
rect 20680 31832 20686 31844
rect 14218 31807 14276 31813
rect 14218 31773 14230 31807
rect 14264 31773 14276 31807
rect 14218 31767 14276 31773
rect 15286 31764 15292 31816
rect 15344 31764 15350 31816
rect 15470 31764 15476 31816
rect 15528 31804 15534 31816
rect 15933 31807 15991 31813
rect 15933 31804 15945 31807
rect 15528 31776 15945 31804
rect 15528 31764 15534 31776
rect 15933 31773 15945 31776
rect 15979 31773 15991 31807
rect 15933 31767 15991 31773
rect 16298 31764 16304 31816
rect 16356 31764 16362 31816
rect 16390 31764 16396 31816
rect 16448 31764 16454 31816
rect 18616 31776 19288 31804
rect 16758 31736 16764 31748
rect 14016 31708 16764 31736
rect 11480 31696 11486 31708
rect 16758 31696 16764 31708
rect 16816 31696 16822 31748
rect 17954 31736 17960 31748
rect 17880 31708 17960 31736
rect 8389 31671 8447 31677
rect 8389 31668 8401 31671
rect 8352 31640 8401 31668
rect 8352 31628 8358 31640
rect 8389 31637 8401 31640
rect 8435 31637 8447 31671
rect 8389 31631 8447 31637
rect 8557 31671 8615 31677
rect 8557 31637 8569 31671
rect 8603 31668 8615 31671
rect 9030 31668 9036 31680
rect 8603 31640 9036 31668
rect 8603 31637 8615 31640
rect 8557 31631 8615 31637
rect 9030 31628 9036 31640
rect 9088 31628 9094 31680
rect 10502 31628 10508 31680
rect 10560 31628 10566 31680
rect 10597 31671 10655 31677
rect 10597 31637 10609 31671
rect 10643 31668 10655 31671
rect 11882 31668 11888 31680
rect 10643 31640 11888 31668
rect 10643 31637 10655 31640
rect 10597 31631 10655 31637
rect 11882 31628 11888 31640
rect 11940 31628 11946 31680
rect 12621 31671 12679 31677
rect 12621 31637 12633 31671
rect 12667 31668 12679 31671
rect 12986 31668 12992 31680
rect 12667 31640 12992 31668
rect 12667 31637 12679 31640
rect 12621 31631 12679 31637
rect 12986 31628 12992 31640
rect 13044 31628 13050 31680
rect 13630 31628 13636 31680
rect 13688 31668 13694 31680
rect 14277 31671 14335 31677
rect 14277 31668 14289 31671
rect 13688 31640 14289 31668
rect 13688 31628 13694 31640
rect 14277 31637 14289 31640
rect 14323 31637 14335 31671
rect 17880 31668 17908 31708
rect 17954 31696 17960 31708
rect 18012 31696 18018 31748
rect 18506 31668 18512 31680
rect 17880 31640 18512 31668
rect 14277 31631 14335 31637
rect 18506 31628 18512 31640
rect 18564 31668 18570 31680
rect 18616 31668 18644 31776
rect 19260 31748 19288 31776
rect 19242 31696 19248 31748
rect 19300 31696 19306 31748
rect 19610 31696 19616 31748
rect 19668 31696 19674 31748
rect 20916 31736 20944 31844
rect 21085 31841 21097 31875
rect 21131 31872 21143 31875
rect 21729 31875 21787 31881
rect 21729 31872 21741 31875
rect 21131 31844 21741 31872
rect 21131 31841 21143 31844
rect 21085 31835 21143 31841
rect 21729 31841 21741 31844
rect 21775 31872 21787 31875
rect 22094 31872 22100 31884
rect 21775 31844 22100 31872
rect 21775 31841 21787 31844
rect 21729 31835 21787 31841
rect 22094 31832 22100 31844
rect 22152 31832 22158 31884
rect 22186 31764 22192 31816
rect 22244 31764 22250 31816
rect 21358 31736 21364 31748
rect 20838 31708 21364 31736
rect 21358 31696 21364 31708
rect 21416 31696 21422 31748
rect 18564 31640 18644 31668
rect 18969 31671 19027 31677
rect 18564 31628 18570 31640
rect 18969 31637 18981 31671
rect 19015 31668 19027 31671
rect 19058 31668 19064 31680
rect 19015 31640 19064 31668
rect 19015 31637 19027 31640
rect 18969 31631 19027 31637
rect 19058 31628 19064 31640
rect 19116 31628 19122 31680
rect 21174 31628 21180 31680
rect 21232 31628 21238 31680
rect 22186 31628 22192 31680
rect 22244 31668 22250 31680
rect 22388 31677 22416 31912
rect 22646 31832 22652 31884
rect 22704 31872 22710 31884
rect 22940 31881 22968 31912
rect 25593 31909 25605 31943
rect 25639 31940 25651 31943
rect 25774 31940 25780 31952
rect 25639 31912 25780 31940
rect 25639 31909 25651 31912
rect 25593 31903 25651 31909
rect 25774 31900 25780 31912
rect 25832 31900 25838 31952
rect 22833 31875 22891 31881
rect 22833 31872 22845 31875
rect 22704 31844 22845 31872
rect 22704 31832 22710 31844
rect 22833 31841 22845 31844
rect 22879 31841 22891 31875
rect 22833 31835 22891 31841
rect 22925 31875 22983 31881
rect 22925 31841 22937 31875
rect 22971 31841 22983 31875
rect 23750 31872 23756 31884
rect 22925 31835 22983 31841
rect 23436 31844 23756 31872
rect 22733 31807 22791 31813
rect 22733 31773 22745 31807
rect 22779 31804 22791 31807
rect 22779 31776 22876 31804
rect 22779 31773 22791 31776
rect 22733 31767 22791 31773
rect 22848 31680 22876 31776
rect 23014 31764 23020 31816
rect 23072 31764 23078 31816
rect 23436 31813 23464 31844
rect 23750 31832 23756 31844
rect 23808 31872 23814 31884
rect 24854 31872 24860 31884
rect 23808 31844 24860 31872
rect 23808 31832 23814 31844
rect 24854 31832 24860 31844
rect 24912 31832 24918 31884
rect 25041 31875 25099 31881
rect 25041 31841 25053 31875
rect 25087 31872 25099 31875
rect 25501 31875 25559 31881
rect 25501 31872 25513 31875
rect 25087 31844 25513 31872
rect 25087 31841 25099 31844
rect 25041 31835 25099 31841
rect 25501 31841 25513 31844
rect 25547 31841 25559 31875
rect 25501 31835 25559 31841
rect 23385 31807 23464 31813
rect 23385 31773 23397 31807
rect 23431 31778 23464 31807
rect 23569 31807 23627 31813
rect 23431 31773 23443 31778
rect 23385 31767 23443 31773
rect 23569 31773 23581 31807
rect 23615 31804 23627 31807
rect 23842 31804 23848 31816
rect 23615 31776 23848 31804
rect 23615 31773 23627 31776
rect 23569 31767 23627 31773
rect 23842 31764 23848 31776
rect 23900 31764 23906 31816
rect 24949 31807 25007 31813
rect 24949 31804 24961 31807
rect 23952 31776 24961 31804
rect 23753 31739 23811 31745
rect 23753 31705 23765 31739
rect 23799 31736 23811 31739
rect 23860 31736 23888 31764
rect 23952 31745 23980 31776
rect 24949 31773 24961 31776
rect 24995 31773 25007 31807
rect 24949 31767 25007 31773
rect 25222 31764 25228 31816
rect 25280 31764 25286 31816
rect 25409 31807 25467 31813
rect 25409 31773 25421 31807
rect 25455 31804 25467 31807
rect 25590 31804 25596 31816
rect 25455 31776 25596 31804
rect 25455 31773 25467 31776
rect 25409 31767 25467 31773
rect 25590 31764 25596 31776
rect 25648 31764 25654 31816
rect 25682 31764 25688 31816
rect 25740 31764 25746 31816
rect 25884 31813 25912 31980
rect 26602 31968 26608 31980
rect 26660 31968 26666 32020
rect 27890 32008 27896 32020
rect 27632 31980 27896 32008
rect 26418 31900 26424 31952
rect 26476 31900 26482 31952
rect 27433 31943 27491 31949
rect 27433 31909 27445 31943
rect 27479 31909 27491 31943
rect 27433 31903 27491 31909
rect 25961 31875 26019 31881
rect 25961 31841 25973 31875
rect 26007 31872 26019 31875
rect 26436 31872 26464 31900
rect 27338 31872 27344 31884
rect 26007 31844 26464 31872
rect 27172 31844 27344 31872
rect 26007 31841 26019 31844
rect 25961 31835 26019 31841
rect 25869 31807 25927 31813
rect 25869 31773 25881 31807
rect 25915 31773 25927 31807
rect 25869 31767 25927 31773
rect 26053 31807 26111 31813
rect 26053 31773 26065 31807
rect 26099 31773 26111 31807
rect 26053 31767 26111 31773
rect 23799 31708 23888 31736
rect 23937 31739 23995 31745
rect 23799 31705 23811 31708
rect 23753 31699 23811 31705
rect 23937 31705 23949 31739
rect 23983 31705 23995 31739
rect 23937 31699 23995 31705
rect 22373 31671 22431 31677
rect 22373 31668 22385 31671
rect 22244 31640 22385 31668
rect 22244 31628 22250 31640
rect 22373 31637 22385 31640
rect 22419 31637 22431 31671
rect 22373 31631 22431 31637
rect 22830 31628 22836 31680
rect 22888 31628 22894 31680
rect 23198 31628 23204 31680
rect 23256 31628 23262 31680
rect 23290 31628 23296 31680
rect 23348 31668 23354 31680
rect 23952 31668 23980 31699
rect 24118 31696 24124 31748
rect 24176 31696 24182 31748
rect 24578 31696 24584 31748
rect 24636 31736 24642 31748
rect 26068 31736 26096 31767
rect 26142 31764 26148 31816
rect 26200 31804 26206 31816
rect 26424 31807 26482 31813
rect 26424 31804 26436 31807
rect 26200 31776 26436 31804
rect 26200 31764 26206 31776
rect 26424 31773 26436 31776
rect 26470 31804 26482 31807
rect 27172 31804 27200 31844
rect 27338 31832 27344 31844
rect 27396 31832 27402 31884
rect 26470 31776 27200 31804
rect 26470 31773 26482 31776
rect 26424 31767 26482 31773
rect 27246 31764 27252 31816
rect 27304 31804 27310 31816
rect 27448 31804 27476 31903
rect 27632 31813 27660 31980
rect 27890 31968 27896 31980
rect 27948 31968 27954 32020
rect 29825 32011 29883 32017
rect 29825 32008 29837 32011
rect 28276 31980 29837 32008
rect 27709 31943 27767 31949
rect 27709 31909 27721 31943
rect 27755 31940 27767 31943
rect 27982 31940 27988 31952
rect 27755 31912 27988 31940
rect 27755 31909 27767 31912
rect 27709 31903 27767 31909
rect 27982 31900 27988 31912
rect 28040 31900 28046 31952
rect 28276 31940 28304 31980
rect 29825 31977 29837 31980
rect 29871 31977 29883 32011
rect 29825 31971 29883 31977
rect 30466 31968 30472 32020
rect 30524 32008 30530 32020
rect 30929 32011 30987 32017
rect 30929 32008 30941 32011
rect 30524 31980 30941 32008
rect 30524 31968 30530 31980
rect 30929 31977 30941 31980
rect 30975 31977 30987 32011
rect 30929 31971 30987 31977
rect 31662 31968 31668 32020
rect 31720 32008 31726 32020
rect 31720 31980 31800 32008
rect 31720 31968 31726 31980
rect 28092 31912 28304 31940
rect 28721 31943 28779 31949
rect 28092 31872 28120 31912
rect 28721 31909 28733 31943
rect 28767 31940 28779 31943
rect 28994 31940 29000 31952
rect 28767 31912 29000 31940
rect 28767 31909 28779 31912
rect 28721 31903 28779 31909
rect 28994 31900 29000 31912
rect 29052 31900 29058 31952
rect 31386 31900 31392 31952
rect 31444 31940 31450 31952
rect 31444 31912 31708 31940
rect 31444 31900 31450 31912
rect 27724 31844 28120 31872
rect 28445 31875 28503 31881
rect 27304 31776 27476 31804
rect 27617 31807 27675 31813
rect 27304 31764 27310 31776
rect 27617 31773 27629 31807
rect 27663 31773 27675 31807
rect 27617 31767 27675 31773
rect 27724 31736 27752 31844
rect 28445 31841 28457 31875
rect 28491 31872 28503 31875
rect 29086 31872 29092 31884
rect 28491 31844 29092 31872
rect 28491 31841 28503 31844
rect 28445 31835 28503 31841
rect 29086 31832 29092 31844
rect 29144 31832 29150 31884
rect 31570 31872 31576 31884
rect 31220 31844 31576 31872
rect 27847 31807 27905 31813
rect 27847 31773 27859 31807
rect 27893 31773 27905 31807
rect 27847 31767 27905 31773
rect 27862 31736 27890 31767
rect 28074 31764 28080 31816
rect 28132 31764 28138 31816
rect 28258 31804 28264 31816
rect 28219 31776 28264 31804
rect 28258 31764 28264 31776
rect 28316 31764 28322 31816
rect 28353 31807 28411 31813
rect 28353 31773 28365 31807
rect 28399 31804 28411 31807
rect 28534 31804 28540 31816
rect 28399 31776 28540 31804
rect 28399 31773 28411 31776
rect 28353 31767 28411 31773
rect 28534 31764 28540 31776
rect 28592 31764 28598 31816
rect 28626 31764 28632 31816
rect 28684 31764 28690 31816
rect 28810 31764 28816 31816
rect 28868 31764 28874 31816
rect 28905 31807 28963 31813
rect 28905 31773 28917 31807
rect 28951 31773 28963 31807
rect 28905 31767 28963 31773
rect 24636 31708 26096 31736
rect 26436 31708 27752 31736
rect 27816 31708 27890 31736
rect 27985 31739 28043 31745
rect 24636 31696 24642 31708
rect 23348 31640 23980 31668
rect 23348 31628 23354 31640
rect 24210 31628 24216 31680
rect 24268 31668 24274 31680
rect 26142 31668 26148 31680
rect 24268 31640 26148 31668
rect 24268 31628 24274 31640
rect 26142 31628 26148 31640
rect 26200 31668 26206 31680
rect 26436 31677 26464 31708
rect 26421 31671 26479 31677
rect 26421 31668 26433 31671
rect 26200 31640 26433 31668
rect 26200 31628 26206 31640
rect 26421 31637 26433 31640
rect 26467 31637 26479 31671
rect 26421 31631 26479 31637
rect 27062 31628 27068 31680
rect 27120 31628 27126 31680
rect 27338 31628 27344 31680
rect 27396 31668 27402 31680
rect 27816 31668 27844 31708
rect 27985 31705 27997 31739
rect 28031 31736 28043 31739
rect 28276 31736 28304 31764
rect 28920 31736 28948 31767
rect 28994 31764 29000 31816
rect 29052 31804 29058 31816
rect 29549 31807 29607 31813
rect 29549 31804 29561 31807
rect 29052 31776 29561 31804
rect 29052 31764 29058 31776
rect 29549 31773 29561 31776
rect 29595 31773 29607 31807
rect 29733 31807 29791 31813
rect 29733 31804 29745 31807
rect 29549 31767 29607 31773
rect 29656 31776 29745 31804
rect 28031 31708 28120 31736
rect 28276 31708 28948 31736
rect 28031 31705 28043 31708
rect 27985 31699 28043 31705
rect 28092 31680 28120 31708
rect 27396 31640 27844 31668
rect 27396 31628 27402 31640
rect 28074 31628 28080 31680
rect 28132 31628 28138 31680
rect 28626 31628 28632 31680
rect 28684 31668 28690 31680
rect 29656 31668 29684 31776
rect 29733 31773 29745 31776
rect 29779 31773 29791 31807
rect 29733 31767 29791 31773
rect 30006 31764 30012 31816
rect 30064 31804 30070 31816
rect 30469 31807 30527 31813
rect 30469 31804 30481 31807
rect 30064 31776 30481 31804
rect 30064 31764 30070 31776
rect 30469 31773 30481 31776
rect 30515 31773 30527 31807
rect 30469 31767 30527 31773
rect 31018 31764 31024 31816
rect 31076 31804 31082 31816
rect 31220 31813 31248 31844
rect 31570 31832 31576 31844
rect 31628 31832 31634 31884
rect 31680 31881 31708 31912
rect 31665 31875 31723 31881
rect 31665 31841 31677 31875
rect 31711 31841 31723 31875
rect 31772 31872 31800 31980
rect 32122 31968 32128 32020
rect 32180 31968 32186 32020
rect 32214 31968 32220 32020
rect 32272 31968 32278 32020
rect 32398 32008 32404 32020
rect 32324 31980 32404 32008
rect 32324 31940 32352 31980
rect 32398 31968 32404 31980
rect 32456 32008 32462 32020
rect 33134 32008 33140 32020
rect 32456 31980 33140 32008
rect 32456 31968 32462 31980
rect 33134 31968 33140 31980
rect 33192 31968 33198 32020
rect 34606 31968 34612 32020
rect 34664 32008 34670 32020
rect 34664 31980 36032 32008
rect 34664 31968 34670 31980
rect 32232 31912 32352 31940
rect 31849 31875 31907 31881
rect 31849 31872 31861 31875
rect 31772 31844 31861 31872
rect 31665 31835 31723 31841
rect 31849 31841 31861 31844
rect 31895 31841 31907 31875
rect 31849 31835 31907 31841
rect 31941 31875 31999 31881
rect 31941 31841 31953 31875
rect 31987 31872 31999 31875
rect 32232 31872 32260 31912
rect 32490 31900 32496 31952
rect 32548 31940 32554 31952
rect 32950 31940 32956 31952
rect 32548 31912 32956 31940
rect 32548 31900 32554 31912
rect 32950 31900 32956 31912
rect 33008 31940 33014 31952
rect 35437 31943 35495 31949
rect 33008 31912 33272 31940
rect 33008 31900 33014 31912
rect 32585 31875 32643 31881
rect 32585 31872 32597 31875
rect 31987 31844 32260 31872
rect 32324 31844 32597 31872
rect 31987 31841 31999 31844
rect 31941 31835 31999 31841
rect 31113 31807 31171 31813
rect 31113 31804 31125 31807
rect 31076 31776 31125 31804
rect 31076 31764 31082 31776
rect 31113 31773 31125 31776
rect 31159 31773 31171 31807
rect 31113 31767 31171 31773
rect 31205 31807 31263 31813
rect 31205 31773 31217 31807
rect 31251 31773 31263 31807
rect 31205 31767 31263 31773
rect 31386 31764 31392 31816
rect 31444 31764 31450 31816
rect 31481 31807 31539 31813
rect 31481 31773 31493 31807
rect 31527 31804 31539 31807
rect 31757 31807 31815 31813
rect 31527 31776 31616 31804
rect 31527 31773 31539 31776
rect 31481 31767 31539 31773
rect 31588 31748 31616 31776
rect 31757 31773 31769 31807
rect 31803 31773 31815 31807
rect 31757 31767 31815 31773
rect 30650 31696 30656 31748
rect 30708 31696 30714 31748
rect 31570 31696 31576 31748
rect 31628 31696 31634 31748
rect 28684 31640 29684 31668
rect 28684 31628 28690 31640
rect 31478 31628 31484 31680
rect 31536 31668 31542 31680
rect 31772 31668 31800 31767
rect 32214 31764 32220 31816
rect 32272 31804 32278 31816
rect 32324 31804 32352 31844
rect 32585 31841 32597 31844
rect 32631 31841 32643 31875
rect 33244 31872 33272 31912
rect 35437 31909 35449 31943
rect 35483 31940 35495 31943
rect 36004 31940 36032 31980
rect 36078 31968 36084 32020
rect 36136 31968 36142 32020
rect 37847 32011 37905 32017
rect 37847 31977 37859 32011
rect 37893 32008 37905 32011
rect 38010 32008 38016 32020
rect 37893 31980 38016 32008
rect 37893 31977 37905 31980
rect 37847 31971 37905 31977
rect 38010 31968 38016 31980
rect 38068 31968 38074 32020
rect 36722 31940 36728 31952
rect 35483 31912 35848 31940
rect 36004 31912 36728 31940
rect 35483 31909 35495 31912
rect 35437 31903 35495 31909
rect 33244 31844 33364 31872
rect 32585 31835 32643 31841
rect 32272 31776 32352 31804
rect 32401 31807 32459 31813
rect 32272 31764 32278 31776
rect 32401 31773 32413 31807
rect 32447 31773 32459 31807
rect 32401 31767 32459 31773
rect 32493 31807 32551 31813
rect 32493 31773 32505 31807
rect 32539 31773 32551 31807
rect 32493 31767 32551 31773
rect 32677 31807 32735 31813
rect 32677 31773 32689 31807
rect 32723 31804 32735 31807
rect 32861 31807 32919 31813
rect 32861 31804 32873 31807
rect 32723 31776 32873 31804
rect 32723 31773 32735 31776
rect 32677 31767 32735 31773
rect 32861 31773 32873 31776
rect 32907 31773 32919 31807
rect 32861 31767 32919 31773
rect 32030 31696 32036 31748
rect 32088 31736 32094 31748
rect 32416 31736 32444 31767
rect 32088 31708 32444 31736
rect 32508 31736 32536 31767
rect 32950 31764 32956 31816
rect 33008 31804 33014 31816
rect 33045 31807 33103 31813
rect 33045 31804 33057 31807
rect 33008 31776 33057 31804
rect 33008 31764 33014 31776
rect 33045 31773 33057 31776
rect 33091 31773 33103 31807
rect 33045 31767 33103 31773
rect 33226 31764 33232 31816
rect 33284 31764 33290 31816
rect 33336 31813 33364 31844
rect 34790 31832 34796 31884
rect 34848 31832 34854 31884
rect 34882 31832 34888 31884
rect 34940 31872 34946 31884
rect 34940 31844 35572 31872
rect 34940 31832 34946 31844
rect 33321 31807 33379 31813
rect 33321 31773 33333 31807
rect 33367 31773 33379 31807
rect 33321 31767 33379 31773
rect 34146 31764 34152 31816
rect 34204 31804 34210 31816
rect 35544 31813 35572 31844
rect 35820 31813 35848 31912
rect 36722 31900 36728 31912
rect 36780 31900 36786 31952
rect 38654 31940 38660 31952
rect 38626 31900 38660 31940
rect 38712 31900 38718 31952
rect 35986 31872 35992 31884
rect 35912 31844 35992 31872
rect 35912 31813 35940 31844
rect 35986 31832 35992 31844
rect 36044 31872 36050 31884
rect 36170 31872 36176 31884
rect 36044 31844 36176 31872
rect 36044 31832 36050 31844
rect 36170 31832 36176 31844
rect 36228 31872 36234 31884
rect 38626 31872 38654 31900
rect 36228 31844 38654 31872
rect 36228 31832 36234 31844
rect 35529 31807 35587 31813
rect 34204 31776 34744 31804
rect 34204 31764 34210 31776
rect 32766 31736 32772 31748
rect 32508 31708 32772 31736
rect 32088 31696 32094 31708
rect 32766 31696 32772 31708
rect 32824 31696 32830 31748
rect 34716 31736 34744 31776
rect 35529 31773 35541 31807
rect 35575 31773 35587 31807
rect 35529 31767 35587 31773
rect 35805 31807 35863 31813
rect 35805 31773 35817 31807
rect 35851 31773 35863 31807
rect 35805 31767 35863 31773
rect 35897 31807 35955 31813
rect 35897 31773 35909 31807
rect 35943 31773 35955 31807
rect 35897 31767 35955 31773
rect 36722 31764 36728 31816
rect 36780 31764 36786 31816
rect 38105 31807 38163 31813
rect 38105 31773 38117 31807
rect 38151 31804 38163 31807
rect 38194 31804 38200 31816
rect 38151 31776 38200 31804
rect 38151 31773 38163 31776
rect 38105 31767 38163 31773
rect 38194 31764 38200 31776
rect 38252 31764 38258 31816
rect 38286 31764 38292 31816
rect 38344 31764 38350 31816
rect 38473 31807 38531 31813
rect 38473 31804 38485 31807
rect 38396 31776 38485 31804
rect 35713 31739 35771 31745
rect 35713 31736 35725 31739
rect 34716 31708 35725 31736
rect 35713 31705 35725 31708
rect 35759 31736 35771 31739
rect 36538 31736 36544 31748
rect 35759 31708 36544 31736
rect 35759 31705 35771 31708
rect 35713 31699 35771 31705
rect 36538 31696 36544 31708
rect 36596 31696 36602 31748
rect 31536 31640 31800 31668
rect 31536 31628 31542 31640
rect 34238 31628 34244 31680
rect 34296 31668 34302 31680
rect 35434 31668 35440 31680
rect 34296 31640 35440 31668
rect 34296 31628 34302 31640
rect 35434 31628 35440 31640
rect 35492 31628 35498 31680
rect 35986 31628 35992 31680
rect 36044 31668 36050 31680
rect 36357 31671 36415 31677
rect 36357 31668 36369 31671
rect 36044 31640 36369 31668
rect 36044 31628 36050 31640
rect 36357 31637 36369 31640
rect 36403 31637 36415 31671
rect 36740 31668 36768 31764
rect 38396 31748 38424 31776
rect 38473 31773 38485 31776
rect 38519 31773 38531 31807
rect 38473 31767 38531 31773
rect 38562 31764 38568 31816
rect 38620 31764 38626 31816
rect 38654 31764 38660 31816
rect 38712 31764 38718 31816
rect 38378 31696 38384 31748
rect 38436 31696 38442 31748
rect 39482 31736 39488 31748
rect 38672 31708 39488 31736
rect 38672 31668 38700 31708
rect 39482 31696 39488 31708
rect 39540 31696 39546 31748
rect 36740 31640 38700 31668
rect 36357 31631 36415 31637
rect 38838 31628 38844 31680
rect 38896 31628 38902 31680
rect 1104 31578 40572 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 40572 31578
rect 1104 31504 40572 31526
rect 2866 31424 2872 31476
rect 2924 31464 2930 31476
rect 5258 31464 5264 31476
rect 2924 31436 5264 31464
rect 2924 31424 2930 31436
rect 5258 31424 5264 31436
rect 5316 31464 5322 31476
rect 5316 31436 5396 31464
rect 5316 31424 5322 31436
rect 2682 31356 2688 31408
rect 2740 31396 2746 31408
rect 5368 31405 5396 31436
rect 5718 31424 5724 31476
rect 5776 31424 5782 31476
rect 7282 31424 7288 31476
rect 7340 31464 7346 31476
rect 7377 31467 7435 31473
rect 7377 31464 7389 31467
rect 7340 31436 7389 31464
rect 7340 31424 7346 31436
rect 7377 31433 7389 31436
rect 7423 31433 7435 31467
rect 7377 31427 7435 31433
rect 7653 31467 7711 31473
rect 7653 31433 7665 31467
rect 7699 31464 7711 31467
rect 8386 31464 8392 31476
rect 7699 31436 8392 31464
rect 7699 31433 7711 31436
rect 7653 31427 7711 31433
rect 8386 31424 8392 31436
rect 8444 31424 8450 31476
rect 8665 31467 8723 31473
rect 8665 31433 8677 31467
rect 8711 31464 8723 31467
rect 10870 31464 10876 31476
rect 8711 31436 10876 31464
rect 8711 31433 8723 31436
rect 8665 31427 8723 31433
rect 10870 31424 10876 31436
rect 10928 31424 10934 31476
rect 10962 31424 10968 31476
rect 11020 31424 11026 31476
rect 11606 31424 11612 31476
rect 11664 31464 11670 31476
rect 11701 31467 11759 31473
rect 11701 31464 11713 31467
rect 11664 31436 11713 31464
rect 11664 31424 11670 31436
rect 11701 31433 11713 31436
rect 11747 31433 11759 31467
rect 11701 31427 11759 31433
rect 12710 31424 12716 31476
rect 12768 31424 12774 31476
rect 13541 31467 13599 31473
rect 13541 31433 13553 31467
rect 13587 31464 13599 31467
rect 13814 31464 13820 31476
rect 13587 31436 13820 31464
rect 13587 31433 13599 31436
rect 13541 31427 13599 31433
rect 13814 31424 13820 31436
rect 13872 31424 13878 31476
rect 14093 31467 14151 31473
rect 14093 31433 14105 31467
rect 14139 31464 14151 31467
rect 14182 31464 14188 31476
rect 14139 31436 14188 31464
rect 14139 31433 14151 31436
rect 14093 31427 14151 31433
rect 14182 31424 14188 31436
rect 14240 31424 14246 31476
rect 16758 31424 16764 31476
rect 16816 31424 16822 31476
rect 17957 31467 18015 31473
rect 17957 31433 17969 31467
rect 18003 31464 18015 31467
rect 18046 31464 18052 31476
rect 18003 31436 18052 31464
rect 18003 31433 18015 31436
rect 17957 31427 18015 31433
rect 18046 31424 18052 31436
rect 18104 31424 18110 31476
rect 19610 31424 19616 31476
rect 19668 31464 19674 31476
rect 19705 31467 19763 31473
rect 19705 31464 19717 31467
rect 19668 31436 19717 31464
rect 19668 31424 19674 31436
rect 19705 31433 19717 31436
rect 19751 31433 19763 31467
rect 19705 31427 19763 31433
rect 20073 31467 20131 31473
rect 20073 31433 20085 31467
rect 20119 31464 20131 31467
rect 21174 31464 21180 31476
rect 20119 31436 21180 31464
rect 20119 31433 20131 31436
rect 20073 31427 20131 31433
rect 21174 31424 21180 31436
rect 21232 31424 21238 31476
rect 21358 31424 21364 31476
rect 21416 31424 21422 31476
rect 21818 31424 21824 31476
rect 21876 31464 21882 31476
rect 22557 31467 22615 31473
rect 21876 31436 22508 31464
rect 21876 31424 21882 31436
rect 5353 31399 5411 31405
rect 2740 31368 3818 31396
rect 2740 31356 2746 31368
rect 5353 31365 5365 31399
rect 5399 31365 5411 31399
rect 5353 31359 5411 31365
rect 5569 31399 5627 31405
rect 5569 31365 5581 31399
rect 5615 31396 5627 31399
rect 5810 31396 5816 31408
rect 5615 31368 5816 31396
rect 5615 31365 5627 31368
rect 5569 31359 5627 31365
rect 5810 31356 5816 31368
rect 5868 31356 5874 31408
rect 6365 31399 6423 31405
rect 6365 31365 6377 31399
rect 6411 31396 6423 31399
rect 8570 31396 8576 31408
rect 6411 31368 8576 31396
rect 6411 31365 6423 31368
rect 6365 31359 6423 31365
rect 5442 31288 5448 31340
rect 5500 31328 5506 31340
rect 6380 31328 6408 31359
rect 8570 31356 8576 31368
rect 8628 31356 8634 31408
rect 8938 31356 8944 31408
rect 8996 31356 9002 31408
rect 9033 31399 9091 31405
rect 9033 31365 9045 31399
rect 9079 31396 9091 31399
rect 9079 31368 11100 31396
rect 9079 31365 9091 31368
rect 9033 31359 9091 31365
rect 5500 31300 6408 31328
rect 5500 31288 5506 31300
rect 7374 31288 7380 31340
rect 7432 31328 7438 31340
rect 8297 31331 8355 31337
rect 8297 31328 8309 31331
rect 7432 31300 8309 31328
rect 7432 31288 7438 31300
rect 8297 31297 8309 31300
rect 8343 31297 8355 31331
rect 8297 31291 8355 31297
rect 9309 31331 9367 31337
rect 9309 31297 9321 31331
rect 9355 31328 9367 31331
rect 9355 31300 9812 31328
rect 9355 31297 9367 31300
rect 9309 31291 9367 31297
rect 3234 31220 3240 31272
rect 3292 31220 3298 31272
rect 4982 31220 4988 31272
rect 5040 31220 5046 31272
rect 5261 31263 5319 31269
rect 5261 31229 5273 31263
rect 5307 31260 5319 31263
rect 5534 31260 5540 31272
rect 5307 31232 5540 31260
rect 5307 31229 5319 31232
rect 5261 31223 5319 31229
rect 5534 31220 5540 31232
rect 5592 31260 5598 31272
rect 5902 31260 5908 31272
rect 5592 31232 5908 31260
rect 5592 31220 5598 31232
rect 5902 31220 5908 31232
rect 5960 31260 5966 31272
rect 7101 31263 7159 31269
rect 7101 31260 7113 31263
rect 5960 31232 7113 31260
rect 5960 31220 5966 31232
rect 7101 31229 7113 31232
rect 7147 31229 7159 31263
rect 7101 31223 7159 31229
rect 7536 31263 7594 31269
rect 7536 31229 7548 31263
rect 7582 31260 7594 31263
rect 7582 31229 7604 31260
rect 7536 31223 7604 31229
rect 7576 31192 7604 31223
rect 7742 31220 7748 31272
rect 7800 31220 7806 31272
rect 7834 31220 7840 31272
rect 7892 31260 7898 31272
rect 8021 31263 8079 31269
rect 8021 31260 8033 31263
rect 7892 31232 8033 31260
rect 7892 31220 7898 31232
rect 8021 31229 8033 31232
rect 8067 31229 8079 31263
rect 8021 31223 8079 31229
rect 8389 31263 8447 31269
rect 8389 31229 8401 31263
rect 8435 31260 8447 31263
rect 8570 31260 8576 31272
rect 8435 31232 8576 31260
rect 8435 31229 8447 31232
rect 8389 31223 8447 31229
rect 8570 31220 8576 31232
rect 8628 31220 8634 31272
rect 9398 31220 9404 31272
rect 9456 31220 9462 31272
rect 9784 31260 9812 31300
rect 9950 31288 9956 31340
rect 10008 31288 10014 31340
rect 10413 31331 10471 31337
rect 10413 31297 10425 31331
rect 10459 31328 10471 31331
rect 10778 31328 10784 31340
rect 10459 31300 10784 31328
rect 10459 31297 10471 31300
rect 10413 31291 10471 31297
rect 10778 31288 10784 31300
rect 10836 31288 10842 31340
rect 10870 31288 10876 31340
rect 10928 31288 10934 31340
rect 11072 31328 11100 31368
rect 11146 31356 11152 31408
rect 11204 31396 11210 31408
rect 11330 31396 11336 31408
rect 11204 31368 11336 31396
rect 11204 31356 11210 31368
rect 11330 31356 11336 31368
rect 11388 31356 11394 31408
rect 11882 31356 11888 31408
rect 11940 31396 11946 31408
rect 11940 31368 12204 31396
rect 11940 31356 11946 31368
rect 11698 31328 11704 31340
rect 11072 31300 11704 31328
rect 9784 31232 10548 31260
rect 8662 31192 8668 31204
rect 7576 31164 8668 31192
rect 8662 31152 8668 31164
rect 8720 31152 8726 31204
rect 9858 31152 9864 31204
rect 9916 31152 9922 31204
rect 10520 31192 10548 31232
rect 10686 31220 10692 31272
rect 10744 31260 10750 31272
rect 10962 31260 10968 31272
rect 10744 31232 10968 31260
rect 10744 31220 10750 31232
rect 10962 31220 10968 31232
rect 11020 31220 11026 31272
rect 11054 31220 11060 31272
rect 11112 31260 11118 31272
rect 11164 31269 11192 31300
rect 11698 31288 11704 31300
rect 11756 31288 11762 31340
rect 12066 31288 12072 31340
rect 12124 31288 12130 31340
rect 12176 31337 12204 31368
rect 12526 31356 12532 31408
rect 12584 31396 12590 31408
rect 14277 31399 14335 31405
rect 14277 31396 14289 31399
rect 12584 31368 13400 31396
rect 12584 31356 12590 31368
rect 12161 31331 12219 31337
rect 12161 31297 12173 31331
rect 12207 31297 12219 31331
rect 12161 31291 12219 31297
rect 12894 31288 12900 31340
rect 12952 31288 12958 31340
rect 12986 31288 12992 31340
rect 13044 31288 13050 31340
rect 13372 31337 13400 31368
rect 13740 31368 14289 31396
rect 13740 31340 13768 31368
rect 14277 31365 14289 31368
rect 14323 31365 14335 31399
rect 15286 31396 15292 31408
rect 14277 31359 14335 31365
rect 15120 31368 15292 31396
rect 13265 31331 13323 31337
rect 13265 31297 13277 31331
rect 13311 31297 13323 31331
rect 13265 31291 13323 31297
rect 13357 31331 13415 31337
rect 13357 31297 13369 31331
rect 13403 31297 13415 31331
rect 13357 31291 13415 31297
rect 13541 31331 13599 31337
rect 13541 31297 13553 31331
rect 13587 31328 13599 31331
rect 13630 31328 13636 31340
rect 13587 31300 13636 31328
rect 13587 31297 13599 31300
rect 13541 31291 13599 31297
rect 11149 31263 11207 31269
rect 11149 31260 11161 31263
rect 11112 31232 11161 31260
rect 11112 31220 11118 31232
rect 11149 31229 11161 31232
rect 11195 31229 11207 31263
rect 11149 31223 11207 31229
rect 11330 31220 11336 31272
rect 11388 31260 11394 31272
rect 12084 31260 12112 31288
rect 11388 31232 12112 31260
rect 13280 31260 13308 31291
rect 13630 31288 13636 31300
rect 13688 31288 13694 31340
rect 13722 31288 13728 31340
rect 13780 31288 13786 31340
rect 13906 31337 13912 31340
rect 13879 31331 13912 31337
rect 13879 31297 13891 31331
rect 13964 31328 13970 31340
rect 13964 31300 14136 31328
rect 13879 31291 13912 31297
rect 13906 31288 13912 31291
rect 13964 31288 13970 31300
rect 14108 31260 14136 31300
rect 14182 31288 14188 31340
rect 14240 31288 14246 31340
rect 14369 31331 14427 31337
rect 14369 31297 14381 31331
rect 14415 31328 14427 31331
rect 14458 31328 14464 31340
rect 14415 31300 14464 31328
rect 14415 31297 14427 31300
rect 14369 31291 14427 31297
rect 14458 31288 14464 31300
rect 14516 31288 14522 31340
rect 14642 31260 14648 31272
rect 13280 31232 13400 31260
rect 14108 31232 14648 31260
rect 11388 31220 11394 31232
rect 13372 31192 13400 31232
rect 14642 31220 14648 31232
rect 14700 31220 14706 31272
rect 15010 31220 15016 31272
rect 15068 31260 15074 31272
rect 15120 31269 15148 31368
rect 15286 31356 15292 31368
rect 15344 31396 15350 31408
rect 19150 31396 19156 31408
rect 15344 31368 16712 31396
rect 15344 31356 15350 31368
rect 15470 31288 15476 31340
rect 15528 31328 15534 31340
rect 15565 31331 15623 31337
rect 15565 31328 15577 31331
rect 15528 31300 15577 31328
rect 15528 31288 15534 31300
rect 15565 31297 15577 31300
rect 15611 31297 15623 31331
rect 15565 31291 15623 31297
rect 15933 31331 15991 31337
rect 15933 31297 15945 31331
rect 15979 31328 15991 31331
rect 16022 31328 16028 31340
rect 15979 31300 16028 31328
rect 15979 31297 15991 31300
rect 15933 31291 15991 31297
rect 16022 31288 16028 31300
rect 16080 31288 16086 31340
rect 16684 31337 16712 31368
rect 17512 31368 19156 31396
rect 17512 31340 17540 31368
rect 19150 31356 19156 31368
rect 19208 31356 19214 31408
rect 19242 31356 19248 31408
rect 19300 31396 19306 31408
rect 21269 31399 21327 31405
rect 21269 31396 21281 31399
rect 19300 31368 21281 31396
rect 19300 31356 19306 31368
rect 21269 31365 21281 31368
rect 21315 31365 21327 31399
rect 21269 31359 21327 31365
rect 21959 31365 22017 31371
rect 16669 31331 16727 31337
rect 16669 31297 16681 31331
rect 16715 31297 16727 31331
rect 16669 31291 16727 31297
rect 16942 31288 16948 31340
rect 17000 31328 17006 31340
rect 17129 31331 17187 31337
rect 17129 31328 17141 31331
rect 17000 31300 17141 31328
rect 17000 31288 17006 31300
rect 17129 31297 17141 31300
rect 17175 31297 17187 31331
rect 17129 31291 17187 31297
rect 17494 31288 17500 31340
rect 17552 31288 17558 31340
rect 18230 31288 18236 31340
rect 18288 31288 18294 31340
rect 18414 31288 18420 31340
rect 18472 31328 18478 31340
rect 18509 31331 18567 31337
rect 18509 31328 18521 31331
rect 18472 31300 18521 31328
rect 18472 31288 18478 31300
rect 18509 31297 18521 31300
rect 18555 31328 18567 31331
rect 20717 31331 20775 31337
rect 20717 31328 20729 31331
rect 18555 31300 20729 31328
rect 18555 31297 18567 31300
rect 18509 31291 18567 31297
rect 20717 31297 20729 31300
rect 20763 31297 20775 31331
rect 20717 31291 20775 31297
rect 20809 31331 20867 31337
rect 20809 31297 20821 31331
rect 20855 31297 20867 31331
rect 20809 31291 20867 31297
rect 20901 31331 20959 31337
rect 20901 31297 20913 31331
rect 20947 31297 20959 31331
rect 20901 31291 20959 31297
rect 15105 31263 15163 31269
rect 15105 31260 15117 31263
rect 15068 31232 15117 31260
rect 15068 31220 15074 31232
rect 15105 31229 15117 31232
rect 15151 31229 15163 31263
rect 15105 31223 15163 31229
rect 15378 31220 15384 31272
rect 15436 31220 15442 31272
rect 15654 31220 15660 31272
rect 15712 31260 15718 31272
rect 15841 31263 15899 31269
rect 15841 31260 15853 31263
rect 15712 31232 15853 31260
rect 15712 31220 15718 31232
rect 15841 31229 15853 31232
rect 15887 31229 15899 31263
rect 15841 31223 15899 31229
rect 15197 31195 15255 31201
rect 15197 31192 15209 31195
rect 10520 31164 15209 31192
rect 15197 31161 15209 31164
rect 15243 31161 15255 31195
rect 15856 31192 15884 31223
rect 17218 31220 17224 31272
rect 17276 31220 17282 31272
rect 17405 31263 17463 31269
rect 17405 31229 17417 31263
rect 17451 31229 17463 31263
rect 17405 31223 17463 31229
rect 16298 31192 16304 31204
rect 15856 31164 16304 31192
rect 15197 31155 15255 31161
rect 16298 31152 16304 31164
rect 16356 31192 16362 31204
rect 17420 31192 17448 31223
rect 17862 31220 17868 31272
rect 17920 31260 17926 31272
rect 18141 31263 18199 31269
rect 18141 31260 18153 31263
rect 17920 31232 18153 31260
rect 17920 31220 17926 31232
rect 18141 31229 18153 31232
rect 18187 31229 18199 31263
rect 18141 31223 18199 31229
rect 18601 31263 18659 31269
rect 18601 31229 18613 31263
rect 18647 31260 18659 31263
rect 18785 31263 18843 31269
rect 18785 31260 18797 31263
rect 18647 31232 18797 31260
rect 18647 31229 18659 31232
rect 18601 31223 18659 31229
rect 18785 31229 18797 31232
rect 18831 31229 18843 31263
rect 18785 31223 18843 31229
rect 16356 31164 17448 31192
rect 18156 31192 18184 31223
rect 19058 31220 19064 31272
rect 19116 31260 19122 31272
rect 19337 31263 19395 31269
rect 19337 31260 19349 31263
rect 19116 31232 19349 31260
rect 19116 31220 19122 31232
rect 19337 31229 19349 31232
rect 19383 31229 19395 31263
rect 19337 31223 19395 31229
rect 20165 31263 20223 31269
rect 20165 31229 20177 31263
rect 20211 31229 20223 31263
rect 20165 31223 20223 31229
rect 20180 31192 20208 31223
rect 20346 31220 20352 31272
rect 20404 31220 20410 31272
rect 20438 31220 20444 31272
rect 20496 31260 20502 31272
rect 20824 31260 20852 31291
rect 20496 31232 20852 31260
rect 20496 31220 20502 31232
rect 20916 31192 20944 31291
rect 20990 31288 20996 31340
rect 21048 31328 21054 31340
rect 21085 31331 21143 31337
rect 21085 31328 21097 31331
rect 21048 31300 21097 31328
rect 21048 31288 21054 31300
rect 21085 31297 21097 31300
rect 21131 31297 21143 31331
rect 21959 31331 21971 31365
rect 22005 31362 22017 31365
rect 22005 31331 22032 31362
rect 22094 31356 22100 31408
rect 22152 31396 22158 31408
rect 22189 31399 22247 31405
rect 22189 31396 22201 31399
rect 22152 31368 22201 31396
rect 22152 31356 22158 31368
rect 22189 31365 22201 31368
rect 22235 31365 22247 31399
rect 22480 31396 22508 31436
rect 22557 31433 22569 31467
rect 22603 31464 22615 31467
rect 22922 31464 22928 31476
rect 22603 31436 22928 31464
rect 22603 31433 22615 31436
rect 22557 31427 22615 31433
rect 22922 31424 22928 31436
rect 22980 31424 22986 31476
rect 23842 31464 23848 31476
rect 23032 31436 23848 31464
rect 23032 31396 23060 31436
rect 23842 31424 23848 31436
rect 23900 31424 23906 31476
rect 24029 31467 24087 31473
rect 24029 31433 24041 31467
rect 24075 31464 24087 31467
rect 24075 31436 25084 31464
rect 24075 31433 24087 31436
rect 24029 31427 24087 31433
rect 24946 31396 24952 31408
rect 22480 31368 23060 31396
rect 23676 31368 24952 31396
rect 22189 31359 22247 31365
rect 21959 31325 22032 31331
rect 21085 31291 21143 31297
rect 22004 31260 22032 31325
rect 22281 31331 22339 31337
rect 22281 31297 22293 31331
rect 22327 31328 22339 31331
rect 22922 31328 22928 31340
rect 22327 31300 22928 31328
rect 22327 31297 22339 31300
rect 22281 31291 22339 31297
rect 22922 31288 22928 31300
rect 22980 31288 22986 31340
rect 23106 31288 23112 31340
rect 23164 31288 23170 31340
rect 23290 31288 23296 31340
rect 23348 31288 23354 31340
rect 23566 31288 23572 31340
rect 23624 31328 23630 31340
rect 23676 31337 23704 31368
rect 24946 31356 24952 31368
rect 25004 31356 25010 31408
rect 23661 31331 23719 31337
rect 23661 31328 23673 31331
rect 23624 31300 23673 31328
rect 23624 31288 23630 31300
rect 23661 31297 23673 31300
rect 23707 31297 23719 31331
rect 24857 31331 24915 31337
rect 24857 31328 24869 31331
rect 23661 31291 23719 31297
rect 24228 31300 24869 31328
rect 22370 31260 22376 31272
rect 22004 31232 22376 31260
rect 22370 31220 22376 31232
rect 22428 31220 22434 31272
rect 22554 31220 22560 31272
rect 22612 31220 22618 31272
rect 23842 31220 23848 31272
rect 23900 31220 23906 31272
rect 24121 31263 24179 31269
rect 24121 31229 24133 31263
rect 24167 31229 24179 31263
rect 24121 31223 24179 31229
rect 22186 31192 22192 31204
rect 18156 31164 20944 31192
rect 21284 31164 22192 31192
rect 16356 31152 16362 31164
rect 4890 31084 4896 31136
rect 4948 31124 4954 31136
rect 5537 31127 5595 31133
rect 5537 31124 5549 31127
rect 4948 31096 5549 31124
rect 4948 31084 4954 31096
rect 5537 31093 5549 31096
rect 5583 31124 5595 31127
rect 7374 31124 7380 31136
rect 5583 31096 7380 31124
rect 5583 31093 5595 31096
rect 5537 31087 5595 31093
rect 7374 31084 7380 31096
rect 7432 31084 7438 31136
rect 9582 31084 9588 31136
rect 9640 31084 9646 31136
rect 9950 31084 9956 31136
rect 10008 31124 10014 31136
rect 11238 31124 11244 31136
rect 10008 31096 11244 31124
rect 10008 31084 10014 31096
rect 11238 31084 11244 31096
rect 11296 31084 11302 31136
rect 11514 31084 11520 31136
rect 11572 31084 11578 31136
rect 13173 31127 13231 31133
rect 13173 31093 13185 31127
rect 13219 31124 13231 31127
rect 13906 31124 13912 31136
rect 13219 31096 13912 31124
rect 13219 31093 13231 31096
rect 13173 31087 13231 31093
rect 13906 31084 13912 31096
rect 13964 31084 13970 31136
rect 16022 31084 16028 31136
rect 16080 31124 16086 31136
rect 19518 31124 19524 31136
rect 16080 31096 19524 31124
rect 16080 31084 16086 31096
rect 19518 31084 19524 31096
rect 19576 31084 19582 31136
rect 20533 31127 20591 31133
rect 20533 31093 20545 31127
rect 20579 31124 20591 31127
rect 20806 31124 20812 31136
rect 20579 31096 20812 31124
rect 20579 31093 20591 31096
rect 20533 31087 20591 31093
rect 20806 31084 20812 31096
rect 20864 31084 20870 31136
rect 20898 31084 20904 31136
rect 20956 31124 20962 31136
rect 21284 31124 21312 31164
rect 20956 31096 21312 31124
rect 20956 31084 20962 31096
rect 21634 31084 21640 31136
rect 21692 31124 21698 31136
rect 22020 31133 22048 31164
rect 22186 31152 22192 31164
rect 22244 31152 22250 31204
rect 23198 31152 23204 31204
rect 23256 31192 23262 31204
rect 24136 31192 24164 31223
rect 23256 31164 24164 31192
rect 23256 31152 23262 31164
rect 21821 31127 21879 31133
rect 21821 31124 21833 31127
rect 21692 31096 21833 31124
rect 21692 31084 21698 31096
rect 21821 31093 21833 31096
rect 21867 31093 21879 31127
rect 21821 31087 21879 31093
rect 22005 31127 22063 31133
rect 22005 31093 22017 31127
rect 22051 31093 22063 31127
rect 22005 31087 22063 31093
rect 22370 31084 22376 31136
rect 22428 31084 22434 31136
rect 23014 31084 23020 31136
rect 23072 31124 23078 31136
rect 24228 31124 24256 31300
rect 24857 31297 24869 31300
rect 24903 31297 24915 31331
rect 24857 31291 24915 31297
rect 23072 31096 24256 31124
rect 23072 31084 23078 31096
rect 24302 31084 24308 31136
rect 24360 31084 24366 31136
rect 24872 31124 24900 31291
rect 24946 31220 24952 31272
rect 25004 31220 25010 31272
rect 25056 31260 25084 31436
rect 25774 31424 25780 31476
rect 25832 31464 25838 31476
rect 25869 31467 25927 31473
rect 25869 31464 25881 31467
rect 25832 31436 25881 31464
rect 25832 31424 25838 31436
rect 25869 31433 25881 31436
rect 25915 31433 25927 31467
rect 25869 31427 25927 31433
rect 26050 31424 26056 31476
rect 26108 31464 26114 31476
rect 26145 31467 26203 31473
rect 26145 31464 26157 31467
rect 26108 31436 26157 31464
rect 26108 31424 26114 31436
rect 26145 31433 26157 31436
rect 26191 31433 26203 31467
rect 28442 31464 28448 31476
rect 26145 31427 26203 31433
rect 26252 31436 28448 31464
rect 25406 31356 25412 31408
rect 25464 31396 25470 31408
rect 26252 31396 26280 31436
rect 27474 31405 27502 31436
rect 28442 31424 28448 31436
rect 28500 31424 28506 31476
rect 29638 31424 29644 31476
rect 29696 31424 29702 31476
rect 34451 31467 34509 31473
rect 33704 31436 34376 31464
rect 27459 31399 27517 31405
rect 25464 31368 26280 31396
rect 26436 31368 27200 31396
rect 25464 31356 25470 31368
rect 25225 31331 25283 31337
rect 25225 31297 25237 31331
rect 25271 31328 25283 31331
rect 25682 31328 25688 31340
rect 25271 31300 25688 31328
rect 25271 31297 25283 31300
rect 25225 31291 25283 31297
rect 25682 31288 25688 31300
rect 25740 31288 25746 31340
rect 25777 31331 25835 31337
rect 25777 31297 25789 31331
rect 25823 31297 25835 31331
rect 25777 31291 25835 31297
rect 25317 31263 25375 31269
rect 25317 31260 25329 31263
rect 25056 31232 25329 31260
rect 25317 31229 25329 31232
rect 25363 31229 25375 31263
rect 25792 31260 25820 31291
rect 25958 31288 25964 31340
rect 26016 31288 26022 31340
rect 26436 31337 26464 31368
rect 27172 31340 27200 31368
rect 27459 31365 27471 31399
rect 27505 31365 27517 31399
rect 27459 31359 27517 31365
rect 28810 31356 28816 31408
rect 28868 31396 28874 31408
rect 28868 31368 33640 31396
rect 28868 31356 28874 31368
rect 26421 31331 26479 31337
rect 26421 31297 26433 31331
rect 26467 31297 26479 31331
rect 26421 31291 26479 31297
rect 26510 31288 26516 31340
rect 26568 31288 26574 31340
rect 26602 31288 26608 31340
rect 26660 31288 26666 31340
rect 26789 31331 26847 31337
rect 26789 31297 26801 31331
rect 26835 31328 26847 31331
rect 27062 31328 27068 31340
rect 26835 31300 27068 31328
rect 26835 31297 26847 31300
rect 26789 31291 26847 31297
rect 27062 31288 27068 31300
rect 27120 31288 27126 31340
rect 27154 31288 27160 31340
rect 27212 31288 27218 31340
rect 27246 31288 27252 31340
rect 27304 31288 27310 31340
rect 27341 31331 27399 31337
rect 27341 31297 27353 31331
rect 27387 31297 27399 31331
rect 27341 31291 27399 31297
rect 27356 31260 27384 31291
rect 28258 31288 28264 31340
rect 28316 31288 28322 31340
rect 28442 31288 28448 31340
rect 28500 31288 28506 31340
rect 29270 31288 29276 31340
rect 29328 31328 29334 31340
rect 29549 31331 29607 31337
rect 29549 31328 29561 31331
rect 29328 31300 29561 31328
rect 29328 31288 29334 31300
rect 29549 31297 29561 31300
rect 29595 31297 29607 31331
rect 29549 31291 29607 31297
rect 29733 31331 29791 31337
rect 29733 31297 29745 31331
rect 29779 31328 29791 31331
rect 30742 31328 30748 31340
rect 29779 31300 30748 31328
rect 29779 31297 29791 31300
rect 29733 31291 29791 31297
rect 30742 31288 30748 31300
rect 30800 31288 30806 31340
rect 30834 31288 30840 31340
rect 30892 31328 30898 31340
rect 32766 31328 32772 31340
rect 30892 31300 32772 31328
rect 30892 31288 30898 31300
rect 32766 31288 32772 31300
rect 32824 31328 32830 31340
rect 33413 31331 33471 31337
rect 33413 31328 33425 31331
rect 32824 31300 33425 31328
rect 32824 31288 32830 31300
rect 33413 31297 33425 31300
rect 33459 31297 33471 31331
rect 33413 31291 33471 31297
rect 25792 31232 27384 31260
rect 25317 31223 25375 31229
rect 26970 31152 26976 31204
rect 27028 31152 27034 31204
rect 26694 31124 26700 31136
rect 24872 31096 26700 31124
rect 26694 31084 26700 31096
rect 26752 31084 26758 31136
rect 27356 31124 27384 31232
rect 27430 31220 27436 31272
rect 27488 31260 27494 31272
rect 27617 31263 27675 31269
rect 27617 31260 27629 31263
rect 27488 31232 27629 31260
rect 27488 31220 27494 31232
rect 27617 31229 27629 31232
rect 27663 31229 27675 31263
rect 27617 31223 27675 31229
rect 27632 31192 27660 31223
rect 27706 31220 27712 31272
rect 27764 31260 27770 31272
rect 28276 31260 28304 31288
rect 28810 31260 28816 31272
rect 27764 31232 28816 31260
rect 27764 31220 27770 31232
rect 28810 31220 28816 31232
rect 28868 31220 28874 31272
rect 31570 31220 31576 31272
rect 31628 31260 31634 31272
rect 33229 31263 33287 31269
rect 33229 31260 33241 31263
rect 31628 31232 33241 31260
rect 31628 31220 31634 31232
rect 33229 31229 33241 31232
rect 33275 31229 33287 31263
rect 33229 31223 33287 31229
rect 27801 31195 27859 31201
rect 27801 31192 27813 31195
rect 27632 31164 27813 31192
rect 27801 31161 27813 31164
rect 27847 31161 27859 31195
rect 27801 31155 27859 31161
rect 27890 31152 27896 31204
rect 27948 31152 27954 31204
rect 28258 31192 28264 31204
rect 28000 31164 28264 31192
rect 28000 31124 28028 31164
rect 28258 31152 28264 31164
rect 28316 31152 28322 31204
rect 33428 31192 33456 31291
rect 33612 31260 33640 31368
rect 33704 31337 33732 31436
rect 33778 31356 33784 31408
rect 33836 31396 33842 31408
rect 34238 31396 34244 31408
rect 33836 31368 34244 31396
rect 33836 31356 33842 31368
rect 34238 31356 34244 31368
rect 34296 31356 34302 31408
rect 34348 31396 34376 31436
rect 34451 31433 34463 31467
rect 34497 31464 34509 31467
rect 34701 31467 34759 31473
rect 34701 31464 34713 31467
rect 34497 31436 34713 31464
rect 34497 31433 34509 31436
rect 34451 31427 34509 31433
rect 34701 31433 34713 31436
rect 34747 31464 34759 31467
rect 34882 31464 34888 31476
rect 34747 31436 34888 31464
rect 34747 31433 34759 31436
rect 34701 31427 34759 31433
rect 34882 31424 34888 31436
rect 34940 31424 34946 31476
rect 35434 31424 35440 31476
rect 35492 31464 35498 31476
rect 37093 31467 37151 31473
rect 35492 31436 36308 31464
rect 35492 31424 35498 31436
rect 34790 31396 34796 31408
rect 34348 31368 34796 31396
rect 34790 31356 34796 31368
rect 34848 31356 34854 31408
rect 36170 31405 36176 31408
rect 36147 31399 36176 31405
rect 36147 31365 36159 31399
rect 36147 31359 36176 31365
rect 36170 31356 36176 31359
rect 36228 31356 36234 31408
rect 36280 31405 36308 31436
rect 37093 31433 37105 31467
rect 37139 31464 37151 31467
rect 37734 31464 37740 31476
rect 37139 31436 37740 31464
rect 37139 31433 37151 31436
rect 37093 31427 37151 31433
rect 37734 31424 37740 31436
rect 37792 31424 37798 31476
rect 37826 31424 37832 31476
rect 37884 31464 37890 31476
rect 38378 31464 38384 31476
rect 37884 31436 38384 31464
rect 37884 31424 37890 31436
rect 38378 31424 38384 31436
rect 38436 31424 38442 31476
rect 38562 31424 38568 31476
rect 38620 31464 38626 31476
rect 40221 31467 40279 31473
rect 40221 31464 40233 31467
rect 38620 31436 40233 31464
rect 38620 31424 38626 31436
rect 40221 31433 40233 31436
rect 40267 31433 40279 31467
rect 40221 31427 40279 31433
rect 36265 31399 36323 31405
rect 36265 31365 36277 31399
rect 36311 31396 36323 31399
rect 36909 31399 36967 31405
rect 36311 31368 36860 31396
rect 36311 31365 36323 31368
rect 36265 31359 36323 31365
rect 33689 31331 33747 31337
rect 33689 31297 33701 31331
rect 33735 31297 33747 31331
rect 33689 31291 33747 31297
rect 34330 31288 34336 31340
rect 34388 31328 34394 31340
rect 34885 31331 34943 31337
rect 34885 31328 34897 31331
rect 34388 31300 34897 31328
rect 34388 31288 34394 31300
rect 34885 31297 34897 31300
rect 34931 31297 34943 31331
rect 35986 31328 35992 31340
rect 34885 31291 34943 31297
rect 34992 31300 35992 31328
rect 34992 31260 35020 31300
rect 35986 31288 35992 31300
rect 36044 31288 36050 31340
rect 36354 31288 36360 31340
rect 36412 31288 36418 31340
rect 36446 31288 36452 31340
rect 36504 31288 36510 31340
rect 36633 31331 36691 31337
rect 36633 31297 36645 31331
rect 36679 31328 36691 31331
rect 36725 31331 36783 31337
rect 36725 31328 36737 31331
rect 36679 31300 36737 31328
rect 36679 31297 36691 31300
rect 36633 31291 36691 31297
rect 36725 31297 36737 31300
rect 36771 31297 36783 31331
rect 36832 31328 36860 31368
rect 36909 31365 36921 31399
rect 36955 31396 36967 31399
rect 37182 31396 37188 31408
rect 36955 31368 37188 31396
rect 36955 31365 36967 31368
rect 36909 31359 36967 31365
rect 37182 31356 37188 31368
rect 37240 31356 37246 31408
rect 37553 31399 37611 31405
rect 37553 31365 37565 31399
rect 37599 31365 37611 31399
rect 37553 31359 37611 31365
rect 38749 31399 38807 31405
rect 38749 31365 38761 31399
rect 38795 31396 38807 31399
rect 38838 31396 38844 31408
rect 38795 31368 38844 31396
rect 38795 31365 38807 31368
rect 38749 31359 38807 31365
rect 37277 31331 37335 31337
rect 37277 31328 37289 31331
rect 36832 31300 37289 31328
rect 36725 31291 36783 31297
rect 37277 31297 37289 31300
rect 37323 31328 37335 31331
rect 37366 31328 37372 31340
rect 37323 31300 37372 31328
rect 37323 31297 37335 31300
rect 37277 31291 37335 31297
rect 37366 31288 37372 31300
rect 37424 31288 37430 31340
rect 37461 31331 37519 31337
rect 37461 31297 37473 31331
rect 37507 31297 37519 31331
rect 37461 31291 37519 31297
rect 33612 31232 35020 31260
rect 35069 31263 35127 31269
rect 35069 31229 35081 31263
rect 35115 31260 35127 31263
rect 35434 31260 35440 31272
rect 35115 31232 35440 31260
rect 35115 31229 35127 31232
rect 35069 31223 35127 31229
rect 35434 31220 35440 31232
rect 35492 31220 35498 31272
rect 37476 31260 37504 31291
rect 37568 31272 37596 31359
rect 38838 31356 38844 31368
rect 38896 31356 38902 31408
rect 39482 31356 39488 31408
rect 39540 31356 39546 31408
rect 37645 31331 37703 31337
rect 37645 31297 37657 31331
rect 37691 31297 37703 31331
rect 37645 31291 37703 31297
rect 36464 31232 37504 31260
rect 36464 31192 36492 31232
rect 37550 31220 37556 31272
rect 37608 31220 37614 31272
rect 33428 31164 36492 31192
rect 37458 31152 37464 31204
rect 37516 31192 37522 31204
rect 37660 31192 37688 31291
rect 38194 31288 38200 31340
rect 38252 31328 38258 31340
rect 38473 31331 38531 31337
rect 38473 31328 38485 31331
rect 38252 31300 38485 31328
rect 38252 31288 38258 31300
rect 38473 31297 38485 31300
rect 38519 31297 38531 31331
rect 38473 31291 38531 31297
rect 37516 31164 37688 31192
rect 37516 31152 37522 31164
rect 27356 31096 28028 31124
rect 28074 31084 28080 31136
rect 28132 31124 28138 31136
rect 28537 31127 28595 31133
rect 28537 31124 28549 31127
rect 28132 31096 28549 31124
rect 28132 31084 28138 31096
rect 28537 31093 28549 31096
rect 28583 31124 28595 31127
rect 28718 31124 28724 31136
rect 28583 31096 28724 31124
rect 28583 31093 28595 31096
rect 28537 31087 28595 31093
rect 28718 31084 28724 31096
rect 28776 31084 28782 31136
rect 31570 31084 31576 31136
rect 31628 31124 31634 31136
rect 33318 31124 33324 31136
rect 31628 31096 33324 31124
rect 31628 31084 31634 31096
rect 33318 31084 33324 31096
rect 33376 31084 33382 31136
rect 33594 31084 33600 31136
rect 33652 31084 33658 31136
rect 34146 31084 34152 31136
rect 34204 31124 34210 31136
rect 34425 31127 34483 31133
rect 34425 31124 34437 31127
rect 34204 31096 34437 31124
rect 34204 31084 34210 31096
rect 34425 31093 34437 31096
rect 34471 31093 34483 31127
rect 34425 31087 34483 31093
rect 34609 31127 34667 31133
rect 34609 31093 34621 31127
rect 34655 31124 34667 31127
rect 34790 31124 34796 31136
rect 34655 31096 34796 31124
rect 34655 31093 34667 31096
rect 34609 31087 34667 31093
rect 34790 31084 34796 31096
rect 34848 31084 34854 31136
rect 37274 31084 37280 31136
rect 37332 31124 37338 31136
rect 37829 31127 37887 31133
rect 37829 31124 37841 31127
rect 37332 31096 37841 31124
rect 37332 31084 37338 31096
rect 37829 31093 37841 31096
rect 37875 31124 37887 31127
rect 38562 31124 38568 31136
rect 37875 31096 38568 31124
rect 37875 31093 37887 31096
rect 37829 31087 37887 31093
rect 38562 31084 38568 31096
rect 38620 31084 38626 31136
rect 1104 31034 40572 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 40572 31034
rect 1104 30960 40572 30982
rect 4157 30923 4215 30929
rect 4157 30889 4169 30923
rect 4203 30920 4215 30923
rect 4982 30920 4988 30932
rect 4203 30892 4988 30920
rect 4203 30889 4215 30892
rect 4157 30883 4215 30889
rect 4982 30880 4988 30892
rect 5040 30880 5046 30932
rect 7929 30923 7987 30929
rect 7929 30889 7941 30923
rect 7975 30920 7987 30923
rect 8018 30920 8024 30932
rect 7975 30892 8024 30920
rect 7975 30889 7987 30892
rect 7929 30883 7987 30889
rect 8018 30880 8024 30892
rect 8076 30880 8082 30932
rect 8570 30880 8576 30932
rect 8628 30880 8634 30932
rect 10778 30880 10784 30932
rect 10836 30880 10842 30932
rect 11330 30880 11336 30932
rect 11388 30880 11394 30932
rect 11882 30880 11888 30932
rect 11940 30920 11946 30932
rect 15197 30923 15255 30929
rect 15197 30920 15209 30923
rect 11940 30892 15209 30920
rect 11940 30880 11946 30892
rect 15197 30889 15209 30892
rect 15243 30889 15255 30923
rect 15197 30883 15255 30889
rect 15470 30880 15476 30932
rect 15528 30880 15534 30932
rect 17402 30880 17408 30932
rect 17460 30920 17466 30932
rect 17862 30920 17868 30932
rect 17460 30892 17868 30920
rect 17460 30880 17466 30892
rect 17862 30880 17868 30892
rect 17920 30880 17926 30932
rect 18414 30880 18420 30932
rect 18472 30880 18478 30932
rect 18690 30880 18696 30932
rect 18748 30880 18754 30932
rect 18877 30923 18935 30929
rect 18877 30889 18889 30923
rect 18923 30920 18935 30923
rect 20990 30920 20996 30932
rect 18923 30892 20996 30920
rect 18923 30889 18935 30892
rect 18877 30883 18935 30889
rect 20990 30880 20996 30892
rect 21048 30880 21054 30932
rect 22830 30880 22836 30932
rect 22888 30880 22894 30932
rect 23109 30923 23167 30929
rect 23109 30889 23121 30923
rect 23155 30920 23167 30923
rect 23198 30920 23204 30932
rect 23155 30892 23204 30920
rect 23155 30889 23167 30892
rect 23109 30883 23167 30889
rect 23198 30880 23204 30892
rect 23256 30880 23262 30932
rect 23293 30923 23351 30929
rect 23293 30889 23305 30923
rect 23339 30920 23351 30923
rect 23658 30920 23664 30932
rect 23339 30892 23664 30920
rect 23339 30889 23351 30892
rect 23293 30883 23351 30889
rect 23658 30880 23664 30892
rect 23716 30880 23722 30932
rect 23842 30880 23848 30932
rect 23900 30920 23906 30932
rect 24581 30923 24639 30929
rect 24581 30920 24593 30923
rect 23900 30892 24593 30920
rect 23900 30880 23906 30892
rect 24581 30889 24593 30892
rect 24627 30889 24639 30923
rect 24581 30883 24639 30889
rect 26510 30880 26516 30932
rect 26568 30920 26574 30932
rect 26605 30923 26663 30929
rect 26605 30920 26617 30923
rect 26568 30892 26617 30920
rect 26568 30880 26574 30892
rect 26605 30889 26617 30892
rect 26651 30889 26663 30923
rect 26605 30883 26663 30889
rect 26694 30880 26700 30932
rect 26752 30920 26758 30932
rect 26752 30892 31340 30920
rect 26752 30880 26758 30892
rect 8386 30852 8392 30864
rect 8036 30824 8392 30852
rect 3234 30744 3240 30796
rect 3292 30784 3298 30796
rect 4617 30787 4675 30793
rect 4617 30784 4629 30787
rect 3292 30756 4629 30784
rect 3292 30744 3298 30756
rect 4617 30753 4629 30756
rect 4663 30753 4675 30787
rect 4617 30747 4675 30753
rect 4798 30744 4804 30796
rect 4856 30744 4862 30796
rect 7377 30787 7435 30793
rect 7377 30753 7389 30787
rect 7423 30753 7435 30787
rect 7377 30747 7435 30753
rect 3605 30719 3663 30725
rect 3605 30685 3617 30719
rect 3651 30716 3663 30719
rect 3786 30716 3792 30728
rect 3651 30688 3792 30716
rect 3651 30685 3663 30688
rect 3605 30679 3663 30685
rect 3786 30676 3792 30688
rect 3844 30676 3850 30728
rect 4525 30719 4583 30725
rect 4525 30685 4537 30719
rect 4571 30716 4583 30719
rect 4890 30716 4896 30728
rect 4571 30688 4896 30716
rect 4571 30685 4583 30688
rect 4525 30679 4583 30685
rect 4890 30676 4896 30688
rect 4948 30676 4954 30728
rect 6086 30676 6092 30728
rect 6144 30716 6150 30728
rect 6546 30716 6552 30728
rect 6144 30688 6552 30716
rect 6144 30676 6150 30688
rect 6546 30676 6552 30688
rect 6604 30676 6610 30728
rect 7392 30716 7420 30747
rect 7650 30716 7656 30728
rect 7392 30688 7656 30716
rect 7650 30676 7656 30688
rect 7708 30676 7714 30728
rect 8036 30725 8064 30824
rect 8386 30812 8392 30824
rect 8444 30852 8450 30864
rect 8754 30852 8760 30864
rect 8444 30824 8760 30852
rect 8444 30812 8450 30824
rect 8754 30812 8760 30824
rect 8812 30852 8818 30864
rect 9122 30852 9128 30864
rect 8812 30824 9128 30852
rect 8812 30812 8818 30824
rect 9122 30812 9128 30824
rect 9180 30812 9186 30864
rect 10502 30852 10508 30864
rect 9876 30824 10508 30852
rect 8294 30744 8300 30796
rect 8352 30784 8358 30796
rect 8352 30756 8616 30784
rect 8352 30744 8358 30756
rect 8021 30719 8079 30725
rect 8021 30685 8033 30719
rect 8067 30685 8079 30719
rect 8021 30679 8079 30685
rect 8202 30676 8208 30728
rect 8260 30676 8266 30728
rect 8588 30725 8616 30756
rect 9674 30744 9680 30796
rect 9732 30744 9738 30796
rect 9876 30725 9904 30824
rect 10502 30812 10508 30824
rect 10560 30852 10566 30864
rect 10962 30852 10968 30864
rect 10560 30824 10968 30852
rect 10560 30812 10566 30824
rect 10962 30812 10968 30824
rect 11020 30812 11026 30864
rect 11514 30784 11520 30796
rect 10336 30756 11520 30784
rect 10336 30725 10364 30756
rect 11514 30744 11520 30756
rect 11572 30744 11578 30796
rect 8389 30719 8447 30725
rect 8389 30685 8401 30719
rect 8435 30685 8447 30719
rect 8389 30679 8447 30685
rect 8573 30719 8631 30725
rect 8573 30685 8585 30719
rect 8619 30685 8631 30719
rect 8573 30679 8631 30685
rect 9861 30719 9919 30725
rect 9861 30685 9873 30719
rect 9907 30685 9919 30719
rect 9861 30679 9919 30685
rect 10321 30719 10379 30725
rect 10321 30685 10333 30719
rect 10367 30685 10379 30719
rect 10321 30679 10379 30685
rect 1578 30608 1584 30660
rect 1636 30608 1642 30660
rect 2682 30608 2688 30660
rect 2740 30608 2746 30660
rect 3326 30608 3332 30660
rect 3384 30608 3390 30660
rect 7561 30651 7619 30657
rect 7561 30617 7573 30651
rect 7607 30648 7619 30651
rect 8113 30651 8171 30657
rect 8113 30648 8125 30651
rect 7607 30620 8125 30648
rect 7607 30617 7619 30620
rect 7561 30611 7619 30617
rect 8113 30617 8125 30620
rect 8159 30648 8171 30651
rect 8404 30648 8432 30679
rect 8159 30620 8432 30648
rect 8159 30617 8171 30620
rect 8113 30611 8171 30617
rect 6178 30540 6184 30592
rect 6236 30540 6242 30592
rect 7469 30583 7527 30589
rect 7469 30549 7481 30583
rect 7515 30580 7527 30583
rect 8588 30580 8616 30679
rect 10686 30676 10692 30728
rect 10744 30676 10750 30728
rect 10962 30719 11020 30725
rect 10962 30685 10974 30719
rect 11008 30716 11020 30719
rect 11054 30716 11060 30728
rect 11008 30688 11060 30716
rect 11008 30685 11020 30688
rect 10962 30679 11020 30685
rect 11054 30676 11060 30688
rect 11112 30676 11118 30728
rect 11422 30676 11428 30728
rect 11480 30676 11486 30728
rect 13078 30676 13084 30728
rect 13136 30676 13142 30728
rect 13265 30719 13323 30725
rect 13265 30685 13277 30719
rect 13311 30716 13323 30719
rect 14182 30716 14188 30728
rect 13311 30688 14188 30716
rect 13311 30685 13323 30688
rect 13265 30679 13323 30685
rect 12158 30608 12164 30660
rect 12216 30648 12222 30660
rect 13280 30648 13308 30679
rect 14182 30676 14188 30688
rect 14240 30676 14246 30728
rect 15010 30676 15016 30728
rect 15068 30716 15074 30728
rect 15488 30725 15516 30880
rect 17957 30855 18015 30861
rect 17957 30821 17969 30855
rect 18003 30852 18015 30855
rect 18003 30824 18736 30852
rect 18003 30821 18015 30824
rect 17957 30815 18015 30821
rect 16666 30784 16672 30796
rect 15580 30756 16672 30784
rect 15580 30728 15608 30756
rect 16666 30744 16672 30756
rect 16724 30744 16730 30796
rect 15197 30719 15255 30725
rect 15197 30716 15209 30719
rect 15068 30688 15209 30716
rect 15068 30676 15074 30688
rect 15197 30685 15209 30688
rect 15243 30685 15255 30719
rect 15197 30679 15255 30685
rect 15289 30719 15347 30725
rect 15289 30685 15301 30719
rect 15335 30685 15347 30719
rect 15289 30679 15347 30685
rect 15473 30719 15531 30725
rect 15473 30685 15485 30719
rect 15519 30685 15531 30719
rect 15473 30679 15531 30685
rect 12216 30620 13308 30648
rect 15304 30648 15332 30679
rect 15562 30676 15568 30728
rect 15620 30676 15626 30728
rect 15654 30676 15660 30728
rect 15712 30676 15718 30728
rect 17773 30719 17831 30725
rect 17773 30685 17785 30719
rect 17819 30685 17831 30719
rect 17773 30679 17831 30685
rect 17957 30719 18015 30725
rect 17957 30685 17969 30719
rect 18003 30716 18015 30719
rect 18049 30719 18107 30725
rect 18049 30716 18061 30719
rect 18003 30688 18061 30716
rect 18003 30685 18015 30688
rect 17957 30679 18015 30685
rect 18049 30685 18061 30688
rect 18095 30716 18107 30719
rect 18322 30716 18328 30728
rect 18095 30688 18328 30716
rect 18095 30685 18107 30688
rect 18049 30679 18107 30685
rect 15304 30620 17632 30648
rect 12216 30608 12222 30620
rect 7515 30552 8616 30580
rect 7515 30549 7527 30552
rect 7469 30543 7527 30549
rect 10318 30540 10324 30592
rect 10376 30580 10382 30592
rect 10594 30580 10600 30592
rect 10376 30552 10600 30580
rect 10376 30540 10382 30552
rect 10594 30540 10600 30552
rect 10652 30580 10658 30592
rect 10965 30583 11023 30589
rect 10965 30580 10977 30583
rect 10652 30552 10977 30580
rect 10652 30540 10658 30552
rect 10965 30549 10977 30552
rect 11011 30549 11023 30583
rect 10965 30543 11023 30549
rect 12894 30540 12900 30592
rect 12952 30580 12958 30592
rect 13262 30580 13268 30592
rect 12952 30552 13268 30580
rect 12952 30540 12958 30552
rect 13262 30540 13268 30552
rect 13320 30540 13326 30592
rect 15286 30540 15292 30592
rect 15344 30580 15350 30592
rect 16482 30580 16488 30592
rect 15344 30552 16488 30580
rect 15344 30540 15350 30552
rect 16482 30540 16488 30552
rect 16540 30540 16546 30592
rect 17604 30580 17632 30620
rect 17678 30608 17684 30660
rect 17736 30648 17742 30660
rect 17788 30648 17816 30679
rect 18322 30676 18328 30688
rect 18380 30676 18386 30728
rect 18233 30651 18291 30657
rect 18233 30648 18245 30651
rect 17736 30620 18245 30648
rect 17736 30608 17742 30620
rect 18233 30617 18245 30620
rect 18279 30617 18291 30651
rect 18233 30611 18291 30617
rect 18509 30651 18567 30657
rect 18509 30617 18521 30651
rect 18555 30648 18567 30651
rect 18598 30648 18604 30660
rect 18555 30620 18604 30648
rect 18555 30617 18567 30620
rect 18509 30611 18567 30617
rect 18598 30608 18604 30620
rect 18656 30608 18662 30660
rect 18708 30657 18736 30824
rect 22922 30812 22928 30864
rect 22980 30852 22986 30864
rect 27522 30852 27528 30864
rect 22980 30824 27528 30852
rect 22980 30812 22986 30824
rect 27522 30812 27528 30824
rect 27580 30812 27586 30864
rect 27706 30812 27712 30864
rect 27764 30812 27770 30864
rect 27798 30812 27804 30864
rect 27856 30812 27862 30864
rect 28350 30812 28356 30864
rect 28408 30852 28414 30864
rect 28902 30852 28908 30864
rect 28408 30824 28908 30852
rect 28408 30812 28414 30824
rect 28902 30812 28908 30824
rect 28960 30852 28966 30864
rect 30377 30855 30435 30861
rect 30377 30852 30389 30855
rect 28960 30824 30389 30852
rect 28960 30812 28966 30824
rect 30377 30821 30389 30824
rect 30423 30821 30435 30855
rect 30377 30815 30435 30821
rect 31312 30852 31340 30892
rect 33594 30880 33600 30932
rect 33652 30880 33658 30932
rect 34698 30920 34704 30932
rect 33704 30892 34704 30920
rect 33704 30852 33732 30892
rect 34698 30880 34704 30892
rect 34756 30920 34762 30932
rect 35161 30923 35219 30929
rect 35161 30920 35173 30923
rect 34756 30892 35173 30920
rect 34756 30880 34762 30892
rect 35161 30889 35173 30892
rect 35207 30889 35219 30923
rect 35161 30883 35219 30889
rect 35713 30923 35771 30929
rect 35713 30889 35725 30923
rect 35759 30920 35771 30923
rect 36354 30920 36360 30932
rect 35759 30892 36360 30920
rect 35759 30889 35771 30892
rect 35713 30883 35771 30889
rect 36354 30880 36360 30892
rect 36412 30880 36418 30932
rect 36909 30923 36967 30929
rect 36909 30889 36921 30923
rect 36955 30920 36967 30923
rect 37458 30920 37464 30932
rect 36955 30892 37464 30920
rect 36955 30889 36967 30892
rect 36909 30883 36967 30889
rect 37458 30880 37464 30892
rect 37516 30880 37522 30932
rect 38013 30923 38071 30929
rect 38013 30889 38025 30923
rect 38059 30920 38071 30923
rect 38286 30920 38292 30932
rect 38059 30892 38292 30920
rect 38059 30889 38071 30892
rect 38013 30883 38071 30889
rect 38286 30880 38292 30892
rect 38344 30880 38350 30932
rect 31312 30824 33732 30852
rect 19337 30787 19395 30793
rect 19337 30753 19349 30787
rect 19383 30784 19395 30787
rect 20438 30784 20444 30796
rect 19383 30756 20444 30784
rect 19383 30753 19395 30756
rect 19337 30747 19395 30753
rect 20438 30744 20444 30756
rect 20496 30744 20502 30796
rect 20806 30744 20812 30796
rect 20864 30744 20870 30796
rect 21082 30744 21088 30796
rect 21140 30744 21146 30796
rect 23860 30756 25912 30784
rect 21726 30676 21732 30728
rect 21784 30676 21790 30728
rect 23198 30676 23204 30728
rect 23256 30676 23262 30728
rect 23566 30676 23572 30728
rect 23624 30676 23630 30728
rect 23750 30676 23756 30728
rect 23808 30716 23814 30728
rect 23860 30725 23888 30756
rect 23845 30719 23903 30725
rect 23845 30716 23857 30719
rect 23808 30688 23857 30716
rect 23808 30676 23814 30688
rect 23845 30685 23857 30688
rect 23891 30685 23903 30719
rect 23845 30679 23903 30685
rect 23937 30719 23995 30725
rect 23937 30685 23949 30719
rect 23983 30685 23995 30719
rect 23937 30679 23995 30685
rect 18708 30651 18783 30657
rect 18708 30620 18737 30651
rect 18725 30617 18737 30620
rect 18771 30648 18783 30651
rect 19426 30648 19432 30660
rect 18771 30620 19432 30648
rect 18771 30617 18783 30620
rect 18725 30611 18783 30617
rect 19426 30608 19432 30620
rect 19484 30608 19490 30660
rect 21358 30648 21364 30660
rect 20378 30620 21364 30648
rect 21358 30608 21364 30620
rect 21416 30608 21422 30660
rect 21818 30648 21824 30660
rect 21560 30620 21824 30648
rect 17770 30580 17776 30592
rect 17604 30552 17776 30580
rect 17770 30540 17776 30552
rect 17828 30540 17834 30592
rect 20990 30540 20996 30592
rect 21048 30580 21054 30592
rect 21560 30580 21588 30620
rect 21818 30608 21824 30620
rect 21876 30648 21882 30660
rect 21913 30651 21971 30657
rect 21913 30648 21925 30651
rect 21876 30620 21925 30648
rect 21876 30608 21882 30620
rect 21913 30617 21925 30620
rect 21959 30617 21971 30651
rect 23952 30648 23980 30679
rect 25884 30660 25912 30756
rect 26510 30744 26516 30796
rect 26568 30784 26574 30796
rect 27724 30784 27752 30812
rect 28626 30784 28632 30796
rect 26568 30756 27752 30784
rect 27816 30756 28632 30784
rect 26568 30744 26574 30756
rect 26234 30676 26240 30728
rect 26292 30716 26298 30728
rect 26292 30688 26832 30716
rect 26292 30676 26298 30688
rect 21913 30611 21971 30617
rect 23492 30620 23980 30648
rect 24489 30651 24547 30657
rect 21048 30552 21588 30580
rect 21637 30583 21695 30589
rect 21048 30540 21054 30552
rect 21637 30549 21649 30583
rect 21683 30580 21695 30583
rect 22094 30580 22100 30592
rect 21683 30552 22100 30580
rect 21683 30549 21695 30552
rect 21637 30543 21695 30549
rect 22094 30540 22100 30552
rect 22152 30540 22158 30592
rect 23382 30540 23388 30592
rect 23440 30580 23446 30592
rect 23492 30589 23520 30620
rect 24489 30617 24501 30651
rect 24535 30617 24547 30651
rect 24489 30611 24547 30617
rect 23477 30583 23535 30589
rect 23477 30580 23489 30583
rect 23440 30552 23489 30580
rect 23440 30540 23446 30552
rect 23477 30549 23489 30552
rect 23523 30549 23535 30583
rect 23477 30543 23535 30549
rect 23842 30540 23848 30592
rect 23900 30580 23906 30592
rect 24504 30580 24532 30611
rect 25866 30608 25872 30660
rect 25924 30648 25930 30660
rect 26804 30657 26832 30688
rect 26878 30676 26884 30728
rect 26936 30676 26942 30728
rect 27540 30725 27568 30756
rect 27525 30719 27583 30725
rect 27525 30685 27537 30719
rect 27571 30685 27583 30719
rect 27525 30679 27583 30685
rect 27614 30676 27620 30728
rect 27672 30716 27678 30728
rect 27709 30719 27767 30725
rect 27709 30716 27721 30719
rect 27672 30688 27721 30716
rect 27672 30676 27678 30688
rect 27709 30685 27721 30688
rect 27755 30685 27767 30719
rect 27709 30679 27767 30685
rect 26605 30651 26663 30657
rect 26605 30648 26617 30651
rect 25924 30620 26617 30648
rect 25924 30608 25930 30620
rect 26605 30617 26617 30620
rect 26651 30617 26663 30651
rect 26605 30611 26663 30617
rect 26789 30651 26847 30657
rect 26789 30617 26801 30651
rect 26835 30648 26847 30651
rect 27816 30648 27844 30756
rect 28626 30744 28632 30756
rect 28684 30744 28690 30796
rect 30466 30744 30472 30796
rect 30524 30784 30530 30796
rect 30524 30756 31248 30784
rect 30524 30744 30530 30756
rect 31220 30728 31248 30756
rect 27890 30676 27896 30728
rect 27948 30716 27954 30728
rect 28721 30719 28779 30725
rect 28721 30716 28733 30719
rect 27948 30688 28733 30716
rect 27948 30676 27954 30688
rect 28721 30685 28733 30688
rect 28767 30685 28779 30719
rect 28721 30679 28779 30685
rect 26835 30620 27844 30648
rect 26835 30617 26847 30620
rect 26789 30611 26847 30617
rect 28166 30608 28172 30660
rect 28224 30648 28230 30660
rect 28353 30651 28411 30657
rect 28353 30648 28365 30651
rect 28224 30620 28365 30648
rect 28224 30608 28230 30620
rect 28353 30617 28365 30620
rect 28399 30617 28411 30651
rect 28353 30611 28411 30617
rect 28537 30651 28595 30657
rect 28537 30617 28549 30651
rect 28583 30648 28595 30651
rect 28626 30648 28632 30660
rect 28583 30620 28632 30648
rect 28583 30617 28595 30620
rect 28537 30611 28595 30617
rect 28626 30608 28632 30620
rect 28684 30608 28690 30660
rect 28184 30580 28212 30608
rect 23900 30552 28212 30580
rect 28736 30580 28764 30679
rect 28994 30676 29000 30728
rect 29052 30676 29058 30728
rect 29546 30676 29552 30728
rect 29604 30676 29610 30728
rect 30374 30676 30380 30728
rect 30432 30716 30438 30728
rect 30742 30716 30748 30728
rect 30432 30688 30748 30716
rect 30432 30676 30438 30688
rect 30742 30676 30748 30688
rect 30800 30716 30806 30728
rect 30837 30719 30895 30725
rect 30837 30716 30849 30719
rect 30800 30688 30849 30716
rect 30800 30676 30806 30688
rect 30837 30685 30849 30688
rect 30883 30685 30895 30719
rect 30837 30679 30895 30685
rect 31113 30719 31171 30725
rect 31113 30685 31125 30719
rect 31159 30685 31171 30719
rect 31113 30679 31171 30685
rect 30098 30608 30104 30660
rect 30156 30648 30162 30660
rect 30558 30648 30564 30660
rect 30156 30620 30564 30648
rect 30156 30608 30162 30620
rect 30558 30608 30564 30620
rect 30616 30648 30622 30660
rect 30653 30651 30711 30657
rect 30653 30648 30665 30651
rect 30616 30620 30665 30648
rect 30616 30608 30622 30620
rect 30653 30617 30665 30620
rect 30699 30617 30711 30651
rect 31128 30648 31156 30679
rect 31202 30676 31208 30728
rect 31260 30676 31266 30728
rect 31312 30725 31340 30824
rect 34606 30812 34612 30864
rect 34664 30852 34670 30864
rect 34977 30855 35035 30861
rect 34977 30852 34989 30855
rect 34664 30824 34989 30852
rect 34664 30812 34670 30824
rect 34977 30821 34989 30824
rect 35023 30821 35035 30855
rect 36078 30852 36084 30864
rect 34977 30815 35035 30821
rect 35176 30824 36084 30852
rect 32122 30784 32128 30796
rect 31496 30756 32128 30784
rect 31496 30725 31524 30756
rect 32122 30744 32128 30756
rect 32180 30784 32186 30796
rect 32674 30784 32680 30796
rect 32180 30756 32680 30784
rect 32180 30744 32186 30756
rect 32674 30744 32680 30756
rect 32732 30744 32738 30796
rect 33686 30744 33692 30796
rect 33744 30784 33750 30796
rect 35176 30784 35204 30824
rect 36078 30812 36084 30824
rect 36136 30852 36142 30864
rect 36814 30852 36820 30864
rect 36136 30824 36820 30852
rect 36136 30812 36142 30824
rect 36814 30812 36820 30824
rect 36872 30812 36878 30864
rect 36998 30812 37004 30864
rect 37056 30852 37062 30864
rect 38197 30855 38255 30861
rect 38197 30852 38209 30855
rect 37056 30824 38209 30852
rect 37056 30812 37062 30824
rect 38197 30821 38209 30824
rect 38243 30821 38255 30855
rect 38197 30815 38255 30821
rect 33744 30756 35204 30784
rect 33744 30744 33750 30756
rect 31297 30719 31355 30725
rect 31297 30685 31309 30719
rect 31343 30685 31355 30719
rect 31297 30679 31355 30685
rect 31481 30719 31539 30725
rect 31481 30685 31493 30719
rect 31527 30685 31539 30719
rect 31481 30679 31539 30685
rect 31570 30676 31576 30728
rect 31628 30676 31634 30728
rect 31757 30719 31815 30725
rect 31757 30685 31769 30719
rect 31803 30685 31815 30719
rect 31757 30679 31815 30685
rect 31662 30648 31668 30660
rect 31128 30620 31668 30648
rect 30653 30611 30711 30617
rect 31662 30608 31668 30620
rect 31720 30608 31726 30660
rect 28813 30583 28871 30589
rect 28813 30580 28825 30583
rect 28736 30552 28825 30580
rect 23900 30540 23906 30552
rect 28813 30549 28825 30552
rect 28859 30549 28871 30583
rect 28813 30543 28871 30549
rect 30193 30583 30251 30589
rect 30193 30549 30205 30583
rect 30239 30580 30251 30583
rect 30282 30580 30288 30592
rect 30239 30552 30288 30580
rect 30239 30549 30251 30552
rect 30193 30543 30251 30549
rect 30282 30540 30288 30552
rect 30340 30540 30346 30592
rect 31110 30540 31116 30592
rect 31168 30580 31174 30592
rect 31389 30583 31447 30589
rect 31389 30580 31401 30583
rect 31168 30552 31401 30580
rect 31168 30540 31174 30552
rect 31389 30549 31401 30552
rect 31435 30549 31447 30583
rect 31772 30580 31800 30679
rect 32030 30676 32036 30728
rect 32088 30716 32094 30728
rect 33781 30719 33839 30725
rect 33781 30716 33793 30719
rect 32088 30688 33793 30716
rect 32088 30676 32094 30688
rect 33781 30685 33793 30688
rect 33827 30685 33839 30719
rect 33781 30679 33839 30685
rect 33870 30676 33876 30728
rect 33928 30676 33934 30728
rect 34241 30719 34299 30725
rect 34241 30685 34253 30719
rect 34287 30716 34299 30719
rect 34330 30716 34336 30728
rect 34287 30688 34336 30716
rect 34287 30685 34299 30688
rect 34241 30679 34299 30685
rect 34330 30676 34336 30688
rect 34388 30676 34394 30728
rect 35176 30725 35204 30756
rect 35345 30787 35403 30793
rect 35345 30753 35357 30787
rect 35391 30784 35403 30787
rect 36262 30784 36268 30796
rect 35391 30756 36268 30784
rect 35391 30753 35403 30756
rect 35345 30747 35403 30753
rect 36262 30744 36268 30756
rect 36320 30784 36326 30796
rect 37550 30784 37556 30796
rect 36320 30756 37556 30784
rect 36320 30744 36326 30756
rect 35161 30719 35219 30725
rect 35161 30685 35173 30719
rect 35207 30685 35219 30719
rect 35713 30719 35771 30725
rect 35713 30716 35725 30719
rect 35161 30679 35219 30685
rect 35268 30688 35725 30716
rect 32306 30608 32312 30660
rect 32364 30648 32370 30660
rect 32582 30648 32588 30660
rect 32364 30620 32588 30648
rect 32364 30608 32370 30620
rect 32582 30608 32588 30620
rect 32640 30608 32646 30660
rect 33318 30608 33324 30660
rect 33376 30648 33382 30660
rect 33965 30651 34023 30657
rect 33965 30648 33977 30651
rect 33376 30620 33977 30648
rect 33376 30608 33382 30620
rect 33965 30617 33977 30620
rect 34011 30617 34023 30651
rect 33965 30611 34023 30617
rect 34103 30651 34161 30657
rect 34103 30617 34115 30651
rect 34149 30648 34161 30651
rect 34348 30648 34376 30676
rect 35268 30648 35296 30688
rect 35713 30685 35725 30688
rect 35759 30685 35771 30719
rect 35713 30679 35771 30685
rect 35897 30719 35955 30725
rect 35897 30685 35909 30719
rect 35943 30685 35955 30719
rect 35897 30679 35955 30685
rect 34149 30620 34284 30648
rect 34348 30620 35296 30648
rect 35621 30651 35679 30657
rect 34149 30617 34161 30620
rect 34103 30611 34161 30617
rect 34256 30592 34284 30620
rect 35621 30617 35633 30651
rect 35667 30617 35679 30651
rect 35912 30648 35940 30679
rect 36170 30676 36176 30728
rect 36228 30716 36234 30728
rect 36633 30719 36691 30725
rect 36633 30716 36645 30719
rect 36228 30688 36645 30716
rect 36228 30676 36234 30688
rect 36633 30685 36645 30688
rect 36679 30685 36691 30719
rect 36633 30679 36691 30685
rect 36814 30676 36820 30728
rect 36872 30676 36878 30728
rect 37108 30725 37136 30756
rect 37550 30744 37556 30756
rect 37608 30784 37614 30796
rect 37737 30787 37795 30793
rect 37737 30784 37749 30787
rect 37608 30756 37749 30784
rect 37608 30744 37614 30756
rect 37737 30753 37749 30756
rect 37783 30753 37795 30787
rect 37737 30747 37795 30753
rect 36909 30719 36967 30725
rect 36909 30685 36921 30719
rect 36955 30685 36967 30719
rect 36909 30679 36967 30685
rect 37093 30719 37151 30725
rect 37093 30685 37105 30719
rect 37139 30685 37151 30719
rect 37093 30679 37151 30685
rect 36924 30648 36952 30679
rect 37366 30676 37372 30728
rect 37424 30676 37430 30728
rect 37642 30676 37648 30728
rect 37700 30716 37706 30728
rect 37700 30688 38148 30716
rect 37700 30676 37706 30688
rect 38120 30660 38148 30688
rect 38286 30676 38292 30728
rect 38344 30716 38350 30728
rect 38473 30719 38531 30725
rect 38473 30716 38485 30719
rect 38344 30688 38485 30716
rect 38344 30676 38350 30688
rect 38473 30685 38485 30688
rect 38519 30685 38531 30719
rect 38473 30679 38531 30685
rect 35912 30620 36952 30648
rect 35621 30611 35679 30617
rect 33594 30580 33600 30592
rect 31772 30552 33600 30580
rect 31389 30543 31447 30549
rect 33594 30540 33600 30552
rect 33652 30540 33658 30592
rect 34238 30540 34244 30592
rect 34296 30540 34302 30592
rect 35636 30580 35664 30611
rect 36170 30580 36176 30592
rect 35636 30552 36176 30580
rect 36170 30540 36176 30552
rect 36228 30540 36234 30592
rect 36648 30589 36676 30620
rect 37458 30608 37464 30660
rect 37516 30648 37522 30660
rect 37854 30651 37912 30657
rect 37854 30648 37866 30651
rect 37516 30620 37866 30648
rect 37516 30608 37522 30620
rect 37854 30617 37866 30620
rect 37900 30617 37912 30651
rect 37854 30611 37912 30617
rect 38102 30608 38108 30660
rect 38160 30648 38166 30660
rect 38381 30651 38439 30657
rect 38381 30648 38393 30651
rect 38160 30620 38393 30648
rect 38160 30608 38166 30620
rect 38381 30617 38393 30620
rect 38427 30617 38439 30651
rect 38381 30611 38439 30617
rect 38746 30608 38752 30660
rect 38804 30648 38810 30660
rect 38933 30651 38991 30657
rect 38933 30648 38945 30651
rect 38804 30620 38945 30648
rect 38804 30608 38810 30620
rect 38933 30617 38945 30620
rect 38979 30648 38991 30651
rect 39022 30648 39028 30660
rect 38979 30620 39028 30648
rect 38979 30617 38991 30620
rect 38933 30611 38991 30617
rect 39022 30608 39028 30620
rect 39080 30608 39086 30660
rect 36633 30583 36691 30589
rect 36633 30549 36645 30583
rect 36679 30580 36691 30583
rect 36722 30580 36728 30592
rect 36679 30552 36728 30580
rect 36679 30549 36691 30552
rect 36633 30543 36691 30549
rect 36722 30540 36728 30552
rect 36780 30540 36786 30592
rect 37642 30540 37648 30592
rect 37700 30540 37706 30592
rect 1104 30490 40572 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 40572 30490
rect 1104 30416 40572 30438
rect 1578 30336 1584 30388
rect 1636 30376 1642 30388
rect 3053 30379 3111 30385
rect 3053 30376 3065 30379
rect 1636 30348 3065 30376
rect 1636 30336 1642 30348
rect 3053 30345 3065 30348
rect 3099 30345 3111 30379
rect 3053 30339 3111 30345
rect 4525 30379 4583 30385
rect 4525 30345 4537 30379
rect 4571 30376 4583 30379
rect 4571 30348 4936 30376
rect 4571 30345 4583 30348
rect 4525 30339 4583 30345
rect 4908 30320 4936 30348
rect 7834 30336 7840 30388
rect 7892 30376 7898 30388
rect 8570 30376 8576 30388
rect 7892 30348 8576 30376
rect 7892 30336 7898 30348
rect 8570 30336 8576 30348
rect 8628 30336 8634 30388
rect 10597 30379 10655 30385
rect 10597 30345 10609 30379
rect 10643 30376 10655 30379
rect 10686 30376 10692 30388
rect 10643 30348 10692 30376
rect 10643 30345 10655 30348
rect 10597 30339 10655 30345
rect 10686 30336 10692 30348
rect 10744 30336 10750 30388
rect 13078 30336 13084 30388
rect 13136 30376 13142 30388
rect 14274 30376 14280 30388
rect 13136 30348 14280 30376
rect 13136 30336 13142 30348
rect 14274 30336 14280 30348
rect 14332 30376 14338 30388
rect 14461 30379 14519 30385
rect 14461 30376 14473 30379
rect 14332 30348 14473 30376
rect 14332 30336 14338 30348
rect 14461 30345 14473 30348
rect 14507 30345 14519 30379
rect 14461 30339 14519 30345
rect 15580 30348 16528 30376
rect 2685 30311 2743 30317
rect 2685 30277 2697 30311
rect 2731 30308 2743 30311
rect 3326 30308 3332 30320
rect 2731 30280 3332 30308
rect 2731 30277 2743 30280
rect 2685 30271 2743 30277
rect 3326 30268 3332 30280
rect 3384 30268 3390 30320
rect 4798 30308 4804 30320
rect 4448 30280 4804 30308
rect 842 30200 848 30252
rect 900 30240 906 30252
rect 1489 30243 1547 30249
rect 1489 30240 1501 30243
rect 900 30212 1501 30240
rect 900 30200 906 30212
rect 1489 30209 1501 30212
rect 1535 30209 1547 30243
rect 1489 30203 1547 30209
rect 2866 30200 2872 30252
rect 2924 30200 2930 30252
rect 3145 30243 3203 30249
rect 3145 30209 3157 30243
rect 3191 30240 3203 30243
rect 4448 30240 4476 30280
rect 4798 30268 4804 30280
rect 4856 30268 4862 30320
rect 4890 30268 4896 30320
rect 4948 30268 4954 30320
rect 9398 30268 9404 30320
rect 9456 30308 9462 30320
rect 11330 30308 11336 30320
rect 9456 30280 11336 30308
rect 9456 30268 9462 30280
rect 11330 30268 11336 30280
rect 11388 30308 11394 30320
rect 11606 30308 11612 30320
rect 11388 30280 11612 30308
rect 11388 30268 11394 30280
rect 11606 30268 11612 30280
rect 11664 30268 11670 30320
rect 11698 30268 11704 30320
rect 11756 30308 11762 30320
rect 12345 30311 12403 30317
rect 11756 30280 12112 30308
rect 11756 30268 11762 30280
rect 3191 30212 4476 30240
rect 3191 30209 3203 30212
rect 3145 30203 3203 30209
rect 7374 30200 7380 30252
rect 7432 30200 7438 30252
rect 10870 30200 10876 30252
rect 10928 30200 10934 30252
rect 12084 30249 12112 30280
rect 12345 30277 12357 30311
rect 12391 30308 12403 30311
rect 12391 30280 13124 30308
rect 12391 30277 12403 30280
rect 12345 30271 12403 30277
rect 12043 30243 12112 30249
rect 12043 30209 12055 30243
rect 12089 30240 12112 30243
rect 12089 30212 12204 30240
rect 12089 30209 12101 30212
rect 12043 30203 12101 30209
rect 4614 30132 4620 30184
rect 4672 30132 4678 30184
rect 4798 30132 4804 30184
rect 4856 30132 4862 30184
rect 4890 30132 4896 30184
rect 4948 30172 4954 30184
rect 5258 30172 5264 30184
rect 4948 30144 5264 30172
rect 4948 30132 4954 30144
rect 5258 30132 5264 30144
rect 5316 30172 5322 30184
rect 9858 30172 9864 30184
rect 5316 30144 9864 30172
rect 5316 30132 5322 30144
rect 9858 30132 9864 30144
rect 9916 30132 9922 30184
rect 11882 30132 11888 30184
rect 11940 30132 11946 30184
rect 12176 30172 12204 30212
rect 12434 30200 12440 30252
rect 12492 30200 12498 30252
rect 12897 30243 12955 30249
rect 12897 30240 12909 30243
rect 12543 30212 12909 30240
rect 12543 30172 12571 30212
rect 12897 30209 12909 30212
rect 12943 30209 12955 30243
rect 12897 30203 12955 30209
rect 12176 30144 12571 30172
rect 12713 30175 12771 30181
rect 12713 30141 12725 30175
rect 12759 30141 12771 30175
rect 12713 30135 12771 30141
rect 1765 30107 1823 30113
rect 1765 30073 1777 30107
rect 1811 30104 1823 30107
rect 5902 30104 5908 30116
rect 1811 30076 5908 30104
rect 1811 30073 1823 30076
rect 1765 30067 1823 30073
rect 5902 30064 5908 30076
rect 5960 30064 5966 30116
rect 6178 30064 6184 30116
rect 6236 30104 6242 30116
rect 7834 30104 7840 30116
rect 6236 30076 7840 30104
rect 6236 30064 6242 30076
rect 7834 30064 7840 30076
rect 7892 30064 7898 30116
rect 11974 30064 11980 30116
rect 12032 30104 12038 30116
rect 12526 30104 12532 30116
rect 12032 30076 12532 30104
rect 12032 30064 12038 30076
rect 12526 30064 12532 30076
rect 12584 30064 12590 30116
rect 12728 30104 12756 30135
rect 12894 30104 12900 30116
rect 12728 30076 12900 30104
rect 12894 30064 12900 30076
rect 12952 30064 12958 30116
rect 13096 30104 13124 30280
rect 13262 30268 13268 30320
rect 13320 30308 13326 30320
rect 15580 30308 15608 30348
rect 13320 30280 13952 30308
rect 13320 30268 13326 30280
rect 13924 30249 13952 30280
rect 15212 30280 15608 30308
rect 13449 30243 13507 30249
rect 13449 30209 13461 30243
rect 13495 30240 13507 30243
rect 13725 30243 13783 30249
rect 13725 30240 13737 30243
rect 13495 30212 13737 30240
rect 13495 30209 13507 30212
rect 13449 30203 13507 30209
rect 13725 30209 13737 30212
rect 13771 30209 13783 30243
rect 13725 30203 13783 30209
rect 13909 30243 13967 30249
rect 13909 30209 13921 30243
rect 13955 30209 13967 30243
rect 13909 30203 13967 30209
rect 14001 30243 14059 30249
rect 14001 30209 14013 30243
rect 14047 30240 14059 30243
rect 14182 30240 14188 30252
rect 14047 30212 14188 30240
rect 14047 30209 14059 30212
rect 14001 30203 14059 30209
rect 14182 30200 14188 30212
rect 14240 30200 14246 30252
rect 14277 30243 14335 30249
rect 14277 30209 14289 30243
rect 14323 30240 14335 30243
rect 14366 30240 14372 30252
rect 14323 30212 14372 30240
rect 14323 30209 14335 30212
rect 14277 30203 14335 30209
rect 14366 30200 14372 30212
rect 14424 30200 14430 30252
rect 14642 30200 14648 30252
rect 14700 30200 14706 30252
rect 14921 30243 14979 30249
rect 14921 30209 14933 30243
rect 14967 30240 14979 30243
rect 15010 30240 15016 30252
rect 14967 30212 15016 30240
rect 14967 30209 14979 30212
rect 14921 30203 14979 30209
rect 15010 30200 15016 30212
rect 15068 30200 15074 30252
rect 15102 30200 15108 30252
rect 15160 30240 15166 30252
rect 15212 30249 15240 30280
rect 15654 30268 15660 30320
rect 15712 30308 15718 30320
rect 16500 30308 16528 30348
rect 18230 30336 18236 30388
rect 18288 30376 18294 30388
rect 18325 30379 18383 30385
rect 18325 30376 18337 30379
rect 18288 30348 18337 30376
rect 18288 30336 18294 30348
rect 18325 30345 18337 30348
rect 18371 30345 18383 30379
rect 23290 30376 23296 30388
rect 18325 30339 18383 30345
rect 23216 30348 23296 30376
rect 21174 30308 21180 30320
rect 15712 30280 16441 30308
rect 16500 30280 21180 30308
rect 15712 30268 15718 30280
rect 15197 30243 15255 30249
rect 15197 30240 15209 30243
rect 15160 30212 15209 30240
rect 15160 30200 15166 30212
rect 15197 30209 15209 30212
rect 15243 30209 15255 30243
rect 15197 30203 15255 30209
rect 15381 30243 15439 30249
rect 15381 30209 15393 30243
rect 15427 30209 15439 30243
rect 15381 30203 15439 30209
rect 13170 30132 13176 30184
rect 13228 30172 13234 30184
rect 13357 30175 13415 30181
rect 13357 30172 13369 30175
rect 13228 30144 13369 30172
rect 13228 30132 13234 30144
rect 13357 30141 13369 30144
rect 13403 30141 13415 30175
rect 15396 30172 15424 30203
rect 15562 30200 15568 30252
rect 15620 30240 15626 30252
rect 15948 30249 15976 30280
rect 16413 30255 16441 30280
rect 21174 30268 21180 30280
rect 21232 30268 21238 30320
rect 22370 30268 22376 30320
rect 22428 30308 22434 30320
rect 23216 30317 23244 30348
rect 23290 30336 23296 30348
rect 23348 30376 23354 30388
rect 23348 30348 25452 30376
rect 23348 30336 23354 30348
rect 23201 30311 23259 30317
rect 23201 30308 23213 30311
rect 22428 30280 23213 30308
rect 22428 30268 22434 30280
rect 23201 30277 23213 30280
rect 23247 30277 23259 30311
rect 24210 30308 24216 30320
rect 23201 30271 23259 30277
rect 23308 30280 24216 30308
rect 15749 30243 15807 30249
rect 15749 30240 15761 30243
rect 15620 30212 15761 30240
rect 15620 30200 15626 30212
rect 15749 30209 15761 30212
rect 15795 30209 15807 30243
rect 15749 30203 15807 30209
rect 15933 30243 15991 30249
rect 15933 30209 15945 30243
rect 15979 30209 15991 30243
rect 15933 30203 15991 30209
rect 16022 30200 16028 30252
rect 16080 30200 16086 30252
rect 16209 30243 16267 30249
rect 16209 30209 16221 30243
rect 16255 30209 16267 30243
rect 16209 30203 16267 30209
rect 15470 30172 15476 30184
rect 13357 30135 13415 30141
rect 13464 30144 15148 30172
rect 15396 30144 15476 30172
rect 13464 30104 13492 30144
rect 15013 30107 15071 30113
rect 15013 30104 15025 30107
rect 13096 30076 13492 30104
rect 13556 30076 15025 30104
rect 4062 29996 4068 30048
rect 4120 30036 4126 30048
rect 4157 30039 4215 30045
rect 4157 30036 4169 30039
rect 4120 30008 4169 30036
rect 4120 29996 4126 30008
rect 4157 30005 4169 30008
rect 4203 30005 4215 30039
rect 4157 29999 4215 30005
rect 7469 30039 7527 30045
rect 7469 30005 7481 30039
rect 7515 30036 7527 30039
rect 7650 30036 7656 30048
rect 7515 30008 7656 30036
rect 7515 30005 7527 30008
rect 7469 29999 7527 30005
rect 7650 29996 7656 30008
rect 7708 29996 7714 30048
rect 9766 29996 9772 30048
rect 9824 30036 9830 30048
rect 12342 30036 12348 30048
rect 9824 30008 12348 30036
rect 9824 29996 9830 30008
rect 12342 29996 12348 30008
rect 12400 30036 12406 30048
rect 13556 30036 13584 30076
rect 15013 30073 15025 30076
rect 15059 30073 15071 30107
rect 15120 30104 15148 30144
rect 15470 30132 15476 30144
rect 15528 30172 15534 30184
rect 16224 30172 16252 30203
rect 16298 30200 16304 30252
rect 16356 30200 16362 30252
rect 16413 30249 16471 30255
rect 16413 30215 16425 30249
rect 16459 30246 16471 30249
rect 16459 30240 16528 30246
rect 16758 30240 16764 30252
rect 16459 30218 16764 30240
rect 16459 30215 16471 30218
rect 16413 30209 16471 30215
rect 16500 30212 16764 30218
rect 16758 30200 16764 30212
rect 16816 30200 16822 30252
rect 16945 30243 17003 30249
rect 16945 30209 16957 30243
rect 16991 30240 17003 30243
rect 17126 30240 17132 30252
rect 16991 30212 17132 30240
rect 16991 30209 17003 30212
rect 16945 30203 17003 30209
rect 17126 30200 17132 30212
rect 17184 30200 17190 30252
rect 18414 30200 18420 30252
rect 18472 30240 18478 30252
rect 18693 30243 18751 30249
rect 18693 30240 18705 30243
rect 18472 30212 18705 30240
rect 18472 30200 18478 30212
rect 18693 30209 18705 30212
rect 18739 30209 18751 30243
rect 18693 30203 18751 30209
rect 22094 30200 22100 30252
rect 22152 30240 22158 30252
rect 23106 30249 23112 30252
rect 23063 30243 23112 30249
rect 23063 30240 23075 30243
rect 22152 30212 23075 30240
rect 22152 30200 22158 30212
rect 23063 30209 23075 30212
rect 23109 30209 23112 30243
rect 23063 30203 23112 30209
rect 23106 30200 23112 30203
rect 23164 30200 23170 30252
rect 23308 30249 23336 30280
rect 24210 30268 24216 30280
rect 24268 30268 24274 30320
rect 23293 30243 23351 30249
rect 23293 30209 23305 30243
rect 23339 30209 23351 30243
rect 23293 30203 23351 30209
rect 23382 30200 23388 30252
rect 23440 30249 23446 30252
rect 23440 30243 23479 30249
rect 23467 30209 23479 30243
rect 23440 30203 23479 30209
rect 23569 30243 23627 30249
rect 23569 30209 23581 30243
rect 23615 30240 23627 30243
rect 23658 30240 23664 30252
rect 23615 30212 23664 30240
rect 23615 30209 23627 30212
rect 23569 30203 23627 30209
rect 23440 30200 23446 30203
rect 23658 30200 23664 30212
rect 23716 30200 23722 30252
rect 25424 30240 25452 30348
rect 27522 30336 27528 30388
rect 27580 30376 27586 30388
rect 29270 30376 29276 30388
rect 27580 30348 29276 30376
rect 27580 30336 27586 30348
rect 29270 30336 29276 30348
rect 29328 30336 29334 30388
rect 29914 30336 29920 30388
rect 29972 30376 29978 30388
rect 29972 30348 32260 30376
rect 29972 30336 29978 30348
rect 25866 30268 25872 30320
rect 25924 30268 25930 30320
rect 28074 30308 28080 30320
rect 26436 30280 28080 30308
rect 26436 30252 26464 30280
rect 28074 30268 28080 30280
rect 28132 30268 28138 30320
rect 28902 30268 28908 30320
rect 28960 30268 28966 30320
rect 30653 30311 30711 30317
rect 30653 30277 30665 30311
rect 30699 30308 30711 30311
rect 31021 30311 31079 30317
rect 31021 30308 31033 30311
rect 30699 30280 31033 30308
rect 30699 30277 30711 30280
rect 30653 30271 30711 30277
rect 31021 30277 31033 30280
rect 31067 30277 31079 30311
rect 31021 30271 31079 30277
rect 31649 30311 31707 30317
rect 31649 30277 31661 30311
rect 31695 30308 31707 30311
rect 31754 30308 31760 30320
rect 31695 30280 31760 30308
rect 31695 30277 31707 30280
rect 31649 30271 31707 30277
rect 31754 30268 31760 30280
rect 31812 30268 31818 30320
rect 31849 30311 31907 30317
rect 31849 30277 31861 30311
rect 31895 30308 31907 30311
rect 31938 30308 31944 30320
rect 31895 30280 31944 30308
rect 31895 30277 31907 30280
rect 31849 30271 31907 30277
rect 31938 30268 31944 30280
rect 31996 30268 32002 30320
rect 26418 30240 26424 30252
rect 25424 30212 26424 30240
rect 26418 30200 26424 30212
rect 26476 30200 26482 30252
rect 26513 30243 26571 30249
rect 26513 30209 26525 30243
rect 26559 30209 26571 30243
rect 26513 30203 26571 30209
rect 16669 30175 16727 30181
rect 15528 30144 16344 30172
rect 15528 30132 15534 30144
rect 16316 30104 16344 30144
rect 16669 30141 16681 30175
rect 16715 30172 16727 30175
rect 17678 30172 17684 30184
rect 16715 30144 17684 30172
rect 16715 30141 16727 30144
rect 16669 30135 16727 30141
rect 17678 30132 17684 30144
rect 17736 30132 17742 30184
rect 18598 30132 18604 30184
rect 18656 30132 18662 30184
rect 21726 30132 21732 30184
rect 21784 30172 21790 30184
rect 24486 30172 24492 30184
rect 21784 30144 24492 30172
rect 21784 30132 21790 30144
rect 24486 30132 24492 30144
rect 24544 30132 24550 30184
rect 24670 30132 24676 30184
rect 24728 30172 24734 30184
rect 25501 30175 25559 30181
rect 25501 30172 25513 30175
rect 24728 30144 25513 30172
rect 24728 30132 24734 30144
rect 25501 30141 25513 30144
rect 25547 30172 25559 30175
rect 25590 30172 25596 30184
rect 25547 30144 25596 30172
rect 25547 30141 25559 30144
rect 25501 30135 25559 30141
rect 25590 30132 25596 30144
rect 25648 30172 25654 30184
rect 26050 30172 26056 30184
rect 25648 30144 26056 30172
rect 25648 30132 25654 30144
rect 26050 30132 26056 30144
rect 26108 30172 26114 30184
rect 26234 30172 26240 30184
rect 26108 30144 26240 30172
rect 26108 30132 26114 30144
rect 26234 30132 26240 30144
rect 26292 30132 26298 30184
rect 26528 30172 26556 30203
rect 30282 30200 30288 30252
rect 30340 30200 30346 30252
rect 30466 30249 30472 30252
rect 30443 30243 30472 30249
rect 30443 30209 30455 30243
rect 30443 30203 30472 30209
rect 30466 30200 30472 30203
rect 30524 30200 30530 30252
rect 30558 30200 30564 30252
rect 30616 30200 30622 30252
rect 30745 30243 30803 30249
rect 30745 30209 30757 30243
rect 30791 30240 30803 30243
rect 31110 30240 31116 30252
rect 30791 30212 31116 30240
rect 30791 30209 30803 30212
rect 30745 30203 30803 30209
rect 31110 30200 31116 30212
rect 31168 30200 31174 30252
rect 31205 30243 31263 30249
rect 31205 30209 31217 30243
rect 31251 30209 31263 30243
rect 31205 30203 31263 30209
rect 26878 30172 26884 30184
rect 26528 30144 26884 30172
rect 26878 30132 26884 30144
rect 26936 30172 26942 30184
rect 28445 30175 28503 30181
rect 28445 30172 28457 30175
rect 26936 30144 28457 30172
rect 26936 30132 26942 30144
rect 28445 30141 28457 30144
rect 28491 30172 28503 30175
rect 29546 30172 29552 30184
rect 28491 30144 29552 30172
rect 28491 30141 28503 30144
rect 28445 30135 28503 30141
rect 29546 30132 29552 30144
rect 29604 30132 29610 30184
rect 29917 30175 29975 30181
rect 29917 30141 29929 30175
rect 29963 30172 29975 30175
rect 29963 30144 30144 30172
rect 29963 30141 29975 30144
rect 29917 30135 29975 30141
rect 16942 30104 16948 30116
rect 15120 30076 16160 30104
rect 16316 30076 16948 30104
rect 15013 30067 15071 30073
rect 12400 30008 13584 30036
rect 14185 30039 14243 30045
rect 12400 29996 12406 30008
rect 14185 30005 14197 30039
rect 14231 30036 14243 30039
rect 14274 30036 14280 30048
rect 14231 30008 14280 30036
rect 14231 30005 14243 30008
rect 14185 29999 14243 30005
rect 14274 29996 14280 30008
rect 14332 29996 14338 30048
rect 15562 29996 15568 30048
rect 15620 30036 15626 30048
rect 15930 30036 15936 30048
rect 15620 30008 15936 30036
rect 15620 29996 15626 30008
rect 15930 29996 15936 30008
rect 15988 29996 15994 30048
rect 16022 29996 16028 30048
rect 16080 29996 16086 30048
rect 16132 30036 16160 30076
rect 16942 30064 16948 30076
rect 17000 30064 17006 30116
rect 18233 30107 18291 30113
rect 18233 30073 18245 30107
rect 18279 30104 18291 30107
rect 18690 30104 18696 30116
rect 18279 30076 18696 30104
rect 18279 30073 18291 30076
rect 18233 30067 18291 30073
rect 16574 30036 16580 30048
rect 16132 30008 16580 30036
rect 16574 29996 16580 30008
rect 16632 29996 16638 30048
rect 16758 29996 16764 30048
rect 16816 29996 16822 30048
rect 17034 29996 17040 30048
rect 17092 30036 17098 30048
rect 18616 30045 18644 30076
rect 18690 30064 18696 30076
rect 18748 30104 18754 30116
rect 25774 30104 25780 30116
rect 18748 30076 25780 30104
rect 18748 30064 18754 30076
rect 25774 30064 25780 30076
rect 25832 30064 25838 30116
rect 25958 30064 25964 30116
rect 26016 30104 26022 30116
rect 26329 30107 26387 30113
rect 26329 30104 26341 30107
rect 26016 30076 26341 30104
rect 26016 30064 26022 30076
rect 26329 30073 26341 30076
rect 26375 30073 26387 30107
rect 30116 30104 30144 30144
rect 30190 30132 30196 30184
rect 30248 30132 30254 30184
rect 31220 30172 31248 30203
rect 31294 30200 31300 30252
rect 31352 30240 31358 30252
rect 31389 30243 31447 30249
rect 31389 30240 31401 30243
rect 31352 30212 31401 30240
rect 31352 30200 31358 30212
rect 31389 30209 31401 30212
rect 31435 30209 31447 30243
rect 31389 30203 31447 30209
rect 31496 30212 31984 30240
rect 31496 30172 31524 30212
rect 31772 30184 31800 30212
rect 31220 30144 31524 30172
rect 31754 30132 31760 30184
rect 31812 30132 31818 30184
rect 31956 30172 31984 30212
rect 32122 30200 32128 30252
rect 32180 30200 32186 30252
rect 32232 30240 32260 30348
rect 32674 30336 32680 30388
rect 32732 30376 32738 30388
rect 36354 30376 36360 30388
rect 32732 30348 36360 30376
rect 32732 30336 32738 30348
rect 36354 30336 36360 30348
rect 36412 30336 36418 30388
rect 36538 30336 36544 30388
rect 36596 30376 36602 30388
rect 37918 30376 37924 30388
rect 36596 30348 37924 30376
rect 36596 30336 36602 30348
rect 37918 30336 37924 30348
rect 37976 30336 37982 30388
rect 38856 30348 39804 30376
rect 33686 30268 33692 30320
rect 33744 30308 33750 30320
rect 33781 30311 33839 30317
rect 33781 30308 33793 30311
rect 33744 30280 33793 30308
rect 33744 30268 33750 30280
rect 33781 30277 33793 30280
rect 33827 30277 33839 30311
rect 38013 30311 38071 30317
rect 38013 30308 38025 30311
rect 33781 30271 33839 30277
rect 37568 30280 38025 30308
rect 37568 30252 37596 30280
rect 38013 30277 38025 30280
rect 38059 30277 38071 30311
rect 38856 30308 38884 30348
rect 38013 30271 38071 30277
rect 38120 30280 38884 30308
rect 32306 30240 32312 30252
rect 32232 30212 32312 30240
rect 32306 30200 32312 30212
rect 32364 30240 32370 30252
rect 32401 30243 32459 30249
rect 32401 30240 32413 30243
rect 32364 30212 32413 30240
rect 32364 30200 32370 30212
rect 32401 30209 32413 30212
rect 32447 30209 32459 30243
rect 32401 30203 32459 30209
rect 32493 30243 32551 30249
rect 32493 30209 32505 30243
rect 32539 30240 32551 30243
rect 33134 30240 33140 30252
rect 32539 30212 33140 30240
rect 32539 30209 32551 30212
rect 32493 30203 32551 30209
rect 33134 30200 33140 30212
rect 33192 30200 33198 30252
rect 34425 30243 34483 30249
rect 34425 30240 34437 30243
rect 33796 30212 34437 30240
rect 32217 30175 32275 30181
rect 32217 30172 32229 30175
rect 31956 30144 32229 30172
rect 32217 30141 32229 30144
rect 32263 30141 32275 30175
rect 32217 30135 32275 30141
rect 30929 30107 30987 30113
rect 30929 30104 30941 30107
rect 30116 30076 30941 30104
rect 26329 30067 26387 30073
rect 30929 30073 30941 30076
rect 30975 30073 30987 30107
rect 30929 30067 30987 30073
rect 31386 30064 31392 30116
rect 31444 30104 31450 30116
rect 31481 30107 31539 30113
rect 31481 30104 31493 30107
rect 31444 30076 31493 30104
rect 31444 30064 31450 30076
rect 31481 30073 31493 30076
rect 31527 30073 31539 30107
rect 31481 30067 31539 30073
rect 32030 30064 32036 30116
rect 32088 30104 32094 30116
rect 32125 30107 32183 30113
rect 32125 30104 32137 30107
rect 32088 30076 32137 30104
rect 32088 30064 32094 30076
rect 32125 30073 32137 30076
rect 32171 30073 32183 30107
rect 32125 30067 32183 30073
rect 33410 30064 33416 30116
rect 33468 30064 33474 30116
rect 17129 30039 17187 30045
rect 17129 30036 17141 30039
rect 17092 30008 17141 30036
rect 17092 29996 17098 30008
rect 17129 30005 17141 30008
rect 17175 30005 17187 30039
rect 17129 29999 17187 30005
rect 18601 30039 18659 30045
rect 18601 30005 18613 30039
rect 18647 30005 18659 30039
rect 18601 29999 18659 30005
rect 22925 30039 22983 30045
rect 22925 30005 22937 30039
rect 22971 30036 22983 30039
rect 23382 30036 23388 30048
rect 22971 30008 23388 30036
rect 22971 30005 22983 30008
rect 22925 29999 22983 30005
rect 23382 29996 23388 30008
rect 23440 29996 23446 30048
rect 24210 29996 24216 30048
rect 24268 30036 24274 30048
rect 25038 30036 25044 30048
rect 24268 30008 25044 30036
rect 24268 29996 24274 30008
rect 25038 29996 25044 30008
rect 25096 29996 25102 30048
rect 25406 29996 25412 30048
rect 25464 30036 25470 30048
rect 25869 30039 25927 30045
rect 25869 30036 25881 30039
rect 25464 30008 25881 30036
rect 25464 29996 25470 30008
rect 25869 30005 25881 30008
rect 25915 30005 25927 30039
rect 25869 29999 25927 30005
rect 26053 30039 26111 30045
rect 26053 30005 26065 30039
rect 26099 30036 26111 30039
rect 26234 30036 26240 30048
rect 26099 30008 26240 30036
rect 26099 30005 26111 30008
rect 26053 29999 26111 30005
rect 26234 29996 26240 30008
rect 26292 29996 26298 30048
rect 26970 29996 26976 30048
rect 27028 30036 27034 30048
rect 31570 30036 31576 30048
rect 27028 30008 31576 30036
rect 27028 29996 27034 30008
rect 31570 29996 31576 30008
rect 31628 29996 31634 30048
rect 31662 29996 31668 30048
rect 31720 29996 31726 30048
rect 32585 30039 32643 30045
rect 32585 30005 32597 30039
rect 32631 30036 32643 30039
rect 32674 30036 32680 30048
rect 32631 30008 32680 30036
rect 32631 30005 32643 30008
rect 32585 29999 32643 30005
rect 32674 29996 32680 30008
rect 32732 29996 32738 30048
rect 33594 29996 33600 30048
rect 33652 30036 33658 30048
rect 33796 30045 33824 30212
rect 34425 30209 34437 30212
rect 34471 30240 34483 30243
rect 34471 30212 34560 30240
rect 34471 30209 34483 30212
rect 34425 30203 34483 30209
rect 34054 30132 34060 30184
rect 34112 30172 34118 30184
rect 34241 30175 34299 30181
rect 34241 30172 34253 30175
rect 34112 30144 34253 30172
rect 34112 30132 34118 30144
rect 34241 30141 34253 30144
rect 34287 30141 34299 30175
rect 34241 30135 34299 30141
rect 34146 30064 34152 30116
rect 34204 30104 34210 30116
rect 34532 30104 34560 30212
rect 36262 30200 36268 30252
rect 36320 30200 36326 30252
rect 36814 30200 36820 30252
rect 36872 30240 36878 30252
rect 37277 30243 37335 30249
rect 37277 30240 37289 30243
rect 36872 30212 37289 30240
rect 36872 30200 36878 30212
rect 37277 30209 37289 30212
rect 37323 30240 37335 30243
rect 37366 30240 37372 30252
rect 37323 30212 37372 30240
rect 37323 30209 37335 30212
rect 37277 30203 37335 30209
rect 37366 30200 37372 30212
rect 37424 30200 37430 30252
rect 37550 30200 37556 30252
rect 37608 30200 37614 30252
rect 38120 30249 38148 30280
rect 39482 30268 39488 30320
rect 39540 30268 39546 30320
rect 39776 30308 39804 30348
rect 40034 30308 40040 30320
rect 39776 30280 40040 30308
rect 40034 30268 40040 30280
rect 40092 30268 40098 30320
rect 37921 30243 37979 30249
rect 37921 30209 37933 30243
rect 37967 30209 37979 30243
rect 37921 30203 37979 30209
rect 38105 30243 38163 30249
rect 38105 30209 38117 30243
rect 38151 30209 38163 30243
rect 38105 30203 38163 30209
rect 36170 30132 36176 30184
rect 36228 30172 36234 30184
rect 36357 30175 36415 30181
rect 36357 30172 36369 30175
rect 36228 30144 36369 30172
rect 36228 30132 36234 30144
rect 36357 30141 36369 30144
rect 36403 30141 36415 30175
rect 37936 30172 37964 30203
rect 36357 30135 36415 30141
rect 36464 30144 37964 30172
rect 36464 30104 36492 30144
rect 38010 30132 38016 30184
rect 38068 30172 38074 30184
rect 38120 30172 38148 30203
rect 38194 30200 38200 30252
rect 38252 30200 38258 30252
rect 38068 30144 38148 30172
rect 38068 30132 38074 30144
rect 38470 30132 38476 30184
rect 38528 30132 38534 30184
rect 40221 30175 40279 30181
rect 40221 30172 40233 30175
rect 39500 30144 40233 30172
rect 34204 30076 34494 30104
rect 34532 30076 36492 30104
rect 34204 30064 34210 30076
rect 33781 30039 33839 30045
rect 33781 30036 33793 30039
rect 33652 30008 33793 30036
rect 33652 29996 33658 30008
rect 33781 30005 33793 30008
rect 33827 30005 33839 30039
rect 33781 29999 33839 30005
rect 33965 30039 34023 30045
rect 33965 30005 33977 30039
rect 34011 30036 34023 30039
rect 34330 30036 34336 30048
rect 34011 30008 34336 30036
rect 34011 30005 34023 30008
rect 33965 29999 34023 30005
rect 34330 29996 34336 30008
rect 34388 29996 34394 30048
rect 34466 30036 34494 30076
rect 34609 30039 34667 30045
rect 34609 30036 34621 30039
rect 34466 30008 34621 30036
rect 34609 30005 34621 30008
rect 34655 30036 34667 30039
rect 35342 30036 35348 30048
rect 34655 30008 35348 30036
rect 34655 30005 34667 30008
rect 34609 29999 34667 30005
rect 35342 29996 35348 30008
rect 35400 29996 35406 30048
rect 36078 29996 36084 30048
rect 36136 30036 36142 30048
rect 36265 30039 36323 30045
rect 36265 30036 36277 30039
rect 36136 30008 36277 30036
rect 36136 29996 36142 30008
rect 36265 30005 36277 30008
rect 36311 30005 36323 30039
rect 36265 29999 36323 30005
rect 36354 29996 36360 30048
rect 36412 30036 36418 30048
rect 36633 30039 36691 30045
rect 36633 30036 36645 30039
rect 36412 30008 36645 30036
rect 36412 29996 36418 30008
rect 36633 30005 36645 30008
rect 36679 30036 36691 30039
rect 37274 30036 37280 30048
rect 36679 30008 37280 30036
rect 36679 30005 36691 30008
rect 36633 29999 36691 30005
rect 37274 29996 37280 30008
rect 37332 29996 37338 30048
rect 37366 29996 37372 30048
rect 37424 29996 37430 30048
rect 37826 29996 37832 30048
rect 37884 29996 37890 30048
rect 38286 29996 38292 30048
rect 38344 30036 38350 30048
rect 39500 30036 39528 30144
rect 40221 30141 40233 30144
rect 40267 30141 40279 30175
rect 40221 30135 40279 30141
rect 38344 30008 39528 30036
rect 38344 29996 38350 30008
rect 1104 29946 40572 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 40572 29946
rect 1104 29872 40572 29894
rect 4614 29792 4620 29844
rect 4672 29832 4678 29844
rect 5537 29835 5595 29841
rect 5537 29832 5549 29835
rect 4672 29804 5549 29832
rect 4672 29792 4678 29804
rect 5537 29801 5549 29804
rect 5583 29832 5595 29835
rect 6822 29832 6828 29844
rect 5583 29804 6828 29832
rect 5583 29801 5595 29804
rect 5537 29795 5595 29801
rect 6822 29792 6828 29804
rect 6880 29792 6886 29844
rect 10505 29835 10563 29841
rect 10505 29801 10517 29835
rect 10551 29832 10563 29835
rect 11054 29832 11060 29844
rect 10551 29804 11060 29832
rect 10551 29801 10563 29804
rect 10505 29795 10563 29801
rect 11054 29792 11060 29804
rect 11112 29832 11118 29844
rect 12250 29832 12256 29844
rect 11112 29804 12256 29832
rect 11112 29792 11118 29804
rect 12250 29792 12256 29804
rect 12308 29792 12314 29844
rect 14550 29792 14556 29844
rect 14608 29832 14614 29844
rect 16298 29832 16304 29844
rect 14608 29804 16304 29832
rect 14608 29792 14614 29804
rect 16298 29792 16304 29804
rect 16356 29792 16362 29844
rect 18322 29792 18328 29844
rect 18380 29792 18386 29844
rect 18506 29792 18512 29844
rect 18564 29832 18570 29844
rect 21450 29832 21456 29844
rect 18564 29804 21456 29832
rect 18564 29792 18570 29804
rect 21450 29792 21456 29804
rect 21508 29792 21514 29844
rect 21910 29792 21916 29844
rect 21968 29832 21974 29844
rect 21968 29804 27292 29832
rect 21968 29792 21974 29804
rect 10686 29764 10692 29776
rect 10244 29736 10692 29764
rect 4062 29656 4068 29708
rect 4120 29656 4126 29708
rect 4798 29656 4804 29708
rect 4856 29696 4862 29708
rect 6273 29699 6331 29705
rect 6273 29696 6285 29699
rect 4856 29668 6285 29696
rect 4856 29656 4862 29668
rect 6273 29665 6285 29668
rect 6319 29696 6331 29699
rect 6546 29696 6552 29708
rect 6319 29668 6552 29696
rect 6319 29665 6331 29668
rect 6273 29659 6331 29665
rect 6546 29656 6552 29668
rect 6604 29656 6610 29708
rect 9398 29656 9404 29708
rect 9456 29696 9462 29708
rect 10244 29705 10272 29736
rect 10686 29724 10692 29736
rect 10744 29724 10750 29776
rect 12529 29767 12587 29773
rect 12529 29733 12541 29767
rect 12575 29764 12587 29767
rect 13446 29764 13452 29776
rect 12575 29736 13452 29764
rect 12575 29733 12587 29736
rect 12529 29727 12587 29733
rect 13446 29724 13452 29736
rect 13504 29724 13510 29776
rect 13541 29767 13599 29773
rect 13541 29733 13553 29767
rect 13587 29764 13599 29767
rect 14369 29767 14427 29773
rect 14369 29764 14381 29767
rect 13587 29736 14381 29764
rect 13587 29733 13599 29736
rect 13541 29727 13599 29733
rect 14369 29733 14381 29736
rect 14415 29733 14427 29767
rect 14369 29727 14427 29733
rect 14734 29724 14740 29776
rect 14792 29764 14798 29776
rect 19150 29764 19156 29776
rect 14792 29736 19156 29764
rect 14792 29724 14798 29736
rect 19150 29724 19156 29736
rect 19208 29764 19214 29776
rect 19613 29767 19671 29773
rect 19613 29764 19625 29767
rect 19208 29736 19625 29764
rect 19208 29724 19214 29736
rect 19613 29733 19625 29736
rect 19659 29733 19671 29767
rect 23474 29764 23480 29776
rect 19613 29727 19671 29733
rect 23124 29736 23480 29764
rect 9861 29699 9919 29705
rect 9861 29696 9873 29699
rect 9456 29668 9873 29696
rect 9456 29656 9462 29668
rect 9861 29665 9873 29668
rect 9907 29665 9919 29699
rect 9861 29659 9919 29665
rect 10229 29699 10287 29705
rect 10229 29665 10241 29699
rect 10275 29665 10287 29699
rect 10229 29659 10287 29665
rect 10321 29699 10379 29705
rect 10321 29665 10333 29699
rect 10367 29696 10379 29699
rect 10778 29696 10784 29708
rect 10367 29668 10784 29696
rect 10367 29665 10379 29668
rect 10321 29659 10379 29665
rect 10778 29656 10784 29668
rect 10836 29656 10842 29708
rect 12161 29699 12219 29705
rect 11164 29668 11928 29696
rect 3786 29588 3792 29640
rect 3844 29588 3850 29640
rect 5994 29588 6000 29640
rect 6052 29628 6058 29640
rect 6089 29631 6147 29637
rect 6089 29628 6101 29631
rect 6052 29600 6101 29628
rect 6052 29588 6058 29600
rect 6089 29597 6101 29600
rect 6135 29597 6147 29631
rect 6089 29591 6147 29597
rect 9950 29588 9956 29640
rect 10008 29628 10014 29640
rect 10597 29631 10655 29637
rect 10597 29628 10609 29631
rect 10008 29600 10609 29628
rect 10008 29588 10014 29600
rect 10597 29597 10609 29600
rect 10643 29597 10655 29631
rect 10597 29591 10655 29597
rect 10686 29588 10692 29640
rect 10744 29628 10750 29640
rect 11164 29637 11192 29668
rect 11149 29631 11207 29637
rect 11149 29628 11161 29631
rect 10744 29600 11161 29628
rect 10744 29588 10750 29600
rect 11149 29597 11161 29600
rect 11195 29597 11207 29631
rect 11149 29591 11207 29597
rect 11330 29588 11336 29640
rect 11388 29628 11394 29640
rect 11425 29631 11483 29637
rect 11425 29628 11437 29631
rect 11388 29600 11437 29628
rect 11388 29588 11394 29600
rect 11425 29597 11437 29600
rect 11471 29597 11483 29631
rect 11425 29591 11483 29597
rect 11790 29588 11796 29640
rect 11848 29588 11854 29640
rect 11900 29628 11928 29668
rect 12161 29665 12173 29699
rect 12207 29696 12219 29699
rect 13078 29696 13084 29708
rect 12207 29668 13084 29696
rect 12207 29665 12219 29668
rect 12161 29659 12219 29665
rect 11958 29631 12016 29637
rect 11958 29628 11970 29631
rect 11900 29600 11970 29628
rect 11958 29597 11970 29600
rect 12004 29597 12016 29631
rect 11958 29591 12016 29597
rect 12069 29631 12127 29637
rect 12069 29597 12081 29631
rect 12115 29597 12127 29631
rect 12069 29591 12127 29597
rect 7190 29560 7196 29572
rect 5290 29532 7196 29560
rect 7190 29520 7196 29532
rect 7248 29520 7254 29572
rect 9674 29560 9680 29572
rect 7300 29532 9680 29560
rect 5629 29495 5687 29501
rect 5629 29461 5641 29495
rect 5675 29492 5687 29495
rect 5718 29492 5724 29504
rect 5675 29464 5724 29492
rect 5675 29461 5687 29464
rect 5629 29455 5687 29461
rect 5718 29452 5724 29464
rect 5776 29452 5782 29504
rect 5997 29495 6055 29501
rect 5997 29461 6009 29495
rect 6043 29492 6055 29495
rect 6178 29492 6184 29504
rect 6043 29464 6184 29492
rect 6043 29461 6055 29464
rect 5997 29455 6055 29461
rect 6178 29452 6184 29464
rect 6236 29492 6242 29504
rect 7300 29492 7328 29532
rect 9674 29520 9680 29532
rect 9732 29520 9738 29572
rect 11514 29520 11520 29572
rect 11572 29560 11578 29572
rect 11701 29563 11759 29569
rect 11701 29560 11713 29563
rect 11572 29532 11713 29560
rect 11572 29520 11578 29532
rect 11701 29529 11713 29532
rect 11747 29529 11759 29563
rect 11701 29523 11759 29529
rect 6236 29464 7328 29492
rect 6236 29452 6242 29464
rect 9490 29452 9496 29504
rect 9548 29492 9554 29504
rect 12084 29492 12112 29591
rect 12176 29504 12204 29659
rect 12544 29640 12572 29668
rect 13078 29656 13084 29668
rect 13136 29656 13142 29708
rect 14185 29699 14243 29705
rect 14185 29696 14197 29699
rect 13372 29668 13584 29696
rect 12342 29588 12348 29640
rect 12400 29588 12406 29640
rect 12526 29588 12532 29640
rect 12584 29588 12590 29640
rect 12713 29631 12771 29637
rect 12713 29597 12725 29631
rect 12759 29597 12771 29631
rect 12713 29591 12771 29597
rect 9548 29464 12112 29492
rect 9548 29452 9554 29464
rect 12158 29452 12164 29504
rect 12216 29452 12222 29504
rect 12342 29452 12348 29504
rect 12400 29492 12406 29504
rect 12728 29492 12756 29591
rect 12894 29588 12900 29640
rect 12952 29588 12958 29640
rect 13372 29637 13400 29668
rect 13357 29631 13415 29637
rect 13357 29597 13369 29631
rect 13403 29597 13415 29631
rect 13357 29591 13415 29597
rect 13449 29631 13507 29637
rect 13449 29597 13461 29631
rect 13495 29597 13507 29631
rect 13449 29591 13507 29597
rect 12805 29563 12863 29569
rect 12805 29529 12817 29563
rect 12851 29560 12863 29563
rect 13464 29560 13492 29591
rect 12851 29532 13492 29560
rect 13556 29560 13584 29668
rect 13648 29668 14197 29696
rect 13648 29637 13676 29668
rect 14185 29665 14197 29668
rect 14231 29665 14243 29699
rect 14185 29659 14243 29665
rect 15470 29656 15476 29708
rect 15528 29656 15534 29708
rect 19978 29696 19984 29708
rect 15580 29668 16896 29696
rect 13633 29631 13691 29637
rect 13633 29597 13645 29631
rect 13679 29597 13691 29631
rect 13633 29591 13691 29597
rect 14090 29588 14096 29640
rect 14148 29588 14154 29640
rect 14277 29631 14335 29637
rect 14277 29628 14289 29631
rect 14200 29600 14289 29628
rect 14108 29560 14136 29588
rect 14200 29572 14228 29600
rect 14277 29597 14289 29600
rect 14323 29597 14335 29631
rect 14277 29591 14335 29597
rect 14366 29588 14372 29640
rect 14424 29588 14430 29640
rect 14553 29631 14611 29637
rect 14553 29597 14565 29631
rect 14599 29628 14611 29631
rect 14642 29628 14648 29640
rect 14599 29600 14648 29628
rect 14599 29597 14611 29600
rect 14553 29591 14611 29597
rect 14642 29588 14648 29600
rect 14700 29628 14706 29640
rect 14918 29628 14924 29640
rect 14700 29600 14924 29628
rect 14700 29588 14706 29600
rect 14918 29588 14924 29600
rect 14976 29588 14982 29640
rect 15010 29588 15016 29640
rect 15068 29628 15074 29640
rect 15580 29637 15608 29668
rect 15105 29631 15163 29637
rect 15105 29628 15117 29631
rect 15068 29600 15117 29628
rect 15068 29588 15074 29600
rect 15105 29597 15117 29600
rect 15151 29628 15163 29631
rect 15565 29631 15623 29637
rect 15151 29600 15424 29628
rect 15151 29597 15163 29600
rect 15105 29591 15163 29597
rect 13556 29532 14136 29560
rect 12851 29529 12863 29532
rect 12805 29523 12863 29529
rect 14182 29520 14188 29572
rect 14240 29520 14246 29572
rect 15396 29560 15424 29600
rect 15565 29597 15577 29631
rect 15611 29597 15623 29631
rect 15565 29591 15623 29597
rect 15746 29588 15752 29640
rect 15804 29628 15810 29640
rect 15933 29631 15991 29637
rect 15933 29628 15945 29631
rect 15804 29600 15945 29628
rect 15804 29588 15810 29600
rect 15933 29597 15945 29600
rect 15979 29597 15991 29631
rect 15933 29591 15991 29597
rect 16117 29631 16175 29637
rect 16117 29597 16129 29631
rect 16163 29628 16175 29631
rect 16482 29628 16488 29640
rect 16163 29600 16488 29628
rect 16163 29597 16175 29600
rect 16117 29591 16175 29597
rect 16482 29588 16488 29600
rect 16540 29588 16546 29640
rect 16868 29637 16896 29668
rect 17880 29668 19984 29696
rect 16853 29631 16911 29637
rect 16853 29597 16865 29631
rect 16899 29628 16911 29631
rect 16942 29628 16948 29640
rect 16899 29600 16948 29628
rect 16899 29597 16911 29600
rect 16853 29591 16911 29597
rect 16942 29588 16948 29600
rect 17000 29588 17006 29640
rect 17126 29588 17132 29640
rect 17184 29588 17190 29640
rect 17880 29637 17908 29668
rect 19978 29656 19984 29668
rect 20036 29656 20042 29708
rect 23014 29696 23020 29708
rect 22066 29668 23020 29696
rect 17865 29631 17923 29637
rect 17865 29597 17877 29631
rect 17911 29597 17923 29631
rect 17865 29591 17923 29597
rect 15396 29532 16160 29560
rect 12400 29464 12756 29492
rect 12400 29452 12406 29464
rect 13170 29452 13176 29504
rect 13228 29452 13234 29504
rect 13814 29452 13820 29504
rect 13872 29492 13878 29504
rect 15197 29495 15255 29501
rect 15197 29492 15209 29495
rect 13872 29464 15209 29492
rect 13872 29452 13878 29464
rect 15197 29461 15209 29464
rect 15243 29461 15255 29495
rect 16132 29492 16160 29532
rect 16758 29520 16764 29572
rect 16816 29560 16822 29572
rect 17880 29560 17908 29591
rect 18506 29588 18512 29640
rect 18564 29588 18570 29640
rect 18782 29588 18788 29640
rect 18840 29588 18846 29640
rect 18874 29588 18880 29640
rect 18932 29588 18938 29640
rect 18966 29588 18972 29640
rect 19024 29628 19030 29640
rect 19061 29631 19119 29637
rect 19061 29628 19073 29631
rect 19024 29600 19073 29628
rect 19024 29588 19030 29600
rect 19061 29597 19073 29600
rect 19107 29597 19119 29631
rect 19061 29591 19119 29597
rect 16816 29532 17908 29560
rect 18892 29560 18920 29588
rect 19245 29563 19303 29569
rect 19245 29560 19257 29563
rect 18892 29532 19257 29560
rect 16816 29520 16822 29532
rect 19245 29529 19257 29532
rect 19291 29529 19303 29563
rect 19245 29523 19303 29529
rect 19426 29520 19432 29572
rect 19484 29560 19490 29572
rect 22066 29560 22094 29668
rect 23014 29656 23020 29668
rect 23072 29656 23078 29708
rect 22278 29588 22284 29640
rect 22336 29588 22342 29640
rect 22646 29588 22652 29640
rect 22704 29588 22710 29640
rect 22738 29588 22744 29640
rect 22796 29628 22802 29640
rect 23124 29637 23152 29736
rect 23474 29724 23480 29736
rect 23532 29724 23538 29776
rect 23842 29764 23848 29776
rect 23584 29736 23848 29764
rect 23584 29696 23612 29736
rect 23842 29724 23848 29736
rect 23900 29724 23906 29776
rect 24118 29724 24124 29776
rect 24176 29764 24182 29776
rect 24176 29736 24808 29764
rect 24176 29724 24182 29736
rect 24210 29696 24216 29708
rect 23216 29668 23612 29696
rect 23768 29668 24216 29696
rect 23216 29637 23244 29668
rect 22833 29631 22891 29637
rect 22833 29628 22845 29631
rect 22796 29600 22845 29628
rect 22796 29588 22802 29600
rect 22833 29597 22845 29600
rect 22879 29597 22891 29631
rect 22833 29591 22891 29597
rect 23109 29631 23167 29637
rect 23109 29597 23121 29631
rect 23155 29597 23167 29631
rect 23109 29591 23167 29597
rect 23201 29631 23259 29637
rect 23201 29597 23213 29631
rect 23247 29597 23259 29631
rect 23201 29591 23259 29597
rect 23382 29588 23388 29640
rect 23440 29588 23446 29640
rect 23477 29631 23535 29637
rect 23477 29597 23489 29631
rect 23523 29628 23535 29631
rect 23566 29628 23572 29640
rect 23523 29600 23572 29628
rect 23523 29597 23535 29600
rect 23477 29591 23535 29597
rect 23566 29588 23572 29600
rect 23624 29588 23630 29640
rect 23768 29637 23796 29668
rect 24210 29656 24216 29668
rect 24268 29656 24274 29708
rect 23753 29631 23811 29637
rect 23753 29597 23765 29631
rect 23799 29628 23811 29631
rect 23842 29628 23848 29640
rect 23799 29600 23848 29628
rect 23799 29597 23811 29600
rect 23753 29591 23811 29597
rect 23842 29588 23848 29600
rect 23900 29588 23906 29640
rect 23937 29631 23995 29637
rect 23937 29597 23949 29631
rect 23983 29628 23995 29631
rect 24026 29628 24032 29640
rect 23983 29600 24032 29628
rect 23983 29597 23995 29600
rect 23937 29591 23995 29597
rect 24026 29588 24032 29600
rect 24084 29628 24090 29640
rect 24780 29637 24808 29736
rect 26418 29724 26424 29776
rect 26476 29764 26482 29776
rect 27264 29773 27292 29804
rect 27430 29792 27436 29844
rect 27488 29832 27494 29844
rect 33870 29832 33876 29844
rect 27488 29804 33876 29832
rect 27488 29792 27494 29804
rect 33870 29792 33876 29804
rect 33928 29792 33934 29844
rect 35250 29792 35256 29844
rect 35308 29832 35314 29844
rect 35805 29835 35863 29841
rect 35805 29832 35817 29835
rect 35308 29804 35817 29832
rect 35308 29792 35314 29804
rect 35805 29801 35817 29804
rect 35851 29801 35863 29835
rect 35805 29795 35863 29801
rect 35989 29835 36047 29841
rect 35989 29801 36001 29835
rect 36035 29832 36047 29835
rect 36446 29832 36452 29844
rect 36035 29804 36452 29832
rect 36035 29801 36047 29804
rect 35989 29795 36047 29801
rect 36446 29792 36452 29804
rect 36504 29792 36510 29844
rect 38378 29792 38384 29844
rect 38436 29792 38442 29844
rect 27157 29767 27215 29773
rect 27157 29764 27169 29767
rect 26476 29736 27169 29764
rect 26476 29724 26482 29736
rect 27157 29733 27169 29736
rect 27203 29733 27215 29767
rect 27157 29727 27215 29733
rect 27249 29767 27307 29773
rect 27249 29733 27261 29767
rect 27295 29733 27307 29767
rect 27249 29727 27307 29733
rect 27798 29724 27804 29776
rect 27856 29724 27862 29776
rect 27890 29724 27896 29776
rect 27948 29764 27954 29776
rect 31018 29764 31024 29776
rect 27948 29736 31024 29764
rect 27948 29724 27954 29736
rect 31018 29724 31024 29736
rect 31076 29724 31082 29776
rect 33594 29764 33600 29776
rect 32411 29736 33600 29764
rect 25038 29656 25044 29708
rect 25096 29696 25102 29708
rect 25225 29699 25283 29705
rect 25225 29696 25237 29699
rect 25096 29668 25237 29696
rect 25096 29656 25102 29668
rect 25225 29665 25237 29668
rect 25271 29665 25283 29699
rect 27816 29696 27844 29724
rect 25225 29659 25283 29665
rect 25332 29668 26004 29696
rect 27816 29668 28396 29696
rect 25332 29640 25360 29668
rect 24765 29631 24823 29637
rect 24084 29600 24716 29628
rect 24084 29588 24090 29600
rect 19484 29532 22094 29560
rect 22373 29563 22431 29569
rect 19484 29520 19490 29532
rect 22373 29529 22385 29563
rect 22419 29560 22431 29563
rect 22554 29560 22560 29572
rect 22419 29532 22560 29560
rect 22419 29529 22431 29532
rect 22373 29523 22431 29529
rect 22554 29520 22560 29532
rect 22612 29520 22618 29572
rect 24581 29563 24639 29569
rect 24581 29529 24593 29563
rect 24627 29529 24639 29563
rect 24688 29560 24716 29600
rect 24765 29597 24777 29631
rect 24811 29597 24823 29631
rect 24765 29591 24823 29597
rect 25130 29588 25136 29640
rect 25188 29588 25194 29640
rect 25314 29588 25320 29640
rect 25372 29588 25378 29640
rect 25976 29637 26004 29668
rect 28368 29640 28396 29668
rect 28534 29656 28540 29708
rect 28592 29696 28598 29708
rect 30561 29699 30619 29705
rect 28592 29668 28856 29696
rect 28592 29656 28598 29668
rect 25777 29631 25835 29637
rect 25777 29597 25789 29631
rect 25823 29597 25835 29631
rect 25777 29591 25835 29597
rect 25961 29631 26019 29637
rect 25961 29597 25973 29631
rect 26007 29597 26019 29631
rect 25961 29591 26019 29597
rect 24854 29560 24860 29572
rect 24688 29532 24860 29560
rect 24581 29523 24639 29529
rect 16301 29495 16359 29501
rect 16301 29492 16313 29495
rect 16132 29464 16313 29492
rect 15197 29455 15255 29461
rect 16301 29461 16313 29464
rect 16347 29461 16359 29495
rect 16301 29455 16359 29461
rect 18601 29495 18659 29501
rect 18601 29461 18613 29495
rect 18647 29492 18659 29495
rect 19518 29492 19524 29504
rect 18647 29464 19524 29492
rect 18647 29461 18659 29464
rect 18601 29455 18659 29461
rect 19518 29452 19524 29464
rect 19576 29452 19582 29504
rect 20714 29452 20720 29504
rect 20772 29492 20778 29504
rect 21910 29492 21916 29504
rect 20772 29464 21916 29492
rect 20772 29452 20778 29464
rect 21910 29452 21916 29464
rect 21968 29452 21974 29504
rect 22462 29452 22468 29504
rect 22520 29492 22526 29504
rect 22925 29495 22983 29501
rect 22925 29492 22937 29495
rect 22520 29464 22937 29492
rect 22520 29452 22526 29464
rect 22925 29461 22937 29464
rect 22971 29461 22983 29495
rect 22925 29455 22983 29461
rect 23566 29452 23572 29504
rect 23624 29452 23630 29504
rect 24210 29452 24216 29504
rect 24268 29492 24274 29504
rect 24489 29495 24547 29501
rect 24489 29492 24501 29495
rect 24268 29464 24501 29492
rect 24268 29452 24274 29464
rect 24489 29461 24501 29464
rect 24535 29461 24547 29495
rect 24596 29492 24624 29523
rect 24854 29520 24860 29532
rect 24912 29560 24918 29572
rect 25682 29560 25688 29572
rect 24912 29532 25688 29560
rect 24912 29520 24918 29532
rect 25682 29520 25688 29532
rect 25740 29520 25746 29572
rect 25792 29560 25820 29591
rect 26234 29588 26240 29640
rect 26292 29588 26298 29640
rect 26510 29588 26516 29640
rect 26568 29588 26574 29640
rect 26605 29631 26663 29637
rect 26605 29597 26617 29631
rect 26651 29628 26663 29631
rect 26878 29628 26884 29640
rect 26651 29600 26884 29628
rect 26651 29597 26663 29600
rect 26605 29591 26663 29597
rect 26878 29588 26884 29600
rect 26936 29588 26942 29640
rect 27801 29631 27859 29637
rect 27801 29597 27813 29631
rect 27847 29597 27859 29631
rect 27801 29591 27859 29597
rect 28169 29631 28227 29637
rect 28169 29597 28181 29631
rect 28215 29628 28227 29631
rect 28258 29628 28264 29640
rect 28215 29600 28264 29628
rect 28215 29597 28227 29600
rect 28169 29591 28227 29597
rect 26142 29560 26148 29572
rect 25792 29532 26148 29560
rect 26142 29520 26148 29532
rect 26200 29520 26206 29572
rect 27065 29563 27123 29569
rect 27065 29529 27077 29563
rect 27111 29560 27123 29563
rect 27522 29560 27528 29572
rect 27111 29532 27528 29560
rect 27111 29529 27123 29532
rect 27065 29523 27123 29529
rect 27522 29520 27528 29532
rect 27580 29520 27586 29572
rect 27816 29560 27844 29591
rect 28258 29588 28264 29600
rect 28316 29588 28322 29640
rect 28350 29588 28356 29640
rect 28408 29588 28414 29640
rect 28828 29637 28856 29668
rect 30561 29665 30573 29699
rect 30607 29696 30619 29699
rect 31754 29696 31760 29708
rect 30607 29668 31760 29696
rect 30607 29665 30619 29668
rect 30561 29659 30619 29665
rect 31754 29656 31760 29668
rect 31812 29656 31818 29708
rect 31846 29656 31852 29708
rect 31904 29696 31910 29708
rect 32411 29696 32439 29736
rect 31904 29668 32439 29696
rect 32493 29699 32551 29705
rect 31904 29656 31910 29668
rect 32493 29665 32505 29699
rect 32539 29696 32551 29699
rect 33042 29696 33048 29708
rect 32539 29668 33048 29696
rect 32539 29665 32551 29668
rect 32493 29659 32551 29665
rect 33042 29656 33048 29668
rect 33100 29656 33106 29708
rect 33152 29705 33180 29736
rect 33594 29724 33600 29736
rect 33652 29724 33658 29776
rect 34238 29724 34244 29776
rect 34296 29764 34302 29776
rect 34882 29764 34888 29776
rect 34296 29736 34888 29764
rect 34296 29724 34302 29736
rect 34882 29724 34888 29736
rect 34940 29724 34946 29776
rect 35158 29724 35164 29776
rect 35216 29724 35222 29776
rect 36078 29724 36084 29776
rect 36136 29764 36142 29776
rect 36357 29767 36415 29773
rect 36357 29764 36369 29767
rect 36136 29736 36369 29764
rect 36136 29724 36142 29736
rect 36357 29733 36369 29736
rect 36403 29733 36415 29767
rect 36538 29764 36544 29776
rect 36357 29727 36415 29733
rect 36464 29736 36544 29764
rect 33137 29699 33195 29705
rect 33137 29665 33149 29699
rect 33183 29665 33195 29699
rect 33137 29659 33195 29665
rect 33229 29699 33287 29705
rect 33229 29665 33241 29699
rect 33275 29696 33287 29699
rect 33502 29696 33508 29708
rect 33275 29668 33508 29696
rect 33275 29665 33287 29668
rect 33229 29659 33287 29665
rect 33502 29656 33508 29668
rect 33560 29656 33566 29708
rect 35069 29699 35127 29705
rect 35069 29696 35081 29699
rect 34072 29668 35081 29696
rect 28813 29631 28871 29637
rect 28813 29597 28825 29631
rect 28859 29597 28871 29631
rect 28813 29591 28871 29597
rect 28534 29560 28540 29572
rect 27816 29532 28540 29560
rect 28534 29520 28540 29532
rect 28592 29520 28598 29572
rect 24670 29492 24676 29504
rect 24596 29464 24676 29492
rect 24489 29455 24547 29461
rect 24670 29452 24676 29464
rect 24728 29492 24734 29504
rect 24949 29495 25007 29501
rect 24949 29492 24961 29495
rect 24728 29464 24961 29492
rect 24728 29452 24734 29464
rect 24949 29461 24961 29464
rect 24995 29461 25007 29495
rect 24949 29455 25007 29461
rect 28258 29452 28264 29504
rect 28316 29492 28322 29504
rect 28828 29492 28856 29591
rect 30466 29588 30472 29640
rect 30524 29588 30530 29640
rect 30653 29631 30711 29637
rect 30653 29597 30665 29631
rect 30699 29628 30711 29631
rect 30699 29600 30880 29628
rect 30699 29597 30711 29600
rect 30653 29591 30711 29597
rect 28316 29464 28856 29492
rect 28316 29452 28322 29464
rect 30742 29452 30748 29504
rect 30800 29452 30806 29504
rect 30852 29492 30880 29600
rect 32766 29588 32772 29640
rect 32824 29588 32830 29640
rect 32858 29588 32864 29640
rect 32916 29628 32922 29640
rect 33318 29628 33324 29640
rect 32916 29600 33324 29628
rect 32916 29588 32922 29600
rect 33318 29588 33324 29600
rect 33376 29588 33382 29640
rect 33962 29588 33968 29640
rect 34020 29628 34026 29640
rect 34072 29637 34100 29668
rect 35069 29665 35081 29668
rect 35115 29665 35127 29699
rect 35176 29696 35204 29724
rect 36170 29696 36176 29708
rect 35176 29668 36176 29696
rect 35069 29659 35127 29665
rect 36170 29656 36176 29668
rect 36228 29696 36234 29708
rect 36228 29668 36308 29696
rect 36228 29656 36234 29668
rect 34057 29631 34115 29637
rect 34057 29628 34069 29631
rect 34020 29600 34069 29628
rect 34020 29588 34026 29600
rect 34057 29597 34069 29600
rect 34103 29597 34115 29631
rect 34057 29591 34115 29597
rect 34146 29588 34152 29640
rect 34204 29588 34210 29640
rect 34238 29588 34244 29640
rect 34296 29628 34302 29640
rect 34296 29600 34652 29628
rect 34296 29588 34302 29600
rect 30926 29520 30932 29572
rect 30984 29560 30990 29572
rect 32217 29563 32275 29569
rect 30984 29532 31050 29560
rect 30984 29520 30990 29532
rect 32217 29529 32229 29563
rect 32263 29560 32275 29563
rect 32585 29563 32643 29569
rect 32585 29560 32597 29563
rect 32263 29532 32597 29560
rect 32263 29529 32275 29532
rect 32217 29523 32275 29529
rect 32585 29529 32597 29532
rect 32631 29529 32643 29563
rect 32585 29523 32643 29529
rect 33042 29520 33048 29572
rect 33100 29560 33106 29572
rect 33873 29563 33931 29569
rect 33873 29560 33885 29563
rect 33100 29532 33885 29560
rect 33100 29520 33106 29532
rect 33873 29529 33885 29532
rect 33919 29529 33931 29563
rect 34425 29563 34483 29569
rect 34425 29560 34437 29563
rect 33873 29523 33931 29529
rect 34072 29532 34437 29560
rect 31846 29492 31852 29504
rect 30852 29464 31852 29492
rect 31846 29452 31852 29464
rect 31904 29452 31910 29504
rect 31938 29452 31944 29504
rect 31996 29492 32002 29504
rect 32953 29495 33011 29501
rect 32953 29492 32965 29495
rect 31996 29464 32965 29492
rect 31996 29452 32002 29464
rect 32953 29461 32965 29464
rect 32999 29461 33011 29495
rect 32953 29455 33011 29461
rect 33226 29452 33232 29504
rect 33284 29492 33290 29504
rect 33778 29492 33784 29504
rect 33284 29464 33784 29492
rect 33284 29452 33290 29464
rect 33778 29452 33784 29464
rect 33836 29492 33842 29504
rect 34072 29492 34100 29532
rect 34425 29529 34437 29532
rect 34471 29529 34483 29563
rect 34624 29560 34652 29600
rect 34698 29588 34704 29640
rect 34756 29588 34762 29640
rect 34885 29631 34943 29637
rect 34885 29597 34897 29631
rect 34931 29597 34943 29631
rect 34885 29591 34943 29597
rect 35161 29631 35219 29637
rect 35161 29597 35173 29631
rect 35207 29628 35219 29631
rect 35434 29628 35440 29640
rect 35207 29600 35440 29628
rect 35207 29597 35219 29600
rect 35161 29591 35219 29597
rect 34900 29560 34928 29591
rect 35434 29588 35440 29600
rect 35492 29628 35498 29640
rect 36280 29637 36308 29668
rect 36464 29637 36492 29736
rect 36538 29724 36544 29736
rect 36596 29764 36602 29776
rect 38010 29764 38016 29776
rect 36596 29736 38016 29764
rect 36596 29724 36602 29736
rect 38010 29724 38016 29736
rect 38068 29724 38074 29776
rect 38473 29767 38531 29773
rect 38473 29733 38485 29767
rect 38519 29733 38531 29767
rect 38473 29727 38531 29733
rect 36630 29656 36636 29708
rect 36688 29696 36694 29708
rect 36688 29668 38240 29696
rect 36688 29656 36694 29668
rect 36265 29631 36323 29637
rect 35492 29600 35880 29628
rect 35492 29588 35498 29600
rect 34624 29532 34928 29560
rect 34425 29523 34483 29529
rect 33836 29464 34100 29492
rect 33836 29452 33842 29464
rect 34146 29452 34152 29504
rect 34204 29492 34210 29504
rect 34241 29495 34299 29501
rect 34241 29492 34253 29495
rect 34204 29464 34253 29492
rect 34204 29452 34210 29464
rect 34241 29461 34253 29464
rect 34287 29461 34299 29495
rect 34900 29492 34928 29532
rect 35066 29520 35072 29572
rect 35124 29560 35130 29572
rect 35618 29560 35624 29572
rect 35124 29532 35624 29560
rect 35124 29520 35130 29532
rect 35618 29520 35624 29532
rect 35676 29520 35682 29572
rect 35852 29569 35880 29600
rect 36265 29597 36277 29631
rect 36311 29597 36323 29631
rect 36265 29591 36323 29597
rect 36449 29631 36507 29637
rect 36449 29597 36461 29631
rect 36495 29597 36507 29631
rect 36449 29591 36507 29597
rect 36541 29631 36599 29637
rect 36541 29597 36553 29631
rect 36587 29628 36599 29631
rect 36814 29628 36820 29640
rect 36587 29600 36820 29628
rect 36587 29597 36599 29600
rect 36541 29591 36599 29597
rect 35837 29563 35895 29569
rect 35837 29529 35849 29563
rect 35883 29560 35895 29563
rect 36081 29563 36139 29569
rect 36081 29560 36093 29563
rect 35883 29532 36093 29560
rect 35883 29529 35895 29532
rect 35837 29523 35895 29529
rect 36081 29529 36093 29532
rect 36127 29529 36139 29563
rect 36280 29560 36308 29591
rect 36814 29588 36820 29600
rect 36872 29628 36878 29640
rect 37458 29628 37464 29640
rect 36872 29600 37464 29628
rect 36872 29588 36878 29600
rect 37458 29588 37464 29600
rect 37516 29628 37522 29640
rect 37642 29628 37648 29640
rect 37516 29600 37648 29628
rect 37516 29588 37522 29600
rect 37642 29588 37648 29600
rect 37700 29588 37706 29640
rect 37826 29588 37832 29640
rect 37884 29628 37890 29640
rect 38105 29631 38163 29637
rect 38105 29628 38117 29631
rect 37884 29600 38117 29628
rect 37884 29588 37890 29600
rect 38105 29597 38117 29600
rect 38151 29597 38163 29631
rect 38212 29628 38240 29668
rect 38378 29656 38384 29708
rect 38436 29696 38442 29708
rect 38488 29696 38516 29727
rect 38436 29668 38516 29696
rect 38672 29668 39528 29696
rect 38436 29656 38442 29668
rect 38672 29640 38700 29668
rect 38212 29600 38516 29628
rect 38105 29591 38163 29597
rect 37366 29560 37372 29572
rect 36280 29532 37372 29560
rect 36081 29523 36139 29529
rect 37366 29520 37372 29532
rect 37424 29560 37430 29572
rect 37553 29563 37611 29569
rect 37553 29560 37565 29563
rect 37424 29532 37565 29560
rect 37424 29520 37430 29532
rect 37553 29529 37565 29532
rect 37599 29529 37611 29563
rect 37553 29523 37611 29529
rect 37921 29563 37979 29569
rect 37921 29529 37933 29563
rect 37967 29560 37979 29563
rect 37967 29532 38332 29560
rect 37967 29529 37979 29532
rect 37921 29523 37979 29529
rect 35986 29492 35992 29504
rect 34900 29464 35992 29492
rect 34241 29455 34299 29461
rect 35986 29452 35992 29464
rect 36044 29452 36050 29504
rect 36170 29452 36176 29504
rect 36228 29492 36234 29504
rect 37936 29492 37964 29523
rect 36228 29464 37964 29492
rect 36228 29452 36234 29464
rect 38010 29452 38016 29504
rect 38068 29492 38074 29504
rect 38197 29495 38255 29501
rect 38197 29492 38209 29495
rect 38068 29464 38209 29492
rect 38068 29452 38074 29464
rect 38197 29461 38209 29464
rect 38243 29461 38255 29495
rect 38304 29492 38332 29532
rect 38378 29520 38384 29572
rect 38436 29520 38442 29572
rect 38488 29560 38516 29600
rect 38654 29588 38660 29640
rect 38712 29588 38718 29640
rect 38930 29588 38936 29640
rect 38988 29628 38994 29640
rect 39025 29631 39083 29637
rect 39025 29628 39037 29631
rect 38988 29600 39037 29628
rect 38988 29588 38994 29600
rect 39025 29597 39037 29600
rect 39071 29597 39083 29631
rect 39025 29591 39083 29597
rect 39114 29588 39120 29640
rect 39172 29588 39178 29640
rect 39500 29637 39528 29668
rect 39485 29631 39543 29637
rect 39485 29597 39497 29631
rect 39531 29597 39543 29631
rect 39485 29591 39543 29597
rect 38749 29563 38807 29569
rect 38749 29560 38761 29563
rect 38488 29532 38761 29560
rect 38749 29529 38761 29532
rect 38795 29529 38807 29563
rect 38749 29523 38807 29529
rect 38654 29492 38660 29504
rect 38304 29464 38660 29492
rect 38197 29455 38255 29461
rect 38654 29452 38660 29464
rect 38712 29452 38718 29504
rect 38764 29492 38792 29523
rect 38838 29520 38844 29572
rect 38896 29520 38902 29572
rect 39132 29560 39160 29588
rect 39577 29563 39635 29569
rect 39577 29560 39589 29563
rect 39132 29532 39589 29560
rect 39577 29529 39589 29532
rect 39623 29529 39635 29563
rect 39577 29523 39635 29529
rect 39206 29492 39212 29504
rect 38764 29464 39212 29492
rect 39206 29452 39212 29464
rect 39264 29452 39270 29504
rect 39298 29452 39304 29504
rect 39356 29452 39362 29504
rect 1104 29402 40572 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 40572 29402
rect 1104 29328 40572 29350
rect 3786 29248 3792 29300
rect 3844 29288 3850 29300
rect 5534 29288 5540 29300
rect 3844 29260 5540 29288
rect 3844 29248 3850 29260
rect 4448 29161 4476 29260
rect 5534 29248 5540 29260
rect 5592 29248 5598 29300
rect 6822 29248 6828 29300
rect 6880 29288 6886 29300
rect 6880 29260 11284 29288
rect 6880 29248 6886 29260
rect 7190 29220 7196 29232
rect 5934 29192 7196 29220
rect 7190 29180 7196 29192
rect 7248 29180 7254 29232
rect 7742 29180 7748 29232
rect 7800 29180 7806 29232
rect 9490 29220 9496 29232
rect 9324 29192 9496 29220
rect 4433 29155 4491 29161
rect 4433 29121 4445 29155
rect 4479 29121 4491 29155
rect 4433 29115 4491 29121
rect 6178 29112 6184 29164
rect 6236 29112 6242 29164
rect 4798 29044 4804 29096
rect 4856 29084 4862 29096
rect 6196 29084 6224 29112
rect 4856 29056 6224 29084
rect 4856 29044 4862 29056
rect 6822 29044 6828 29096
rect 6880 29044 6886 29096
rect 7098 29044 7104 29096
rect 7156 29044 7162 29096
rect 7190 29044 7196 29096
rect 7248 29084 7254 29096
rect 7742 29084 7748 29096
rect 7248 29056 7748 29084
rect 7248 29044 7254 29056
rect 7742 29044 7748 29056
rect 7800 29044 7806 29096
rect 9217 29087 9275 29093
rect 9217 29053 9229 29087
rect 9263 29053 9275 29087
rect 9217 29047 9275 29053
rect 5994 28976 6000 29028
rect 6052 29016 6058 29028
rect 6178 29016 6184 29028
rect 6052 28988 6184 29016
rect 6052 28976 6058 28988
rect 6178 28976 6184 28988
rect 6236 28976 6242 29028
rect 8573 29019 8631 29025
rect 8573 28985 8585 29019
rect 8619 29016 8631 29019
rect 8754 29016 8760 29028
rect 8619 28988 8760 29016
rect 8619 28985 8631 28988
rect 8573 28979 8631 28985
rect 8754 28976 8760 28988
rect 8812 29016 8818 29028
rect 9232 29016 9260 29047
rect 8812 28988 9260 29016
rect 9324 29016 9352 29192
rect 9490 29180 9496 29192
rect 9548 29180 9554 29232
rect 9766 29180 9772 29232
rect 9824 29180 9830 29232
rect 11054 29220 11060 29232
rect 9876 29192 11060 29220
rect 9876 29161 9904 29192
rect 11054 29180 11060 29192
rect 11112 29180 11118 29232
rect 9401 29155 9459 29161
rect 9401 29121 9413 29155
rect 9447 29152 9459 29155
rect 9861 29155 9919 29161
rect 9861 29152 9873 29155
rect 9447 29124 9873 29152
rect 9447 29121 9459 29124
rect 9401 29115 9459 29121
rect 9861 29121 9873 29124
rect 9907 29121 9919 29155
rect 9861 29115 9919 29121
rect 10137 29155 10195 29161
rect 10137 29121 10149 29155
rect 10183 29121 10195 29155
rect 10137 29115 10195 29121
rect 10229 29155 10287 29161
rect 10229 29121 10241 29155
rect 10275 29152 10287 29155
rect 10965 29155 11023 29161
rect 10965 29152 10977 29155
rect 10275 29124 10977 29152
rect 10275 29121 10287 29124
rect 10229 29115 10287 29121
rect 10965 29121 10977 29124
rect 11011 29121 11023 29155
rect 11256 29152 11284 29260
rect 11330 29248 11336 29300
rect 11388 29248 11394 29300
rect 11698 29288 11704 29300
rect 11532 29260 11704 29288
rect 11532 29229 11560 29260
rect 11698 29248 11704 29260
rect 11756 29248 11762 29300
rect 12069 29291 12127 29297
rect 12069 29257 12081 29291
rect 12115 29288 12127 29291
rect 12434 29288 12440 29300
rect 12115 29260 12440 29288
rect 12115 29257 12127 29260
rect 12069 29251 12127 29257
rect 12434 29248 12440 29260
rect 12492 29248 12498 29300
rect 14366 29248 14372 29300
rect 14424 29288 14430 29300
rect 16669 29291 16727 29297
rect 16669 29288 16681 29291
rect 14424 29260 16681 29288
rect 14424 29248 14430 29260
rect 16669 29257 16681 29260
rect 16715 29257 16727 29291
rect 16669 29251 16727 29257
rect 16758 29248 16764 29300
rect 16816 29288 16822 29300
rect 18693 29291 18751 29297
rect 18693 29288 18705 29291
rect 16816 29260 18705 29288
rect 16816 29248 16822 29260
rect 18693 29257 18705 29260
rect 18739 29257 18751 29291
rect 18693 29251 18751 29257
rect 19518 29248 19524 29300
rect 19576 29248 19582 29300
rect 26970 29288 26976 29300
rect 21928 29260 26976 29288
rect 11517 29223 11575 29229
rect 11517 29189 11529 29223
rect 11563 29189 11575 29223
rect 11974 29220 11980 29232
rect 11517 29183 11575 29189
rect 11624 29192 11980 29220
rect 11330 29152 11336 29164
rect 11256 29124 11336 29152
rect 10965 29115 11023 29121
rect 9490 29044 9496 29096
rect 9548 29084 9554 29096
rect 9585 29087 9643 29093
rect 9585 29084 9597 29087
rect 9548 29056 9597 29084
rect 9548 29044 9554 29056
rect 9585 29053 9597 29056
rect 9631 29084 9643 29087
rect 10152 29084 10180 29115
rect 9631 29056 10180 29084
rect 10689 29087 10747 29093
rect 9631 29053 9643 29056
rect 9585 29047 9643 29053
rect 10689 29053 10701 29087
rect 10735 29053 10747 29087
rect 10689 29047 10747 29053
rect 9324 28988 9536 29016
rect 8812 28976 8818 28988
rect 9508 28960 9536 28988
rect 9950 28976 9956 29028
rect 10008 28976 10014 29028
rect 10704 28960 10732 29047
rect 10778 29044 10784 29096
rect 10836 29084 10842 29096
rect 10873 29087 10931 29093
rect 10873 29084 10885 29087
rect 10836 29056 10885 29084
rect 10836 29044 10842 29056
rect 10873 29053 10885 29056
rect 10919 29053 10931 29087
rect 10980 29084 11008 29115
rect 11330 29112 11336 29124
rect 11388 29112 11394 29164
rect 11624 29161 11652 29192
rect 11974 29180 11980 29192
rect 12032 29220 12038 29232
rect 12342 29220 12348 29232
rect 12032 29192 12348 29220
rect 12032 29180 12038 29192
rect 12342 29180 12348 29192
rect 12400 29180 12406 29232
rect 12529 29223 12587 29229
rect 12529 29189 12541 29223
rect 12575 29220 12587 29223
rect 12618 29220 12624 29232
rect 12575 29192 12624 29220
rect 12575 29189 12587 29192
rect 12529 29183 12587 29189
rect 12618 29180 12624 29192
rect 12676 29180 12682 29232
rect 14642 29180 14648 29232
rect 14700 29220 14706 29232
rect 14700 29192 15608 29220
rect 14700 29180 14706 29192
rect 11609 29155 11667 29161
rect 11609 29121 11621 29155
rect 11655 29121 11667 29155
rect 11609 29115 11667 29121
rect 11698 29112 11704 29164
rect 11756 29152 11762 29164
rect 11885 29155 11943 29161
rect 11885 29152 11897 29155
rect 11756 29124 11897 29152
rect 11756 29112 11762 29124
rect 11885 29121 11897 29124
rect 11931 29152 11943 29155
rect 12158 29152 12164 29164
rect 11931 29124 12164 29152
rect 11931 29121 11943 29124
rect 11885 29115 11943 29121
rect 12158 29112 12164 29124
rect 12216 29112 12222 29164
rect 12434 29112 12440 29164
rect 12492 29152 12498 29164
rect 15105 29155 15163 29161
rect 15105 29152 15117 29155
rect 12492 29124 15117 29152
rect 12492 29112 12498 29124
rect 15105 29121 15117 29124
rect 15151 29121 15163 29155
rect 15105 29115 15163 29121
rect 15473 29155 15531 29161
rect 15473 29121 15485 29155
rect 15519 29121 15531 29155
rect 15473 29115 15531 29121
rect 10980 29056 12434 29084
rect 10873 29047 10931 29053
rect 11330 28976 11336 29028
rect 11388 29016 11394 29028
rect 12406 29016 12434 29056
rect 12526 29044 12532 29096
rect 12584 29084 12590 29096
rect 12621 29087 12679 29093
rect 12621 29084 12633 29087
rect 12584 29056 12633 29084
rect 12584 29044 12590 29056
rect 12621 29053 12633 29056
rect 12667 29053 12679 29087
rect 12621 29047 12679 29053
rect 15010 29044 15016 29096
rect 15068 29044 15074 29096
rect 15286 29044 15292 29096
rect 15344 29044 15350 29096
rect 13814 29016 13820 29028
rect 11388 28988 11836 29016
rect 12406 28988 13820 29016
rect 11388 28976 11394 28988
rect 4696 28951 4754 28957
rect 4696 28917 4708 28951
rect 4742 28948 4754 28951
rect 5718 28948 5724 28960
rect 4742 28920 5724 28948
rect 4742 28917 4754 28920
rect 4696 28911 4754 28917
rect 5718 28908 5724 28920
rect 5776 28908 5782 28960
rect 8662 28908 8668 28960
rect 8720 28908 8726 28960
rect 9490 28948 9496 28960
rect 9471 28920 9496 28948
rect 9490 28908 9496 28920
rect 9548 28908 9554 28960
rect 9585 28951 9643 28957
rect 9585 28917 9597 28951
rect 9631 28948 9643 28951
rect 9674 28948 9680 28960
rect 9631 28920 9680 28948
rect 9631 28917 9643 28920
rect 9585 28911 9643 28917
rect 9674 28908 9680 28920
rect 9732 28908 9738 28960
rect 10410 28908 10416 28960
rect 10468 28908 10474 28960
rect 10686 28908 10692 28960
rect 10744 28948 10750 28960
rect 11698 28948 11704 28960
rect 10744 28920 11704 28948
rect 10744 28908 10750 28920
rect 11698 28908 11704 28920
rect 11756 28908 11762 28960
rect 11808 28948 11836 28988
rect 13814 28976 13820 28988
rect 13872 28976 13878 29028
rect 15488 29016 15516 29115
rect 15580 29084 15608 29192
rect 16022 29180 16028 29232
rect 16080 29220 16086 29232
rect 16080 29192 17172 29220
rect 16080 29180 16086 29192
rect 15838 29112 15844 29164
rect 15896 29112 15902 29164
rect 15933 29155 15991 29161
rect 15933 29121 15945 29155
rect 15979 29152 15991 29155
rect 16482 29152 16488 29164
rect 15979 29124 16488 29152
rect 15979 29121 15991 29124
rect 15933 29115 15991 29121
rect 16482 29112 16488 29124
rect 16540 29152 16546 29164
rect 16853 29155 16911 29161
rect 16853 29152 16865 29155
rect 16540 29124 16865 29152
rect 16540 29112 16546 29124
rect 16853 29121 16865 29124
rect 16899 29121 16911 29155
rect 16853 29115 16911 29121
rect 16758 29084 16764 29096
rect 15580 29056 16764 29084
rect 16758 29044 16764 29056
rect 16816 29044 16822 29096
rect 16868 29084 16896 29115
rect 17034 29112 17040 29164
rect 17092 29112 17098 29164
rect 17144 29161 17172 29192
rect 18782 29180 18788 29232
rect 18840 29220 18846 29232
rect 19337 29223 19395 29229
rect 19337 29220 19349 29223
rect 18840 29192 19349 29220
rect 18840 29180 18846 29192
rect 19337 29189 19349 29192
rect 19383 29220 19395 29223
rect 19383 29192 21036 29220
rect 19383 29189 19395 29192
rect 19337 29183 19395 29189
rect 17129 29155 17187 29161
rect 17129 29121 17141 29155
rect 17175 29121 17187 29155
rect 17129 29115 17187 29121
rect 17586 29112 17592 29164
rect 17644 29112 17650 29164
rect 17862 29112 17868 29164
rect 17920 29112 17926 29164
rect 19521 29155 19579 29161
rect 19521 29152 19533 29155
rect 19306 29124 19533 29152
rect 17313 29087 17371 29093
rect 17313 29084 17325 29087
rect 16868 29056 17325 29084
rect 17313 29053 17325 29056
rect 17359 29053 17371 29087
rect 17313 29047 17371 29053
rect 18966 29044 18972 29096
rect 19024 29084 19030 29096
rect 19306 29084 19334 29124
rect 19521 29121 19533 29124
rect 19567 29121 19579 29155
rect 19521 29115 19579 29121
rect 19705 29155 19763 29161
rect 19705 29121 19717 29155
rect 19751 29152 19763 29155
rect 20714 29152 20720 29164
rect 19751 29124 20720 29152
rect 19751 29121 19763 29124
rect 19705 29115 19763 29121
rect 19024 29056 19334 29084
rect 19536 29084 19564 29115
rect 20714 29112 20720 29124
rect 20772 29112 20778 29164
rect 20898 29112 20904 29164
rect 20956 29112 20962 29164
rect 20806 29084 20812 29096
rect 19536 29056 20812 29084
rect 19024 29044 19030 29056
rect 20806 29044 20812 29056
rect 20864 29044 20870 29096
rect 16942 29016 16948 29028
rect 15488 28988 16948 29016
rect 16942 28976 16948 28988
rect 17000 28976 17006 29028
rect 18598 28976 18604 29028
rect 18656 29016 18662 29028
rect 19061 29019 19119 29025
rect 19061 29016 19073 29019
rect 18656 28988 19073 29016
rect 18656 28976 18662 28988
rect 19061 28985 19073 28988
rect 19107 28985 19119 29019
rect 19061 28979 19119 28985
rect 20714 28976 20720 29028
rect 20772 28976 20778 29028
rect 21008 29016 21036 29192
rect 21174 29180 21180 29232
rect 21232 29220 21238 29232
rect 21928 29220 21956 29260
rect 26970 29248 26976 29260
rect 27028 29248 27034 29300
rect 27249 29291 27307 29297
rect 27249 29288 27261 29291
rect 27080 29260 27261 29288
rect 21232 29192 21956 29220
rect 21232 29180 21238 29192
rect 22646 29180 22652 29232
rect 22704 29220 22710 29232
rect 23658 29220 23664 29232
rect 22704 29192 23664 29220
rect 22704 29180 22710 29192
rect 23658 29180 23664 29192
rect 23716 29220 23722 29232
rect 25130 29220 25136 29232
rect 23716 29192 24164 29220
rect 23716 29180 23722 29192
rect 21082 29112 21088 29164
rect 21140 29152 21146 29164
rect 21450 29152 21456 29164
rect 21140 29124 21456 29152
rect 21140 29112 21146 29124
rect 21450 29112 21456 29124
rect 21508 29112 21514 29164
rect 21542 29112 21548 29164
rect 21600 29112 21606 29164
rect 22097 29155 22155 29161
rect 22097 29152 22109 29155
rect 21652 29124 22109 29152
rect 21266 29044 21272 29096
rect 21324 29084 21330 29096
rect 21652 29084 21680 29124
rect 22097 29121 22109 29124
rect 22143 29121 22155 29155
rect 22097 29115 22155 29121
rect 23014 29112 23020 29164
rect 23072 29152 23078 29164
rect 23109 29155 23167 29161
rect 23109 29152 23121 29155
rect 23072 29124 23121 29152
rect 23072 29112 23078 29124
rect 23109 29121 23121 29124
rect 23155 29121 23167 29155
rect 23109 29115 23167 29121
rect 23293 29155 23351 29161
rect 23293 29121 23305 29155
rect 23339 29152 23351 29155
rect 23474 29152 23480 29164
rect 23339 29124 23480 29152
rect 23339 29121 23351 29124
rect 23293 29115 23351 29121
rect 23474 29112 23480 29124
rect 23532 29112 23538 29164
rect 23566 29112 23572 29164
rect 23624 29112 23630 29164
rect 23842 29112 23848 29164
rect 23900 29112 23906 29164
rect 24026 29112 24032 29164
rect 24084 29112 24090 29164
rect 24136 29161 24164 29192
rect 24688 29192 25136 29220
rect 24121 29155 24179 29161
rect 24121 29121 24133 29155
rect 24167 29121 24179 29155
rect 24121 29115 24179 29121
rect 24397 29155 24455 29161
rect 24397 29121 24409 29155
rect 24443 29121 24455 29155
rect 24397 29115 24455 29121
rect 21324 29056 21680 29084
rect 22005 29087 22063 29093
rect 21324 29044 21330 29056
rect 22005 29053 22017 29087
rect 22051 29084 22063 29087
rect 22370 29084 22376 29096
rect 22051 29056 22376 29084
rect 22051 29053 22063 29056
rect 22005 29047 22063 29053
rect 22370 29044 22376 29056
rect 22428 29044 22434 29096
rect 22465 29087 22523 29093
rect 22465 29053 22477 29087
rect 22511 29084 22523 29087
rect 22554 29084 22560 29096
rect 22511 29056 22560 29084
rect 22511 29053 22523 29056
rect 22465 29047 22523 29053
rect 22554 29044 22560 29056
rect 22612 29044 22618 29096
rect 23385 29087 23443 29093
rect 23385 29053 23397 29087
rect 23431 29084 23443 29087
rect 24213 29087 24271 29093
rect 24213 29084 24225 29087
rect 23431 29056 24225 29084
rect 23431 29053 23443 29056
rect 23385 29047 23443 29053
rect 23860 29028 23888 29056
rect 24213 29053 24225 29056
rect 24259 29053 24271 29087
rect 24412 29084 24440 29115
rect 24486 29112 24492 29164
rect 24544 29152 24550 29164
rect 24581 29155 24639 29161
rect 24581 29152 24593 29155
rect 24544 29124 24593 29152
rect 24544 29112 24550 29124
rect 24581 29121 24593 29124
rect 24627 29121 24639 29155
rect 24581 29115 24639 29121
rect 24213 29047 24271 29053
rect 24320 29056 24440 29084
rect 21008 28988 21680 29016
rect 16022 28948 16028 28960
rect 11808 28920 16028 28948
rect 16022 28908 16028 28920
rect 16080 28908 16086 28960
rect 19150 28908 19156 28960
rect 19208 28957 19214 28960
rect 19208 28951 19230 28957
rect 19218 28917 19230 28951
rect 21652 28948 21680 28988
rect 21726 28976 21732 29028
rect 21784 29016 21790 29028
rect 21821 29019 21879 29025
rect 21821 29016 21833 29019
rect 21784 28988 21833 29016
rect 21784 28976 21790 28988
rect 21821 28985 21833 28988
rect 21867 28985 21879 29019
rect 22278 29016 22284 29028
rect 21821 28979 21879 28985
rect 21928 28988 22284 29016
rect 21928 28948 21956 28988
rect 22278 28976 22284 28988
rect 22336 28976 22342 29028
rect 23201 29019 23259 29025
rect 23201 28985 23213 29019
rect 23247 29016 23259 29019
rect 23247 28988 23336 29016
rect 23247 28985 23259 28988
rect 23201 28979 23259 28985
rect 21652 28920 21956 28948
rect 22925 28951 22983 28957
rect 19208 28911 19230 28917
rect 22925 28917 22937 28951
rect 22971 28948 22983 28951
rect 23014 28948 23020 28960
rect 22971 28920 23020 28948
rect 22971 28917 22983 28920
rect 22925 28911 22983 28917
rect 19208 28908 19214 28911
rect 23014 28908 23020 28920
rect 23072 28908 23078 28960
rect 23308 28948 23336 28988
rect 23842 28976 23848 29028
rect 23900 28976 23906 29028
rect 23474 28948 23480 28960
rect 23308 28920 23480 28948
rect 23474 28908 23480 28920
rect 23532 28908 23538 28960
rect 23658 28908 23664 28960
rect 23716 28908 23722 28960
rect 24320 28948 24348 29056
rect 24486 28948 24492 28960
rect 24320 28920 24492 28948
rect 24486 28908 24492 28920
rect 24544 28908 24550 28960
rect 24596 28948 24624 29115
rect 24688 29093 24716 29192
rect 24762 29112 24768 29164
rect 24820 29112 24826 29164
rect 25056 29161 25084 29192
rect 25130 29180 25136 29192
rect 25188 29180 25194 29232
rect 25774 29180 25780 29232
rect 25832 29220 25838 29232
rect 27080 29220 27108 29260
rect 27249 29257 27261 29260
rect 27295 29288 27307 29291
rect 27430 29288 27436 29300
rect 27295 29260 27436 29288
rect 27295 29257 27307 29260
rect 27249 29251 27307 29257
rect 27430 29248 27436 29260
rect 27488 29248 27494 29300
rect 27893 29291 27951 29297
rect 27893 29257 27905 29291
rect 27939 29288 27951 29291
rect 29730 29288 29736 29300
rect 27939 29260 29736 29288
rect 27939 29257 27951 29260
rect 27893 29251 27951 29257
rect 29730 29248 29736 29260
rect 29788 29248 29794 29300
rect 30742 29248 30748 29300
rect 30800 29288 30806 29300
rect 31478 29288 31484 29300
rect 30800 29260 31484 29288
rect 30800 29248 30806 29260
rect 31478 29248 31484 29260
rect 31536 29288 31542 29300
rect 32217 29291 32275 29297
rect 31536 29260 32168 29288
rect 31536 29248 31542 29260
rect 28534 29220 28540 29232
rect 28592 29229 28598 29232
rect 28592 29223 28621 29229
rect 25832 29192 27108 29220
rect 27172 29192 28540 29220
rect 25832 29180 25838 29192
rect 24857 29155 24915 29161
rect 24857 29121 24869 29155
rect 24903 29121 24915 29155
rect 24857 29115 24915 29121
rect 25041 29155 25099 29161
rect 25041 29121 25053 29155
rect 25087 29121 25099 29155
rect 25041 29115 25099 29121
rect 24673 29087 24731 29093
rect 24673 29053 24685 29087
rect 24719 29053 24731 29087
rect 24673 29047 24731 29053
rect 24872 29028 24900 29115
rect 25406 29112 25412 29164
rect 25464 29112 25470 29164
rect 25498 29112 25504 29164
rect 25556 29112 25562 29164
rect 25590 29112 25596 29164
rect 25648 29152 25654 29164
rect 25685 29155 25743 29161
rect 25685 29152 25697 29155
rect 25648 29124 25697 29152
rect 25648 29112 25654 29124
rect 25685 29121 25697 29124
rect 25731 29121 25743 29155
rect 25685 29115 25743 29121
rect 25869 29155 25927 29161
rect 25869 29121 25881 29155
rect 25915 29152 25927 29155
rect 26234 29152 26240 29164
rect 25915 29124 26240 29152
rect 25915 29121 25927 29124
rect 25869 29115 25927 29121
rect 26234 29112 26240 29124
rect 26292 29112 26298 29164
rect 26418 29112 26424 29164
rect 26476 29112 26482 29164
rect 27172 29161 27200 29192
rect 28534 29180 28540 29192
rect 28609 29189 28621 29223
rect 28592 29183 28621 29189
rect 28592 29180 28598 29183
rect 31754 29180 31760 29232
rect 31812 29180 31818 29232
rect 32140 29220 32168 29260
rect 32217 29257 32229 29291
rect 32263 29288 32275 29291
rect 32766 29288 32772 29300
rect 32263 29260 32772 29288
rect 32263 29257 32275 29260
rect 32217 29251 32275 29257
rect 32766 29248 32772 29260
rect 32824 29248 32830 29300
rect 33686 29248 33692 29300
rect 33744 29288 33750 29300
rect 35066 29288 35072 29300
rect 33744 29260 35072 29288
rect 33744 29248 33750 29260
rect 35066 29248 35072 29260
rect 35124 29248 35130 29300
rect 35437 29291 35495 29297
rect 35176 29260 35388 29288
rect 32493 29223 32551 29229
rect 32493 29220 32505 29223
rect 32140 29192 32505 29220
rect 32493 29189 32505 29192
rect 32539 29189 32551 29223
rect 32493 29183 32551 29189
rect 32585 29223 32643 29229
rect 32585 29189 32597 29223
rect 32631 29220 32643 29223
rect 33502 29220 33508 29232
rect 32631 29192 33508 29220
rect 32631 29189 32643 29192
rect 32585 29183 32643 29189
rect 33502 29180 33508 29192
rect 33560 29180 33566 29232
rect 34330 29220 34336 29232
rect 33612 29192 34336 29220
rect 26605 29155 26663 29161
rect 26605 29121 26617 29155
rect 26651 29152 26663 29155
rect 27157 29155 27215 29161
rect 27157 29152 27169 29155
rect 26651 29124 27169 29152
rect 26651 29121 26663 29124
rect 26605 29115 26663 29121
rect 27157 29121 27169 29124
rect 27203 29121 27215 29155
rect 27157 29115 27215 29121
rect 27522 29112 27528 29164
rect 27580 29112 27586 29164
rect 28258 29112 28264 29164
rect 28316 29112 28322 29164
rect 28350 29112 28356 29164
rect 28408 29112 28414 29164
rect 28442 29112 28448 29164
rect 28500 29112 28506 29164
rect 28997 29155 29055 29161
rect 28997 29121 29009 29155
rect 29043 29152 29055 29155
rect 30374 29152 30380 29164
rect 29043 29124 30380 29152
rect 29043 29121 29055 29124
rect 28997 29115 29055 29121
rect 30374 29112 30380 29124
rect 30432 29112 30438 29164
rect 32398 29161 32404 29164
rect 31941 29155 31999 29161
rect 31941 29121 31953 29155
rect 31987 29152 31999 29155
rect 32396 29152 32404 29161
rect 31987 29124 32260 29152
rect 32359 29124 32404 29152
rect 31987 29121 31999 29124
rect 31941 29115 31999 29121
rect 25130 29044 25136 29096
rect 25188 29044 25194 29096
rect 25225 29087 25283 29093
rect 25225 29053 25237 29087
rect 25271 29084 25283 29087
rect 25516 29084 25544 29112
rect 25271 29056 25544 29084
rect 25271 29053 25283 29056
rect 25225 29047 25283 29053
rect 27430 29044 27436 29096
rect 27488 29084 27494 29096
rect 28077 29087 28135 29093
rect 28077 29084 28089 29087
rect 27488 29056 28089 29084
rect 27488 29044 27494 29056
rect 28077 29053 28089 29056
rect 28123 29053 28135 29087
rect 28077 29047 28135 29053
rect 28718 29044 28724 29096
rect 28776 29044 28782 29096
rect 32232 29084 32260 29124
rect 32396 29115 32404 29124
rect 32398 29112 32404 29115
rect 32456 29112 32462 29164
rect 32674 29112 32680 29164
rect 32732 29161 32738 29164
rect 32732 29155 32771 29161
rect 32759 29121 32771 29155
rect 32732 29115 32771 29121
rect 32861 29155 32919 29161
rect 32861 29121 32873 29155
rect 32907 29152 32919 29155
rect 33042 29152 33048 29164
rect 32907 29124 33048 29152
rect 32907 29121 32919 29124
rect 32861 29115 32919 29121
rect 32732 29112 32738 29115
rect 33042 29112 33048 29124
rect 33100 29112 33106 29164
rect 33612 29161 33640 29192
rect 34330 29180 34336 29192
rect 34388 29180 34394 29232
rect 34514 29180 34520 29232
rect 34572 29220 34578 29232
rect 35176 29220 35204 29260
rect 34572 29192 35204 29220
rect 35360 29220 35388 29260
rect 35437 29257 35449 29291
rect 35483 29288 35495 29291
rect 35483 29260 35848 29288
rect 35483 29257 35495 29260
rect 35437 29251 35495 29257
rect 35360 29192 35480 29220
rect 34572 29180 34578 29192
rect 33596 29155 33654 29161
rect 33596 29121 33608 29155
rect 33642 29121 33654 29155
rect 33596 29115 33654 29121
rect 33686 29112 33692 29164
rect 33744 29112 33750 29164
rect 34057 29155 34115 29161
rect 34057 29121 34069 29155
rect 34103 29152 34115 29155
rect 34146 29152 34152 29164
rect 34103 29124 34152 29152
rect 34103 29121 34115 29124
rect 34057 29115 34115 29121
rect 34146 29112 34152 29124
rect 34204 29112 34210 29164
rect 34606 29112 34612 29164
rect 34664 29112 34670 29164
rect 34974 29112 34980 29164
rect 35032 29112 35038 29164
rect 33781 29087 33839 29093
rect 32232 29056 32812 29084
rect 24854 28976 24860 29028
rect 24912 28976 24918 29028
rect 25314 28976 25320 29028
rect 25372 29016 25378 29028
rect 25685 29019 25743 29025
rect 25685 29016 25697 29019
rect 25372 28988 25697 29016
rect 25372 28976 25378 28988
rect 25685 28985 25697 28988
rect 25731 28985 25743 29019
rect 25685 28979 25743 28985
rect 25792 28988 26648 29016
rect 25792 28948 25820 28988
rect 24596 28920 25820 28948
rect 26620 28948 26648 28988
rect 26694 28976 26700 29028
rect 26752 29016 26758 29028
rect 26789 29019 26847 29025
rect 26789 29016 26801 29019
rect 26752 28988 26801 29016
rect 26752 28976 26758 28988
rect 26789 28985 26801 28988
rect 26835 29016 26847 29019
rect 27617 29019 27675 29025
rect 27617 29016 27629 29019
rect 26835 28988 27629 29016
rect 26835 28985 26847 28988
rect 26789 28979 26847 28985
rect 27617 28985 27629 28988
rect 27663 28985 27675 29019
rect 27617 28979 27675 28985
rect 28810 28976 28816 29028
rect 28868 28976 28874 29028
rect 31573 29019 31631 29025
rect 31573 28985 31585 29019
rect 31619 29016 31631 29019
rect 32214 29016 32220 29028
rect 31619 28988 32220 29016
rect 31619 28985 31631 28988
rect 31573 28979 31631 28985
rect 32214 28976 32220 28988
rect 32272 28976 32278 29028
rect 28258 28948 28264 28960
rect 26620 28920 28264 28948
rect 28258 28908 28264 28920
rect 28316 28908 28322 28960
rect 32784 28948 32812 29056
rect 33781 29053 33793 29087
rect 33827 29084 33839 29087
rect 34425 29087 34483 29093
rect 34425 29084 34437 29087
rect 33827 29056 34437 29084
rect 33827 29053 33839 29056
rect 33781 29047 33839 29053
rect 32858 28976 32864 29028
rect 32916 29016 32922 29028
rect 33796 29016 33824 29047
rect 34072 29028 34100 29056
rect 34425 29053 34437 29056
rect 34471 29053 34483 29087
rect 34992 29084 35020 29112
rect 34425 29047 34483 29053
rect 34532 29056 35020 29084
rect 35452 29084 35480 29192
rect 35526 29180 35532 29232
rect 35584 29180 35590 29232
rect 35621 29223 35679 29229
rect 35621 29189 35633 29223
rect 35667 29220 35679 29223
rect 35667 29192 35756 29220
rect 35667 29189 35679 29192
rect 35621 29183 35679 29189
rect 35728 29084 35756 29192
rect 35820 29152 35848 29260
rect 36078 29248 36084 29300
rect 36136 29288 36142 29300
rect 36136 29260 37504 29288
rect 36136 29248 36142 29260
rect 35897 29223 35955 29229
rect 35897 29189 35909 29223
rect 35943 29220 35955 29223
rect 36446 29220 36452 29232
rect 35943 29192 36452 29220
rect 35943 29189 35955 29192
rect 35897 29183 35955 29189
rect 36446 29180 36452 29192
rect 36504 29180 36510 29232
rect 36722 29229 36728 29232
rect 36709 29223 36728 29229
rect 36709 29189 36721 29223
rect 36709 29183 36728 29189
rect 36722 29180 36728 29183
rect 36780 29180 36786 29232
rect 36906 29180 36912 29232
rect 36964 29180 36970 29232
rect 35989 29155 36047 29161
rect 35989 29152 36001 29155
rect 35820 29124 36001 29152
rect 35989 29121 36001 29124
rect 36035 29152 36047 29155
rect 36078 29152 36084 29164
rect 36035 29124 36084 29152
rect 36035 29121 36047 29124
rect 35989 29115 36047 29121
rect 36078 29112 36084 29124
rect 36136 29112 36142 29164
rect 36173 29155 36231 29161
rect 36173 29121 36185 29155
rect 36219 29152 36231 29155
rect 36262 29152 36268 29164
rect 36219 29124 36268 29152
rect 36219 29121 36231 29124
rect 36173 29115 36231 29121
rect 36262 29112 36268 29124
rect 36320 29112 36326 29164
rect 36357 29155 36415 29161
rect 36357 29121 36369 29155
rect 36403 29152 36415 29155
rect 36538 29152 36544 29164
rect 36403 29124 36544 29152
rect 36403 29121 36415 29124
rect 36357 29115 36415 29121
rect 36538 29112 36544 29124
rect 36596 29112 36602 29164
rect 37274 29112 37280 29164
rect 37332 29112 37338 29164
rect 37476 29161 37504 29260
rect 39206 29248 39212 29300
rect 39264 29288 39270 29300
rect 39264 29260 40264 29288
rect 39264 29248 39270 29260
rect 38470 29180 38476 29232
rect 38528 29180 38534 29232
rect 39482 29180 39488 29232
rect 39540 29180 39546 29232
rect 40236 29229 40264 29260
rect 40221 29223 40279 29229
rect 40221 29189 40233 29223
rect 40267 29189 40279 29223
rect 40221 29183 40279 29189
rect 37461 29155 37519 29161
rect 37461 29121 37473 29155
rect 37507 29152 37519 29155
rect 37553 29155 37611 29161
rect 37553 29152 37565 29155
rect 37507 29124 37565 29152
rect 37507 29121 37519 29124
rect 37461 29115 37519 29121
rect 37553 29121 37565 29124
rect 37599 29121 37611 29155
rect 37553 29115 37611 29121
rect 37737 29155 37795 29161
rect 37737 29121 37749 29155
rect 37783 29152 37795 29155
rect 37826 29152 37832 29164
rect 37783 29124 37832 29152
rect 37783 29121 37795 29124
rect 37737 29115 37795 29121
rect 37826 29112 37832 29124
rect 37884 29112 37890 29164
rect 38194 29112 38200 29164
rect 38252 29112 38258 29164
rect 35452 29056 35756 29084
rect 37645 29087 37703 29093
rect 32916 28988 33824 29016
rect 32916 28976 32922 28988
rect 33870 28976 33876 29028
rect 33928 28976 33934 29028
rect 34054 28976 34060 29028
rect 34112 28976 34118 29028
rect 34146 28976 34152 29028
rect 34204 29016 34210 29028
rect 34532 29016 34560 29056
rect 37645 29053 37657 29087
rect 37691 29084 37703 29087
rect 38930 29084 38936 29096
rect 37691 29056 38936 29084
rect 37691 29053 37703 29056
rect 37645 29047 37703 29053
rect 38930 29044 38936 29056
rect 38988 29044 38994 29096
rect 34204 28988 34560 29016
rect 34885 29019 34943 29025
rect 34204 28976 34210 28988
rect 34885 28985 34897 29019
rect 34931 28985 34943 29019
rect 34885 28979 34943 28985
rect 33134 28948 33140 28960
rect 32784 28920 33140 28948
rect 33134 28908 33140 28920
rect 33192 28948 33198 28960
rect 33505 28951 33563 28957
rect 33505 28948 33517 28951
rect 33192 28920 33517 28948
rect 33192 28908 33198 28920
rect 33505 28917 33517 28920
rect 33551 28948 33563 28951
rect 33594 28948 33600 28960
rect 33551 28920 33600 28948
rect 33551 28917 33563 28920
rect 33505 28911 33563 28917
rect 33594 28908 33600 28920
rect 33652 28908 33658 28960
rect 34238 28908 34244 28960
rect 34296 28908 34302 28960
rect 34422 28908 34428 28960
rect 34480 28948 34486 28960
rect 34900 28948 34928 28979
rect 35250 28976 35256 29028
rect 35308 29016 35314 29028
rect 35308 28988 35480 29016
rect 35308 28976 35314 28988
rect 34480 28920 34928 28948
rect 35452 28948 35480 28988
rect 35802 28976 35808 29028
rect 35860 28976 35866 29028
rect 36262 28976 36268 29028
rect 36320 29016 36326 29028
rect 36541 29019 36599 29025
rect 36541 29016 36553 29019
rect 36320 28988 36553 29016
rect 36320 28976 36326 28988
rect 36541 28985 36553 28988
rect 36587 28985 36599 29019
rect 36541 28979 36599 28985
rect 37277 29019 37335 29025
rect 37277 28985 37289 29019
rect 37323 29016 37335 29019
rect 37550 29016 37556 29028
rect 37323 28988 37556 29016
rect 37323 28985 37335 28988
rect 37277 28979 37335 28985
rect 37550 28976 37556 28988
rect 37608 28976 37614 29028
rect 37734 28976 37740 29028
rect 37792 29016 37798 29028
rect 38194 29016 38200 29028
rect 37792 28988 38200 29016
rect 37792 28976 37798 28988
rect 38194 28976 38200 28988
rect 38252 28976 38258 29028
rect 36725 28951 36783 28957
rect 36725 28948 36737 28951
rect 35452 28920 36737 28948
rect 34480 28908 34486 28920
rect 36725 28917 36737 28920
rect 36771 28917 36783 28951
rect 36725 28911 36783 28917
rect 1104 28858 40572 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 40572 28858
rect 1104 28784 40572 28806
rect 6178 28704 6184 28756
rect 6236 28744 6242 28756
rect 6236 28716 6868 28744
rect 6236 28704 6242 28716
rect 6840 28676 6868 28716
rect 7098 28704 7104 28756
rect 7156 28744 7162 28756
rect 7561 28747 7619 28753
rect 7561 28744 7573 28747
rect 7156 28716 7573 28744
rect 7156 28704 7162 28716
rect 7561 28713 7573 28716
rect 7607 28713 7619 28747
rect 11149 28747 11207 28753
rect 7561 28707 7619 28713
rect 7668 28716 11100 28744
rect 7668 28676 7696 28716
rect 6840 28648 7696 28676
rect 9858 28636 9864 28688
rect 9916 28676 9922 28688
rect 10413 28679 10471 28685
rect 10413 28676 10425 28679
rect 9916 28648 10425 28676
rect 9916 28636 9922 28648
rect 10413 28645 10425 28648
rect 10459 28645 10471 28679
rect 11072 28676 11100 28716
rect 11149 28713 11161 28747
rect 11195 28744 11207 28747
rect 11790 28744 11796 28756
rect 11195 28716 11796 28744
rect 11195 28713 11207 28716
rect 11149 28707 11207 28713
rect 11790 28704 11796 28716
rect 11848 28704 11854 28756
rect 11882 28704 11888 28756
rect 11940 28744 11946 28756
rect 12069 28747 12127 28753
rect 12069 28744 12081 28747
rect 11940 28716 12081 28744
rect 11940 28704 11946 28716
rect 12069 28713 12081 28716
rect 12115 28713 12127 28747
rect 12069 28707 12127 28713
rect 14366 28704 14372 28756
rect 14424 28744 14430 28756
rect 16390 28744 16396 28756
rect 14424 28716 16396 28744
rect 14424 28704 14430 28716
rect 16390 28704 16396 28716
rect 16448 28704 16454 28756
rect 20898 28704 20904 28756
rect 20956 28744 20962 28756
rect 21913 28747 21971 28753
rect 21913 28744 21925 28747
rect 20956 28716 21925 28744
rect 20956 28704 20962 28716
rect 21913 28713 21925 28716
rect 21959 28713 21971 28747
rect 21913 28707 21971 28713
rect 24026 28704 24032 28756
rect 24084 28704 24090 28756
rect 24394 28704 24400 28756
rect 24452 28744 24458 28756
rect 24489 28747 24547 28753
rect 24489 28744 24501 28747
rect 24452 28716 24501 28744
rect 24452 28704 24458 28716
rect 24489 28713 24501 28716
rect 24535 28713 24547 28747
rect 24489 28707 24547 28713
rect 26234 28704 26240 28756
rect 26292 28704 26298 28756
rect 26694 28704 26700 28756
rect 26752 28704 26758 28756
rect 27062 28704 27068 28756
rect 27120 28744 27126 28756
rect 29638 28744 29644 28756
rect 27120 28716 29644 28744
rect 27120 28704 27126 28716
rect 29638 28704 29644 28716
rect 29696 28744 29702 28756
rect 29914 28744 29920 28756
rect 29696 28716 29920 28744
rect 29696 28704 29702 28716
rect 29914 28704 29920 28716
rect 29972 28704 29978 28756
rect 32398 28704 32404 28756
rect 32456 28744 32462 28756
rect 32582 28744 32588 28756
rect 32456 28716 32588 28744
rect 32456 28704 32462 28716
rect 32582 28704 32588 28716
rect 32640 28704 32646 28756
rect 34146 28704 34152 28756
rect 34204 28744 34210 28756
rect 34241 28747 34299 28753
rect 34241 28744 34253 28747
rect 34204 28716 34253 28744
rect 34204 28704 34210 28716
rect 34241 28713 34253 28716
rect 34287 28713 34299 28747
rect 34241 28707 34299 28713
rect 34422 28704 34428 28756
rect 34480 28744 34486 28756
rect 35161 28747 35219 28753
rect 35161 28744 35173 28747
rect 34480 28716 35173 28744
rect 34480 28704 34486 28716
rect 35161 28713 35173 28716
rect 35207 28744 35219 28747
rect 36446 28744 36452 28756
rect 35207 28716 36452 28744
rect 35207 28713 35219 28716
rect 35161 28707 35219 28713
rect 36446 28704 36452 28716
rect 36504 28744 36510 28756
rect 38102 28744 38108 28756
rect 36504 28716 38108 28744
rect 36504 28704 36510 28716
rect 38102 28704 38108 28716
rect 38160 28704 38166 28756
rect 38197 28747 38255 28753
rect 38197 28713 38209 28747
rect 38243 28744 38255 28747
rect 38378 28744 38384 28756
rect 38243 28716 38384 28744
rect 38243 28713 38255 28716
rect 38197 28707 38255 28713
rect 38378 28704 38384 28716
rect 38436 28704 38442 28756
rect 11072 28648 12020 28676
rect 10413 28639 10471 28645
rect 5534 28568 5540 28620
rect 5592 28608 5598 28620
rect 6822 28608 6828 28620
rect 5592 28580 6828 28608
rect 5592 28568 5598 28580
rect 6822 28568 6828 28580
rect 6880 28568 6886 28620
rect 8205 28611 8263 28617
rect 8205 28577 8217 28611
rect 8251 28608 8263 28611
rect 8478 28608 8484 28620
rect 8251 28580 8484 28608
rect 8251 28577 8263 28580
rect 8205 28571 8263 28577
rect 8478 28568 8484 28580
rect 8536 28568 8542 28620
rect 10045 28611 10103 28617
rect 10045 28577 10057 28611
rect 10091 28608 10103 28611
rect 10597 28611 10655 28617
rect 10597 28608 10609 28611
rect 10091 28580 10609 28608
rect 10091 28577 10103 28580
rect 10045 28571 10103 28577
rect 10597 28577 10609 28580
rect 10643 28608 10655 28611
rect 10643 28580 11192 28608
rect 10643 28577 10655 28580
rect 10597 28571 10655 28577
rect 8021 28543 8079 28549
rect 8021 28509 8033 28543
rect 8067 28540 8079 28543
rect 8662 28540 8668 28552
rect 8067 28512 8668 28540
rect 8067 28509 8079 28512
rect 8021 28503 8079 28509
rect 8662 28500 8668 28512
rect 8720 28500 8726 28552
rect 9674 28500 9680 28552
rect 9732 28540 9738 28552
rect 9769 28543 9827 28549
rect 9769 28540 9781 28543
rect 9732 28512 9781 28540
rect 9732 28500 9738 28512
rect 9769 28509 9781 28512
rect 9815 28509 9827 28543
rect 9769 28503 9827 28509
rect 10410 28500 10416 28552
rect 10468 28500 10474 28552
rect 10686 28500 10692 28552
rect 10744 28540 10750 28552
rect 11164 28549 11192 28580
rect 11606 28568 11612 28620
rect 11664 28608 11670 28620
rect 11992 28608 12020 28648
rect 13906 28636 13912 28688
rect 13964 28676 13970 28688
rect 15562 28676 15568 28688
rect 13964 28648 15568 28676
rect 13964 28636 13970 28648
rect 15562 28636 15568 28648
rect 15620 28636 15626 28688
rect 17586 28636 17592 28688
rect 17644 28676 17650 28688
rect 23845 28679 23903 28685
rect 23845 28676 23857 28679
rect 17644 28648 23857 28676
rect 17644 28636 17650 28648
rect 14734 28608 14740 28620
rect 11664 28580 11928 28608
rect 11992 28580 14740 28608
rect 11664 28568 11670 28580
rect 10873 28543 10931 28549
rect 10873 28540 10885 28543
rect 10744 28512 10885 28540
rect 10744 28500 10750 28512
rect 10873 28509 10885 28512
rect 10919 28509 10931 28543
rect 10873 28503 10931 28509
rect 11149 28543 11207 28549
rect 11149 28509 11161 28543
rect 11195 28540 11207 28543
rect 11698 28540 11704 28552
rect 11195 28512 11704 28540
rect 11195 28509 11207 28512
rect 11149 28503 11207 28509
rect 11698 28500 11704 28512
rect 11756 28500 11762 28552
rect 11900 28549 11928 28580
rect 14734 28568 14740 28580
rect 14792 28568 14798 28620
rect 16942 28568 16948 28620
rect 17000 28608 17006 28620
rect 17313 28611 17371 28617
rect 17313 28608 17325 28611
rect 17000 28580 17325 28608
rect 17000 28568 17006 28580
rect 17313 28577 17325 28580
rect 17359 28577 17371 28611
rect 17313 28571 17371 28577
rect 11793 28543 11851 28549
rect 11793 28509 11805 28543
rect 11839 28509 11851 28543
rect 11793 28503 11851 28509
rect 11885 28543 11943 28549
rect 11885 28509 11897 28543
rect 11931 28509 11943 28543
rect 11885 28503 11943 28509
rect 12161 28543 12219 28549
rect 12161 28509 12173 28543
rect 12207 28540 12219 28543
rect 12250 28540 12256 28552
rect 12207 28512 12256 28540
rect 12207 28509 12219 28512
rect 12161 28503 12219 28509
rect 3878 28432 3884 28484
rect 3936 28472 3942 28484
rect 4614 28472 4620 28484
rect 3936 28444 4620 28472
rect 3936 28432 3942 28444
rect 4614 28432 4620 28444
rect 4672 28432 4678 28484
rect 5810 28432 5816 28484
rect 5868 28432 5874 28484
rect 9475 28475 9533 28481
rect 9475 28472 9487 28475
rect 5920 28444 6302 28472
rect 7116 28444 9487 28472
rect 4062 28364 4068 28416
rect 4120 28404 4126 28416
rect 5920 28404 5948 28444
rect 4120 28376 5948 28404
rect 4120 28364 4126 28376
rect 6454 28364 6460 28416
rect 6512 28404 6518 28416
rect 7116 28404 7144 28444
rect 9475 28441 9487 28444
rect 9521 28441 9533 28475
rect 9475 28435 9533 28441
rect 10778 28432 10784 28484
rect 10836 28432 10842 28484
rect 11057 28475 11115 28481
rect 11057 28441 11069 28475
rect 11103 28441 11115 28475
rect 11808 28472 11836 28503
rect 12250 28500 12256 28512
rect 12308 28500 12314 28552
rect 13354 28500 13360 28552
rect 13412 28540 13418 28552
rect 14274 28540 14280 28552
rect 13412 28512 14280 28540
rect 13412 28500 13418 28512
rect 14274 28500 14280 28512
rect 14332 28500 14338 28552
rect 14642 28500 14648 28552
rect 14700 28500 14706 28552
rect 17788 28549 17816 28648
rect 23845 28645 23857 28648
rect 23891 28645 23903 28679
rect 24670 28676 24676 28688
rect 23845 28639 23903 28645
rect 24412 28648 24676 28676
rect 17862 28568 17868 28620
rect 17920 28608 17926 28620
rect 23566 28608 23572 28620
rect 17920 28580 22324 28608
rect 17920 28568 17926 28580
rect 17773 28543 17831 28549
rect 17773 28509 17785 28543
rect 17819 28509 17831 28543
rect 17773 28503 17831 28509
rect 21174 28500 21180 28552
rect 21232 28500 21238 28552
rect 21358 28500 21364 28552
rect 21416 28540 21422 28552
rect 22094 28540 22100 28552
rect 21416 28512 22100 28540
rect 21416 28500 21422 28512
rect 22094 28500 22100 28512
rect 22152 28500 22158 28552
rect 22189 28543 22247 28549
rect 22189 28509 22201 28543
rect 22235 28509 22247 28543
rect 22189 28503 22247 28509
rect 12434 28472 12440 28484
rect 11808 28444 12440 28472
rect 11057 28435 11115 28441
rect 6512 28376 7144 28404
rect 6512 28364 6518 28376
rect 7282 28364 7288 28416
rect 7340 28364 7346 28416
rect 7929 28407 7987 28413
rect 7929 28373 7941 28407
rect 7975 28404 7987 28407
rect 8294 28404 8300 28416
rect 7975 28376 8300 28404
rect 7975 28373 7987 28376
rect 7929 28367 7987 28373
rect 8294 28364 8300 28376
rect 8352 28404 8358 28416
rect 8846 28404 8852 28416
rect 8352 28376 8852 28404
rect 8352 28364 8358 28376
rect 8846 28364 8852 28376
rect 8904 28364 8910 28416
rect 9953 28407 10011 28413
rect 9953 28373 9965 28407
rect 9999 28404 10011 28407
rect 10226 28404 10232 28416
rect 9999 28376 10232 28404
rect 9999 28373 10011 28376
rect 9953 28367 10011 28373
rect 10226 28364 10232 28376
rect 10284 28404 10290 28416
rect 11072 28404 11100 28435
rect 12434 28432 12440 28444
rect 12492 28432 12498 28484
rect 14369 28475 14427 28481
rect 14369 28441 14381 28475
rect 14415 28441 14427 28475
rect 14369 28435 14427 28441
rect 14461 28475 14519 28481
rect 14461 28441 14473 28475
rect 14507 28472 14519 28475
rect 15010 28472 15016 28484
rect 14507 28444 15016 28472
rect 14507 28441 14519 28444
rect 14461 28435 14519 28441
rect 10284 28376 11100 28404
rect 11609 28407 11667 28413
rect 10284 28364 10290 28376
rect 11609 28373 11621 28407
rect 11655 28404 11667 28407
rect 11698 28404 11704 28416
rect 11655 28376 11704 28404
rect 11655 28373 11667 28376
rect 11609 28367 11667 28373
rect 11698 28364 11704 28376
rect 11756 28364 11762 28416
rect 11790 28364 11796 28416
rect 11848 28404 11854 28416
rect 12066 28404 12072 28416
rect 11848 28376 12072 28404
rect 11848 28364 11854 28376
rect 12066 28364 12072 28376
rect 12124 28364 12130 28416
rect 14090 28364 14096 28416
rect 14148 28364 14154 28416
rect 14384 28404 14412 28435
rect 15010 28432 15016 28444
rect 15068 28432 15074 28484
rect 16114 28404 16120 28416
rect 14384 28376 16120 28404
rect 16114 28364 16120 28376
rect 16172 28364 16178 28416
rect 20898 28364 20904 28416
rect 20956 28404 20962 28416
rect 20993 28407 21051 28413
rect 20993 28404 21005 28407
rect 20956 28376 21005 28404
rect 20956 28364 20962 28376
rect 20993 28373 21005 28376
rect 21039 28404 21051 28407
rect 21082 28404 21088 28416
rect 21039 28376 21088 28404
rect 21039 28373 21051 28376
rect 20993 28367 21051 28373
rect 21082 28364 21088 28376
rect 21140 28364 21146 28416
rect 22204 28404 22232 28503
rect 22296 28472 22324 28580
rect 22388 28580 23572 28608
rect 22388 28549 22416 28580
rect 23566 28568 23572 28580
rect 23624 28568 23630 28620
rect 23661 28611 23719 28617
rect 23661 28577 23673 28611
rect 23707 28608 23719 28611
rect 24412 28608 24440 28648
rect 24670 28636 24676 28648
rect 24728 28636 24734 28688
rect 24780 28648 26020 28676
rect 23707 28580 24440 28608
rect 23707 28577 23719 28580
rect 23661 28571 23719 28577
rect 24780 28552 24808 28648
rect 25225 28611 25283 28617
rect 25225 28608 25237 28611
rect 24872 28580 25237 28608
rect 22373 28543 22431 28549
rect 22373 28509 22385 28543
rect 22419 28509 22431 28543
rect 22373 28503 22431 28509
rect 22462 28500 22468 28552
rect 22520 28500 22526 28552
rect 23017 28543 23075 28549
rect 23017 28509 23029 28543
rect 23063 28540 23075 28543
rect 23293 28543 23351 28549
rect 23293 28540 23305 28543
rect 23063 28512 23305 28540
rect 23063 28509 23075 28512
rect 23017 28503 23075 28509
rect 23293 28509 23305 28512
rect 23339 28540 23351 28543
rect 23382 28540 23388 28552
rect 23339 28512 23388 28540
rect 23339 28509 23351 28512
rect 23293 28503 23351 28509
rect 23382 28500 23388 28512
rect 23440 28500 23446 28552
rect 23474 28500 23480 28552
rect 23532 28540 23538 28552
rect 23750 28540 23756 28552
rect 23532 28512 23756 28540
rect 23532 28500 23538 28512
rect 23750 28500 23756 28512
rect 23808 28500 23814 28552
rect 24670 28540 24676 28552
rect 24136 28512 24676 28540
rect 24136 28472 24164 28512
rect 24670 28500 24676 28512
rect 24728 28500 24734 28552
rect 24762 28500 24768 28552
rect 24820 28500 24826 28552
rect 24872 28549 24900 28580
rect 25225 28577 25237 28580
rect 25271 28577 25283 28611
rect 25590 28608 25596 28620
rect 25225 28571 25283 28577
rect 25424 28580 25596 28608
rect 24857 28543 24915 28549
rect 24857 28509 24869 28543
rect 24903 28509 24915 28543
rect 24857 28503 24915 28509
rect 24949 28543 25007 28549
rect 24949 28509 24961 28543
rect 24995 28540 25007 28543
rect 25038 28540 25044 28552
rect 24995 28512 25044 28540
rect 24995 28509 25007 28512
rect 24949 28503 25007 28509
rect 25038 28500 25044 28512
rect 25096 28500 25102 28552
rect 25130 28500 25136 28552
rect 25188 28500 25194 28552
rect 25424 28549 25452 28580
rect 25590 28568 25596 28580
rect 25648 28568 25654 28620
rect 25685 28611 25743 28617
rect 25685 28577 25697 28611
rect 25731 28608 25743 28611
rect 25866 28608 25872 28620
rect 25731 28580 25872 28608
rect 25731 28577 25743 28580
rect 25685 28571 25743 28577
rect 25866 28568 25872 28580
rect 25924 28568 25930 28620
rect 25992 28608 26020 28648
rect 26237 28611 26295 28617
rect 25992 28580 26096 28608
rect 25409 28543 25467 28549
rect 25409 28509 25421 28543
rect 25455 28509 25467 28543
rect 25409 28503 25467 28509
rect 25498 28500 25504 28552
rect 25556 28500 25562 28552
rect 25774 28500 25780 28552
rect 25832 28500 25838 28552
rect 25884 28540 25912 28568
rect 26068 28549 26096 28580
rect 26237 28577 26249 28611
rect 26283 28608 26295 28611
rect 26712 28608 26740 28704
rect 27338 28636 27344 28688
rect 27396 28676 27402 28688
rect 38286 28676 38292 28688
rect 27396 28648 28028 28676
rect 27396 28636 27402 28648
rect 26283 28580 26740 28608
rect 26835 28611 26893 28617
rect 26283 28577 26295 28580
rect 26237 28571 26295 28577
rect 26835 28577 26847 28611
rect 26881 28608 26893 28611
rect 27522 28608 27528 28620
rect 26881 28580 27528 28608
rect 26881 28577 26893 28580
rect 26835 28571 26893 28577
rect 27522 28568 27528 28580
rect 27580 28568 27586 28620
rect 26053 28543 26111 28549
rect 25884 28512 26004 28540
rect 22296 28444 24164 28472
rect 24210 28432 24216 28484
rect 24268 28432 24274 28484
rect 25976 28472 26004 28512
rect 26053 28509 26065 28543
rect 26099 28509 26111 28543
rect 26053 28503 26111 28509
rect 26142 28500 26148 28552
rect 26200 28540 26206 28552
rect 26329 28543 26387 28549
rect 26329 28540 26341 28543
rect 26200 28512 26341 28540
rect 26200 28500 26206 28512
rect 26329 28509 26341 28512
rect 26375 28509 26387 28543
rect 26329 28503 26387 28509
rect 26510 28500 26516 28552
rect 26568 28500 26574 28552
rect 26973 28543 27031 28549
rect 26973 28509 26985 28543
rect 27019 28540 27031 28543
rect 27430 28540 27436 28552
rect 27019 28512 27436 28540
rect 27019 28509 27031 28512
rect 26973 28503 27031 28509
rect 27430 28500 27436 28512
rect 27488 28500 27494 28552
rect 27617 28543 27675 28549
rect 27617 28509 27629 28543
rect 27663 28540 27675 28543
rect 27890 28540 27896 28552
rect 27663 28512 27896 28540
rect 27663 28509 27675 28512
rect 27617 28503 27675 28509
rect 27890 28500 27896 28512
rect 27948 28500 27954 28552
rect 28000 28549 28028 28648
rect 28092 28648 38292 28676
rect 27985 28543 28043 28549
rect 27985 28509 27997 28543
rect 28031 28509 28043 28543
rect 27985 28503 28043 28509
rect 28092 28472 28120 28648
rect 38286 28636 38292 28648
rect 38344 28676 38350 28688
rect 38344 28648 38424 28676
rect 38344 28636 38350 28648
rect 31938 28608 31944 28620
rect 30116 28580 31944 28608
rect 28258 28500 28264 28552
rect 28316 28500 28322 28552
rect 28629 28543 28687 28549
rect 28629 28509 28641 28543
rect 28675 28540 28687 28543
rect 28810 28540 28816 28552
rect 28675 28512 28816 28540
rect 28675 28509 28687 28512
rect 28629 28503 28687 28509
rect 28810 28500 28816 28512
rect 28868 28500 28874 28552
rect 29730 28500 29736 28552
rect 29788 28500 29794 28552
rect 29914 28500 29920 28552
rect 29972 28500 29978 28552
rect 30116 28549 30144 28580
rect 31938 28568 31944 28580
rect 31996 28568 32002 28620
rect 32674 28568 32680 28620
rect 32732 28608 32738 28620
rect 32861 28611 32919 28617
rect 32861 28608 32873 28611
rect 32732 28580 32873 28608
rect 32732 28568 32738 28580
rect 32861 28577 32873 28580
rect 32907 28608 32919 28611
rect 32950 28608 32956 28620
rect 32907 28580 32956 28608
rect 32907 28577 32919 28580
rect 32861 28571 32919 28577
rect 32950 28568 32956 28580
rect 33008 28568 33014 28620
rect 35434 28568 35440 28620
rect 35492 28608 35498 28620
rect 35802 28608 35808 28620
rect 35492 28580 35808 28608
rect 35492 28568 35498 28580
rect 35802 28568 35808 28580
rect 35860 28568 35866 28620
rect 38396 28617 38424 28648
rect 38381 28611 38439 28617
rect 38381 28577 38393 28611
rect 38427 28577 38439 28611
rect 38381 28571 38439 28577
rect 38838 28568 38844 28620
rect 38896 28608 38902 28620
rect 39758 28608 39764 28620
rect 38896 28580 39764 28608
rect 38896 28568 38902 28580
rect 39758 28568 39764 28580
rect 39816 28568 39822 28620
rect 30101 28543 30159 28549
rect 30101 28509 30113 28543
rect 30147 28509 30159 28543
rect 30101 28503 30159 28509
rect 30193 28543 30251 28549
rect 30193 28509 30205 28543
rect 30239 28509 30251 28543
rect 32125 28543 32183 28549
rect 32125 28540 32137 28543
rect 30193 28503 30251 28509
rect 30300 28512 32137 28540
rect 24412 28444 25912 28472
rect 25976 28444 28120 28472
rect 22646 28404 22652 28416
rect 22204 28376 22652 28404
rect 22646 28364 22652 28376
rect 22704 28364 22710 28416
rect 23106 28364 23112 28416
rect 23164 28364 23170 28416
rect 23385 28407 23443 28413
rect 23385 28373 23397 28407
rect 23431 28404 23443 28407
rect 23750 28404 23756 28416
rect 23431 28376 23756 28404
rect 23431 28373 23443 28376
rect 23385 28367 23443 28373
rect 23750 28364 23756 28376
rect 23808 28364 23814 28416
rect 24013 28407 24071 28413
rect 24013 28373 24025 28407
rect 24059 28404 24071 28407
rect 24412 28404 24440 28444
rect 25884 28413 25912 28444
rect 29270 28432 29276 28484
rect 29328 28472 29334 28484
rect 29328 28444 29776 28472
rect 29328 28432 29334 28444
rect 24059 28376 24440 28404
rect 25869 28407 25927 28413
rect 24059 28373 24071 28376
rect 24013 28367 24071 28373
rect 25869 28373 25881 28407
rect 25915 28373 25927 28407
rect 25869 28367 25927 28373
rect 26510 28364 26516 28416
rect 26568 28364 26574 28416
rect 28534 28364 28540 28416
rect 28592 28364 28598 28416
rect 29178 28364 29184 28416
rect 29236 28404 29242 28416
rect 29549 28407 29607 28413
rect 29549 28404 29561 28407
rect 29236 28376 29561 28404
rect 29236 28364 29242 28376
rect 29549 28373 29561 28376
rect 29595 28373 29607 28407
rect 29748 28404 29776 28444
rect 29822 28432 29828 28484
rect 29880 28432 29886 28484
rect 30006 28432 30012 28484
rect 30064 28472 30070 28484
rect 30208 28472 30236 28503
rect 30064 28444 30236 28472
rect 30064 28432 30070 28444
rect 30300 28404 30328 28512
rect 32125 28509 32137 28512
rect 32171 28509 32183 28543
rect 32125 28503 32183 28509
rect 30469 28475 30527 28481
rect 30469 28441 30481 28475
rect 30515 28472 30527 28475
rect 30650 28472 30656 28484
rect 30515 28444 30656 28472
rect 30515 28441 30527 28444
rect 30469 28435 30527 28441
rect 30650 28432 30656 28444
rect 30708 28432 30714 28484
rect 32140 28472 32168 28503
rect 32214 28500 32220 28552
rect 32272 28540 32278 28552
rect 32582 28540 32588 28552
rect 32272 28512 32588 28540
rect 32272 28500 32278 28512
rect 32582 28500 32588 28512
rect 32640 28500 32646 28552
rect 33594 28500 33600 28552
rect 33652 28500 33658 28552
rect 33873 28543 33931 28549
rect 33873 28509 33885 28543
rect 33919 28540 33931 28543
rect 34238 28540 34244 28552
rect 33919 28512 34244 28540
rect 33919 28509 33931 28512
rect 33873 28503 33931 28509
rect 34238 28500 34244 28512
rect 34296 28500 34302 28552
rect 35526 28500 35532 28552
rect 35584 28540 35590 28552
rect 35713 28543 35771 28549
rect 35713 28540 35725 28543
rect 35584 28512 35725 28540
rect 35584 28500 35590 28512
rect 35713 28509 35725 28512
rect 35759 28509 35771 28543
rect 35713 28503 35771 28509
rect 35986 28500 35992 28552
rect 36044 28500 36050 28552
rect 38010 28500 38016 28552
rect 38068 28540 38074 28552
rect 38473 28543 38531 28549
rect 38473 28540 38485 28543
rect 38068 28512 38485 28540
rect 38068 28500 38074 28512
rect 38473 28509 38485 28512
rect 38519 28540 38531 28543
rect 39206 28540 39212 28552
rect 38519 28512 39212 28540
rect 38519 28509 38531 28512
rect 38473 28503 38531 28509
rect 39206 28500 39212 28512
rect 39264 28500 39270 28552
rect 33502 28472 33508 28484
rect 32140 28444 33508 28472
rect 33502 28432 33508 28444
rect 33560 28432 33566 28484
rect 33686 28432 33692 28484
rect 33744 28472 33750 28484
rect 34149 28475 34207 28481
rect 34149 28472 34161 28475
rect 33744 28444 34161 28472
rect 33744 28432 33750 28444
rect 34149 28441 34161 28444
rect 34195 28441 34207 28475
rect 34149 28435 34207 28441
rect 34330 28432 34336 28484
rect 34388 28472 34394 28484
rect 35161 28475 35219 28481
rect 35161 28472 35173 28475
rect 34388 28444 35173 28472
rect 34388 28432 34394 28444
rect 35161 28441 35173 28444
rect 35207 28441 35219 28475
rect 35161 28435 35219 28441
rect 35345 28475 35403 28481
rect 35345 28441 35357 28475
rect 35391 28472 35403 28475
rect 36170 28472 36176 28484
rect 35391 28444 36176 28472
rect 35391 28441 35403 28444
rect 35345 28435 35403 28441
rect 36170 28432 36176 28444
rect 36228 28432 36234 28484
rect 38102 28432 38108 28484
rect 38160 28472 38166 28484
rect 38749 28475 38807 28481
rect 38749 28472 38761 28475
rect 38160 28444 38761 28472
rect 38160 28432 38166 28444
rect 38749 28441 38761 28444
rect 38795 28441 38807 28475
rect 38749 28435 38807 28441
rect 29748 28376 30328 28404
rect 29549 28367 29607 28373
rect 30374 28364 30380 28416
rect 30432 28404 30438 28416
rect 30561 28407 30619 28413
rect 30561 28404 30573 28407
rect 30432 28376 30573 28404
rect 30432 28364 30438 28376
rect 30561 28373 30573 28376
rect 30607 28373 30619 28407
rect 30561 28367 30619 28373
rect 33410 28364 33416 28416
rect 33468 28404 33474 28416
rect 33597 28407 33655 28413
rect 33597 28404 33609 28407
rect 33468 28376 33609 28404
rect 33468 28364 33474 28376
rect 33597 28373 33609 28376
rect 33643 28373 33655 28407
rect 33597 28367 33655 28373
rect 34238 28364 34244 28416
rect 34296 28404 34302 28416
rect 34977 28407 35035 28413
rect 34977 28404 34989 28407
rect 34296 28376 34989 28404
rect 34296 28364 34302 28376
rect 34977 28373 34989 28376
rect 35023 28373 35035 28407
rect 34977 28367 35035 28373
rect 35618 28364 35624 28416
rect 35676 28404 35682 28416
rect 35897 28407 35955 28413
rect 35897 28404 35909 28407
rect 35676 28376 35909 28404
rect 35676 28364 35682 28376
rect 35897 28373 35909 28376
rect 35943 28404 35955 28407
rect 36078 28404 36084 28416
rect 35943 28376 36084 28404
rect 35943 28373 35955 28376
rect 35897 28367 35955 28373
rect 36078 28364 36084 28376
rect 36136 28364 36142 28416
rect 1104 28314 40572 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 40572 28314
rect 1104 28240 40572 28262
rect 4249 28203 4307 28209
rect 4249 28169 4261 28203
rect 4295 28169 4307 28203
rect 4249 28163 4307 28169
rect 4062 28132 4068 28144
rect 4002 28104 4068 28132
rect 4062 28092 4068 28104
rect 4120 28092 4126 28144
rect 4264 28132 4292 28163
rect 5810 28160 5816 28212
rect 5868 28200 5874 28212
rect 6365 28203 6423 28209
rect 6365 28200 6377 28203
rect 5868 28172 6377 28200
rect 5868 28160 5874 28172
rect 6365 28169 6377 28172
rect 6411 28169 6423 28203
rect 6365 28163 6423 28169
rect 6454 28160 6460 28212
rect 6512 28200 6518 28212
rect 14642 28200 14648 28212
rect 6512 28172 14648 28200
rect 6512 28160 6518 28172
rect 14642 28160 14648 28172
rect 14700 28160 14706 28212
rect 14826 28200 14832 28212
rect 14752 28172 14832 28200
rect 4801 28135 4859 28141
rect 4801 28132 4813 28135
rect 4264 28104 4813 28132
rect 4801 28101 4813 28104
rect 4847 28132 4859 28135
rect 5994 28132 6000 28144
rect 4847 28104 6000 28132
rect 4847 28101 4859 28104
rect 4801 28095 4859 28101
rect 5994 28092 6000 28104
rect 6052 28092 6058 28144
rect 6546 28132 6552 28144
rect 6472 28104 6552 28132
rect 4706 28024 4712 28076
rect 4764 28064 4770 28076
rect 6362 28064 6368 28076
rect 4764 28036 6368 28064
rect 4764 28024 4770 28036
rect 6362 28024 6368 28036
rect 6420 28024 6426 28076
rect 2501 27999 2559 28005
rect 2501 27965 2513 27999
rect 2547 27965 2559 27999
rect 2501 27959 2559 27965
rect 2777 27999 2835 28005
rect 2777 27965 2789 27999
rect 2823 27996 2835 27999
rect 4985 27999 5043 28005
rect 2823 27968 4384 27996
rect 2823 27965 2835 27968
rect 2777 27959 2835 27965
rect 2516 27860 2544 27959
rect 4356 27937 4384 27968
rect 4985 27965 4997 27999
rect 5031 27996 5043 27999
rect 6472 27996 6500 28104
rect 6546 28092 6552 28104
rect 6604 28132 6610 28144
rect 6604 28104 7052 28132
rect 6604 28092 6610 28104
rect 6733 28067 6791 28073
rect 6733 28033 6745 28067
rect 6779 28064 6791 28067
rect 6779 28036 6960 28064
rect 6779 28033 6791 28036
rect 6733 28027 6791 28033
rect 5031 27968 6500 27996
rect 6825 27999 6883 28005
rect 5031 27965 5043 27968
rect 4985 27959 5043 27965
rect 6825 27965 6837 27999
rect 6871 27965 6883 27999
rect 6825 27959 6883 27965
rect 4341 27931 4399 27937
rect 4341 27897 4353 27931
rect 4387 27897 4399 27931
rect 4341 27891 4399 27897
rect 4614 27888 4620 27940
rect 4672 27928 4678 27940
rect 5000 27928 5028 27959
rect 4672 27900 5028 27928
rect 4672 27888 4678 27900
rect 3786 27860 3792 27872
rect 2516 27832 3792 27860
rect 3786 27820 3792 27832
rect 3844 27820 3850 27872
rect 6840 27860 6868 27959
rect 6932 27928 6960 28036
rect 7024 28005 7052 28104
rect 7098 28092 7104 28144
rect 7156 28132 7162 28144
rect 7156 28104 13676 28132
rect 7156 28092 7162 28104
rect 9858 28064 9864 28076
rect 8588 28036 9864 28064
rect 7009 27999 7067 28005
rect 7009 27965 7021 27999
rect 7055 27996 7067 27999
rect 8478 27996 8484 28008
rect 7055 27968 8484 27996
rect 7055 27965 7067 27968
rect 7009 27959 7067 27965
rect 8478 27956 8484 27968
rect 8536 27956 8542 28008
rect 7558 27928 7564 27940
rect 6932 27900 7564 27928
rect 7558 27888 7564 27900
rect 7616 27928 7622 27940
rect 8588 27928 8616 28036
rect 9858 28024 9864 28036
rect 9916 28024 9922 28076
rect 11146 28024 11152 28076
rect 11204 28064 11210 28076
rect 11330 28064 11336 28076
rect 11204 28036 11336 28064
rect 11204 28024 11210 28036
rect 11330 28024 11336 28036
rect 11388 28024 11394 28076
rect 11698 28024 11704 28076
rect 11756 28024 11762 28076
rect 11790 28024 11796 28076
rect 11848 28064 11854 28076
rect 11885 28067 11943 28073
rect 11885 28064 11897 28067
rect 11848 28036 11897 28064
rect 11848 28024 11854 28036
rect 11885 28033 11897 28036
rect 11931 28033 11943 28067
rect 11885 28027 11943 28033
rect 12069 28067 12127 28073
rect 12069 28033 12081 28067
rect 12115 28064 12127 28067
rect 12618 28064 12624 28076
rect 12115 28036 12624 28064
rect 12115 28033 12127 28036
rect 12069 28027 12127 28033
rect 12618 28024 12624 28036
rect 12676 28024 12682 28076
rect 12710 28024 12716 28076
rect 12768 28064 12774 28076
rect 13354 28073 13360 28076
rect 12805 28067 12863 28073
rect 12805 28064 12817 28067
rect 12768 28036 12817 28064
rect 12768 28024 12774 28036
rect 12805 28033 12817 28036
rect 12851 28033 12863 28067
rect 12805 28027 12863 28033
rect 12898 28067 12956 28073
rect 12898 28033 12910 28067
rect 12944 28033 12956 28067
rect 12898 28027 12956 28033
rect 13081 28067 13139 28073
rect 13081 28033 13093 28067
rect 13127 28033 13139 28067
rect 13081 28027 13139 28033
rect 13173 28067 13231 28073
rect 13173 28033 13185 28067
rect 13219 28033 13231 28067
rect 13173 28027 13231 28033
rect 13311 28067 13360 28073
rect 13311 28033 13323 28067
rect 13357 28033 13360 28067
rect 13311 28027 13360 28033
rect 8846 27956 8852 28008
rect 8904 27996 8910 28008
rect 12912 27996 12940 28027
rect 8904 27968 12940 27996
rect 8904 27956 8910 27968
rect 7616 27900 8616 27928
rect 7616 27888 7622 27900
rect 9674 27888 9680 27940
rect 9732 27928 9738 27940
rect 11701 27931 11759 27937
rect 11701 27928 11713 27931
rect 9732 27900 11713 27928
rect 9732 27888 9738 27900
rect 11701 27897 11713 27900
rect 11747 27897 11759 27931
rect 13096 27928 13124 28027
rect 13188 27996 13216 28027
rect 13354 28024 13360 28027
rect 13412 28024 13418 28076
rect 13538 28024 13544 28076
rect 13596 28024 13602 28076
rect 13648 28073 13676 28104
rect 13906 28092 13912 28144
rect 13964 28092 13970 28144
rect 14553 28135 14611 28141
rect 14553 28101 14565 28135
rect 14599 28132 14611 28135
rect 14752 28132 14780 28172
rect 14826 28160 14832 28172
rect 14884 28160 14890 28212
rect 15010 28160 15016 28212
rect 15068 28200 15074 28212
rect 15470 28200 15476 28212
rect 15068 28172 15476 28200
rect 15068 28160 15074 28172
rect 15470 28160 15476 28172
rect 15528 28200 15534 28212
rect 15528 28172 19288 28200
rect 15528 28160 15534 28172
rect 15672 28141 15700 28172
rect 14599 28104 14780 28132
rect 15657 28135 15715 28141
rect 14599 28101 14611 28104
rect 14553 28095 14611 28101
rect 15657 28101 15669 28135
rect 15703 28101 15715 28135
rect 15657 28095 15715 28101
rect 15746 28092 15752 28144
rect 15804 28092 15810 28144
rect 16022 28092 16028 28144
rect 16080 28132 16086 28144
rect 16960 28141 16988 28172
rect 16945 28135 17003 28141
rect 16080 28104 16804 28132
rect 16080 28092 16086 28104
rect 13634 28067 13692 28073
rect 13634 28033 13646 28067
rect 13680 28033 13692 28067
rect 13634 28027 13692 28033
rect 13814 28024 13820 28076
rect 13872 28024 13878 28076
rect 14047 28067 14105 28073
rect 14047 28033 14059 28067
rect 14093 28064 14105 28067
rect 14274 28064 14280 28076
rect 14093 28036 14280 28064
rect 14093 28033 14105 28036
rect 14047 28027 14105 28033
rect 14274 28024 14280 28036
rect 14332 28064 14338 28076
rect 14456 28067 14514 28073
rect 14456 28064 14468 28067
rect 14332 28036 14468 28064
rect 14332 28024 14338 28036
rect 14456 28033 14468 28036
rect 14502 28033 14514 28067
rect 14456 28027 14514 28033
rect 14645 28067 14703 28073
rect 14645 28033 14657 28067
rect 14691 28033 14703 28067
rect 14645 28027 14703 28033
rect 14366 27996 14372 28008
rect 13188 27968 14372 27996
rect 14366 27956 14372 27968
rect 14424 27956 14430 28008
rect 13814 27928 13820 27940
rect 13096 27900 13820 27928
rect 11701 27891 11759 27897
rect 13814 27888 13820 27900
rect 13872 27888 13878 27940
rect 13906 27888 13912 27940
rect 13964 27928 13970 27940
rect 14185 27931 14243 27937
rect 14185 27928 14197 27931
rect 13964 27900 14197 27928
rect 13964 27888 13970 27900
rect 14185 27897 14197 27900
rect 14231 27897 14243 27931
rect 14471 27928 14499 28027
rect 14550 27956 14556 28008
rect 14608 27996 14614 28008
rect 14660 27996 14688 28027
rect 14734 28024 14740 28076
rect 14792 28073 14798 28076
rect 14792 28067 14841 28073
rect 14792 28033 14795 28067
rect 14829 28033 14841 28067
rect 14792 28027 14841 28033
rect 14921 28067 14979 28073
rect 14921 28033 14933 28067
rect 14967 28064 14979 28067
rect 15194 28064 15200 28076
rect 14967 28036 15200 28064
rect 14967 28033 14979 28036
rect 14921 28027 14979 28033
rect 14792 28024 14798 28027
rect 15194 28024 15200 28036
rect 15252 28064 15258 28076
rect 15381 28067 15439 28073
rect 15381 28064 15393 28067
rect 15252 28036 15393 28064
rect 15252 28024 15258 28036
rect 15381 28033 15393 28036
rect 15427 28033 15439 28067
rect 15381 28027 15439 28033
rect 15474 28067 15532 28073
rect 15474 28033 15486 28067
rect 15520 28033 15532 28067
rect 15474 28027 15532 28033
rect 15865 28067 15923 28073
rect 15865 28033 15877 28067
rect 15911 28033 15923 28067
rect 15865 28027 15923 28033
rect 15010 27996 15016 28008
rect 14608 27968 15016 27996
rect 14608 27956 14614 27968
rect 15010 27956 15016 27968
rect 15068 27956 15074 28008
rect 14734 27928 14740 27940
rect 14471 27900 14740 27928
rect 14185 27891 14243 27897
rect 14734 27888 14740 27900
rect 14792 27888 14798 27940
rect 6914 27860 6920 27872
rect 6840 27832 6920 27860
rect 6914 27820 6920 27832
rect 6972 27860 6978 27872
rect 7282 27860 7288 27872
rect 6972 27832 7288 27860
rect 6972 27820 6978 27832
rect 7282 27820 7288 27832
rect 7340 27860 7346 27872
rect 12526 27860 12532 27872
rect 7340 27832 12532 27860
rect 7340 27820 7346 27832
rect 12526 27820 12532 27832
rect 12584 27820 12590 27872
rect 13449 27863 13507 27869
rect 13449 27829 13461 27863
rect 13495 27860 13507 27863
rect 13998 27860 14004 27872
rect 13495 27832 14004 27860
rect 13495 27829 13507 27832
rect 13449 27823 13507 27829
rect 13998 27820 14004 27832
rect 14056 27820 14062 27872
rect 14274 27820 14280 27872
rect 14332 27820 14338 27872
rect 14366 27820 14372 27872
rect 14424 27860 14430 27872
rect 15489 27860 15517 28027
rect 15746 27956 15752 28008
rect 15804 27996 15810 28008
rect 15892 27996 15920 28027
rect 16666 28024 16672 28076
rect 16724 28024 16730 28076
rect 16776 28073 16804 28104
rect 16945 28101 16957 28135
rect 16991 28101 17003 28135
rect 16945 28095 17003 28101
rect 17037 28135 17095 28141
rect 17037 28101 17049 28135
rect 17083 28132 17095 28135
rect 17494 28132 17500 28144
rect 17083 28104 17500 28132
rect 17083 28101 17095 28104
rect 17037 28095 17095 28101
rect 17494 28092 17500 28104
rect 17552 28092 17558 28144
rect 19260 28141 19288 28172
rect 19352 28172 22232 28200
rect 19245 28135 19303 28141
rect 19245 28101 19257 28135
rect 19291 28101 19303 28135
rect 19245 28095 19303 28101
rect 16762 28067 16820 28073
rect 16762 28033 16774 28067
rect 16808 28033 16820 28067
rect 16762 28027 16820 28033
rect 17175 28067 17233 28073
rect 17175 28033 17187 28067
rect 17221 28064 17233 28067
rect 17678 28064 17684 28076
rect 17221 28036 17684 28064
rect 17221 28033 17233 28036
rect 17175 28027 17233 28033
rect 17190 27996 17218 28027
rect 17678 28024 17684 28036
rect 17736 28024 17742 28076
rect 18417 28067 18475 28073
rect 18417 28033 18429 28067
rect 18463 28033 18475 28067
rect 18417 28027 18475 28033
rect 18601 28067 18659 28073
rect 18601 28033 18613 28067
rect 18647 28064 18659 28067
rect 18877 28067 18935 28073
rect 18647 28036 18828 28064
rect 18647 28033 18659 28036
rect 18601 28027 18659 28033
rect 15804 27968 17218 27996
rect 15804 27956 15810 27968
rect 18138 27956 18144 28008
rect 18196 27996 18202 28008
rect 18233 27999 18291 28005
rect 18233 27996 18245 27999
rect 18196 27968 18245 27996
rect 18196 27956 18202 27968
rect 18233 27965 18245 27968
rect 18279 27965 18291 27999
rect 18432 27996 18460 28027
rect 18690 27996 18696 28008
rect 18432 27968 18696 27996
rect 18233 27959 18291 27965
rect 18690 27956 18696 27968
rect 18748 27956 18754 28008
rect 18800 27928 18828 28036
rect 18877 28033 18889 28067
rect 18923 28033 18935 28067
rect 18877 28027 18935 28033
rect 19061 28067 19119 28073
rect 19061 28033 19073 28067
rect 19107 28064 19119 28067
rect 19352 28064 19380 28172
rect 19426 28092 19432 28144
rect 19484 28132 19490 28144
rect 19484 28104 19840 28132
rect 19484 28092 19490 28104
rect 19107 28036 19380 28064
rect 19521 28067 19579 28073
rect 19107 28033 19119 28036
rect 19061 28027 19119 28033
rect 18892 27996 18920 28027
rect 19260 28008 19288 28036
rect 19521 28033 19533 28067
rect 19567 28064 19579 28067
rect 19702 28064 19708 28076
rect 19567 28036 19708 28064
rect 19567 28033 19579 28036
rect 19521 28027 19579 28033
rect 19702 28024 19708 28036
rect 19760 28024 19766 28076
rect 19812 28073 19840 28104
rect 19996 28073 20024 28172
rect 21269 28135 21327 28141
rect 21269 28132 21281 28135
rect 20640 28104 21281 28132
rect 20640 28073 20668 28104
rect 21269 28101 21281 28104
rect 21315 28132 21327 28135
rect 21450 28132 21456 28144
rect 21315 28104 21456 28132
rect 21315 28101 21327 28104
rect 21269 28095 21327 28101
rect 21450 28092 21456 28104
rect 21508 28092 21514 28144
rect 19797 28067 19855 28073
rect 19797 28033 19809 28067
rect 19843 28033 19855 28067
rect 19797 28027 19855 28033
rect 19981 28067 20039 28073
rect 19981 28033 19993 28067
rect 20027 28033 20039 28067
rect 19981 28027 20039 28033
rect 20165 28067 20223 28073
rect 20165 28033 20177 28067
rect 20211 28033 20223 28067
rect 20165 28027 20223 28033
rect 20625 28067 20683 28073
rect 20625 28033 20637 28067
rect 20671 28033 20683 28067
rect 20625 28027 20683 28033
rect 21361 28067 21419 28073
rect 21361 28033 21373 28067
rect 21407 28064 21419 28067
rect 21634 28064 21640 28076
rect 21407 28036 21640 28064
rect 21407 28033 21419 28036
rect 21361 28027 21419 28033
rect 19150 27996 19156 28008
rect 18892 27968 19156 27996
rect 19150 27956 19156 27968
rect 19208 27956 19214 28008
rect 19242 27956 19248 28008
rect 19300 27956 19306 28008
rect 19429 27999 19487 28005
rect 19429 27965 19441 27999
rect 19475 27996 19487 27999
rect 19610 27996 19616 28008
rect 19475 27968 19616 27996
rect 19475 27965 19487 27968
rect 19429 27959 19487 27965
rect 19610 27956 19616 27968
rect 19668 27996 19674 28008
rect 20073 27999 20131 28005
rect 20073 27996 20085 27999
rect 19668 27968 20085 27996
rect 19668 27956 19674 27968
rect 20073 27965 20085 27968
rect 20119 27965 20131 27999
rect 20073 27959 20131 27965
rect 19518 27928 19524 27940
rect 18800 27900 19524 27928
rect 19518 27888 19524 27900
rect 19576 27888 19582 27940
rect 14424 27832 15517 27860
rect 16025 27863 16083 27869
rect 14424 27820 14430 27832
rect 16025 27829 16037 27863
rect 16071 27860 16083 27863
rect 16114 27860 16120 27872
rect 16071 27832 16120 27860
rect 16071 27829 16083 27832
rect 16025 27823 16083 27829
rect 16114 27820 16120 27832
rect 16172 27820 16178 27872
rect 17310 27820 17316 27872
rect 17368 27820 17374 27872
rect 17402 27820 17408 27872
rect 17460 27860 17466 27872
rect 17862 27860 17868 27872
rect 17460 27832 17868 27860
rect 17460 27820 17466 27832
rect 17862 27820 17868 27832
rect 17920 27860 17926 27872
rect 18693 27863 18751 27869
rect 18693 27860 18705 27863
rect 17920 27832 18705 27860
rect 17920 27820 17926 27832
rect 18693 27829 18705 27832
rect 18739 27829 18751 27863
rect 18693 27823 18751 27829
rect 19150 27820 19156 27872
rect 19208 27860 19214 27872
rect 20180 27860 20208 28027
rect 21634 28024 21640 28036
rect 21692 28024 21698 28076
rect 21818 28024 21824 28076
rect 21876 28024 21882 28076
rect 22094 28024 22100 28076
rect 22152 28024 22158 28076
rect 20806 27956 20812 28008
rect 20864 27996 20870 28008
rect 21450 27996 21456 28008
rect 20864 27968 21456 27996
rect 20864 27956 20870 27968
rect 21450 27956 21456 27968
rect 21508 27956 21514 28008
rect 22204 28005 22232 28172
rect 25406 28160 25412 28212
rect 25464 28160 25470 28212
rect 25498 28160 25504 28212
rect 25556 28200 25562 28212
rect 25777 28203 25835 28209
rect 25777 28200 25789 28203
rect 25556 28172 25789 28200
rect 25556 28160 25562 28172
rect 25777 28169 25789 28172
rect 25823 28169 25835 28203
rect 25777 28163 25835 28169
rect 32490 28160 32496 28212
rect 32548 28160 32554 28212
rect 24762 28132 24768 28144
rect 22848 28104 24768 28132
rect 22373 28067 22431 28073
rect 22373 28033 22385 28067
rect 22419 28033 22431 28067
rect 22373 28027 22431 28033
rect 21545 27999 21603 28005
rect 21545 27965 21557 27999
rect 21591 27965 21603 27999
rect 21545 27959 21603 27965
rect 22189 27999 22247 28005
rect 22189 27965 22201 27999
rect 22235 27965 22247 27999
rect 22388 27996 22416 28027
rect 22462 28024 22468 28076
rect 22520 28064 22526 28076
rect 22557 28067 22615 28073
rect 22557 28064 22569 28067
rect 22520 28036 22569 28064
rect 22520 28024 22526 28036
rect 22557 28033 22569 28036
rect 22603 28033 22615 28067
rect 22557 28027 22615 28033
rect 22738 28024 22744 28076
rect 22796 28064 22802 28076
rect 22848 28073 22876 28104
rect 24762 28092 24768 28104
rect 24820 28092 24826 28144
rect 30098 28092 30104 28144
rect 30156 28092 30162 28144
rect 30834 28092 30840 28144
rect 30892 28092 30898 28144
rect 31386 28092 31392 28144
rect 31444 28092 31450 28144
rect 22833 28067 22891 28073
rect 22833 28064 22845 28067
rect 22796 28036 22845 28064
rect 22796 28024 22802 28036
rect 22833 28033 22845 28036
rect 22879 28033 22891 28067
rect 22833 28027 22891 28033
rect 23014 28024 23020 28076
rect 23072 28024 23078 28076
rect 25133 28067 25191 28073
rect 25133 28033 25145 28067
rect 25179 28064 25191 28067
rect 26050 28064 26056 28076
rect 25179 28036 26056 28064
rect 25179 28033 25191 28036
rect 25133 28027 25191 28033
rect 26050 28024 26056 28036
rect 26108 28024 26114 28076
rect 28813 28067 28871 28073
rect 28813 28033 28825 28067
rect 28859 28064 28871 28067
rect 28859 28036 29316 28064
rect 28859 28033 28871 28036
rect 28813 28027 28871 28033
rect 23658 27996 23664 28008
rect 22388 27968 23664 27996
rect 22189 27959 22247 27965
rect 20346 27888 20352 27940
rect 20404 27928 20410 27940
rect 20901 27931 20959 27937
rect 20901 27928 20913 27931
rect 20404 27900 20913 27928
rect 20404 27888 20410 27900
rect 20901 27897 20913 27900
rect 20947 27897 20959 27931
rect 20901 27891 20959 27897
rect 21082 27888 21088 27940
rect 21140 27928 21146 27940
rect 21560 27928 21588 27959
rect 23658 27956 23664 27968
rect 23716 27956 23722 28008
rect 23750 27956 23756 28008
rect 23808 27996 23814 28008
rect 25501 27999 25559 28005
rect 25501 27996 25513 27999
rect 23808 27968 25513 27996
rect 23808 27956 23814 27968
rect 25501 27965 25513 27968
rect 25547 27965 25559 27999
rect 25501 27959 25559 27965
rect 25618 27999 25676 28005
rect 25618 27965 25630 27999
rect 25664 27996 25676 27999
rect 25774 27996 25780 28008
rect 25664 27968 25780 27996
rect 25664 27965 25676 27968
rect 25618 27959 25676 27965
rect 22738 27928 22744 27940
rect 21140 27900 22744 27928
rect 21140 27888 21146 27900
rect 22738 27888 22744 27900
rect 22796 27888 22802 27940
rect 25516 27928 25544 27959
rect 25774 27956 25780 27968
rect 25832 27956 25838 28008
rect 29178 27956 29184 28008
rect 29236 27956 29242 28008
rect 29288 27996 29316 28036
rect 30742 28024 30748 28076
rect 30800 28064 30806 28076
rect 31297 28067 31355 28073
rect 31297 28064 31309 28067
rect 30800 28036 31309 28064
rect 30800 28024 30806 28036
rect 31297 28033 31309 28036
rect 31343 28064 31355 28067
rect 32309 28067 32367 28073
rect 31343 28036 31754 28064
rect 31343 28033 31355 28036
rect 31297 28027 31355 28033
rect 31726 28008 31754 28036
rect 32309 28033 32321 28067
rect 32355 28064 32367 28067
rect 32398 28064 32404 28076
rect 32355 28036 32404 28064
rect 32355 28033 32367 28036
rect 32309 28027 32367 28033
rect 32398 28024 32404 28036
rect 32456 28024 32462 28076
rect 32582 28024 32588 28076
rect 32640 28064 32646 28076
rect 32677 28067 32735 28073
rect 32677 28064 32689 28067
rect 32640 28036 32689 28064
rect 32640 28024 32646 28036
rect 32677 28033 32689 28036
rect 32723 28033 32735 28067
rect 32677 28027 32735 28033
rect 30190 27996 30196 28008
rect 29288 27968 30196 27996
rect 30190 27956 30196 27968
rect 30248 27956 30254 28008
rect 30558 27956 30564 28008
rect 30616 27996 30622 28008
rect 30616 27968 31156 27996
rect 30616 27956 30622 27968
rect 25866 27928 25872 27940
rect 25516 27900 25872 27928
rect 25866 27888 25872 27900
rect 25924 27888 25930 27940
rect 19208 27832 20208 27860
rect 20441 27863 20499 27869
rect 19208 27820 19214 27832
rect 20441 27829 20453 27863
rect 20487 27860 20499 27863
rect 20530 27860 20536 27872
rect 20487 27832 20536 27860
rect 20487 27829 20499 27832
rect 20441 27823 20499 27829
rect 20530 27820 20536 27832
rect 20588 27820 20594 27872
rect 23017 27863 23075 27869
rect 23017 27829 23029 27863
rect 23063 27860 23075 27863
rect 23290 27860 23296 27872
rect 23063 27832 23296 27860
rect 23063 27829 23075 27832
rect 23017 27823 23075 27829
rect 23290 27820 23296 27832
rect 23348 27820 23354 27872
rect 24210 27820 24216 27872
rect 24268 27860 24274 27872
rect 25130 27860 25136 27872
rect 24268 27832 25136 27860
rect 24268 27820 24274 27832
rect 25130 27820 25136 27832
rect 25188 27860 25194 27872
rect 29914 27860 29920 27872
rect 25188 27832 29920 27860
rect 25188 27820 25194 27832
rect 29914 27820 29920 27832
rect 29972 27820 29978 27872
rect 30098 27820 30104 27872
rect 30156 27860 30162 27872
rect 30282 27860 30288 27872
rect 30156 27832 30288 27860
rect 30156 27820 30162 27832
rect 30282 27820 30288 27832
rect 30340 27860 30346 27872
rect 30650 27869 30656 27872
rect 30607 27863 30656 27869
rect 30607 27860 30619 27863
rect 30340 27832 30619 27860
rect 30340 27820 30346 27832
rect 30607 27829 30619 27832
rect 30653 27829 30656 27863
rect 30607 27823 30656 27829
rect 30650 27820 30656 27823
rect 30708 27820 30714 27872
rect 31128 27869 31156 27968
rect 31662 27956 31668 28008
rect 31720 27996 31754 28008
rect 32766 27996 32772 28008
rect 31720 27968 32772 27996
rect 31720 27956 31726 27968
rect 32766 27956 32772 27968
rect 32824 27956 32830 28008
rect 31478 27888 31484 27940
rect 31536 27928 31542 27940
rect 31938 27928 31944 27940
rect 31536 27900 31944 27928
rect 31536 27888 31542 27900
rect 31938 27888 31944 27900
rect 31996 27888 32002 27940
rect 36998 27928 37004 27940
rect 32048 27900 37004 27928
rect 31113 27863 31171 27869
rect 31113 27829 31125 27863
rect 31159 27860 31171 27863
rect 32048 27860 32076 27900
rect 36998 27888 37004 27900
rect 37056 27888 37062 27940
rect 31159 27832 32076 27860
rect 31159 27829 31171 27832
rect 31113 27823 31171 27829
rect 32122 27820 32128 27872
rect 32180 27860 32186 27872
rect 32769 27863 32827 27869
rect 32769 27860 32781 27863
rect 32180 27832 32781 27860
rect 32180 27820 32186 27832
rect 32769 27829 32781 27832
rect 32815 27829 32827 27863
rect 32769 27823 32827 27829
rect 1104 27770 40572 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 40572 27770
rect 1104 27696 40572 27718
rect 7272 27659 7330 27665
rect 7272 27625 7284 27659
rect 7318 27656 7330 27659
rect 8386 27656 8392 27668
rect 7318 27628 8392 27656
rect 7318 27625 7330 27628
rect 7272 27619 7330 27625
rect 8386 27616 8392 27628
rect 8444 27616 8450 27668
rect 11333 27659 11391 27665
rect 11333 27625 11345 27659
rect 11379 27656 11391 27659
rect 11514 27656 11520 27668
rect 11379 27628 11520 27656
rect 11379 27625 11391 27628
rect 11333 27619 11391 27625
rect 5534 27548 5540 27600
rect 5592 27588 5598 27600
rect 6454 27588 6460 27600
rect 5592 27560 6460 27588
rect 5592 27548 5598 27560
rect 6454 27548 6460 27560
rect 6512 27548 6518 27600
rect 3786 27480 3792 27532
rect 3844 27480 3850 27532
rect 6822 27480 6828 27532
rect 6880 27520 6886 27532
rect 7009 27523 7067 27529
rect 7009 27520 7021 27523
rect 6880 27492 7021 27520
rect 6880 27480 6886 27492
rect 7009 27489 7021 27492
rect 7055 27489 7067 27523
rect 7009 27483 7067 27489
rect 8757 27523 8815 27529
rect 8757 27489 8769 27523
rect 8803 27489 8815 27523
rect 8757 27483 8815 27489
rect 8772 27452 8800 27483
rect 9582 27480 9588 27532
rect 9640 27480 9646 27532
rect 9677 27523 9735 27529
rect 9677 27489 9689 27523
rect 9723 27520 9735 27523
rect 11348 27520 11376 27619
rect 11514 27616 11520 27628
rect 11572 27656 11578 27668
rect 11790 27656 11796 27668
rect 11572 27628 11796 27656
rect 11572 27616 11578 27628
rect 11790 27616 11796 27628
rect 11848 27616 11854 27668
rect 12710 27616 12716 27668
rect 12768 27656 12774 27668
rect 12768 27628 13584 27656
rect 12768 27616 12774 27628
rect 13556 27600 13584 27628
rect 13814 27616 13820 27668
rect 13872 27656 13878 27668
rect 14550 27656 14556 27668
rect 13872 27628 14556 27656
rect 13872 27616 13878 27628
rect 14550 27616 14556 27628
rect 14608 27616 14614 27668
rect 14734 27616 14740 27668
rect 14792 27656 14798 27668
rect 15746 27656 15752 27668
rect 14792 27628 15752 27656
rect 14792 27616 14798 27628
rect 15746 27616 15752 27628
rect 15804 27616 15810 27668
rect 17678 27616 17684 27668
rect 17736 27616 17742 27668
rect 17862 27616 17868 27668
rect 17920 27616 17926 27668
rect 18432 27628 28994 27656
rect 12986 27548 12992 27600
rect 13044 27548 13050 27600
rect 13538 27548 13544 27600
rect 13596 27588 13602 27600
rect 15194 27588 15200 27600
rect 13596 27560 15200 27588
rect 13596 27548 13602 27560
rect 9723 27492 11376 27520
rect 9723 27489 9735 27492
rect 9677 27483 9735 27489
rect 12250 27480 12256 27532
rect 12308 27520 12314 27532
rect 12437 27523 12495 27529
rect 12437 27520 12449 27523
rect 12308 27492 12449 27520
rect 12308 27480 12314 27492
rect 12437 27489 12449 27492
rect 12483 27489 12495 27523
rect 12437 27483 12495 27489
rect 9858 27452 9864 27464
rect 8772 27424 9864 27452
rect 9858 27412 9864 27424
rect 9916 27452 9922 27464
rect 10686 27452 10692 27464
rect 9916 27424 10692 27452
rect 9916 27412 9922 27424
rect 10686 27412 10692 27424
rect 10744 27412 10750 27464
rect 10870 27412 10876 27464
rect 10928 27452 10934 27464
rect 11057 27455 11115 27461
rect 11057 27452 11069 27455
rect 10928 27424 11069 27452
rect 10928 27412 10934 27424
rect 11057 27421 11069 27424
rect 11103 27421 11115 27455
rect 11057 27415 11115 27421
rect 11146 27412 11152 27464
rect 11204 27452 11210 27464
rect 12268 27452 12296 27480
rect 11204 27424 12296 27452
rect 12529 27455 12587 27461
rect 11204 27412 11210 27424
rect 12529 27421 12541 27455
rect 12575 27452 12587 27455
rect 13004 27452 13032 27548
rect 13173 27523 13231 27529
rect 13173 27489 13185 27523
rect 13219 27520 13231 27523
rect 13817 27523 13875 27529
rect 13817 27520 13829 27523
rect 13219 27492 13829 27520
rect 13219 27489 13231 27492
rect 13173 27483 13231 27489
rect 13817 27489 13829 27492
rect 13863 27489 13875 27523
rect 13817 27483 13875 27489
rect 12575 27424 13032 27452
rect 12575 27421 12587 27424
rect 12529 27415 12587 27421
rect 13262 27412 13268 27464
rect 13320 27412 13326 27464
rect 13357 27455 13415 27461
rect 13357 27421 13369 27455
rect 13403 27421 13415 27455
rect 13357 27415 13415 27421
rect 4062 27344 4068 27396
rect 4120 27344 4126 27396
rect 7742 27384 7748 27396
rect 5290 27356 7748 27384
rect 7742 27344 7748 27356
rect 7800 27344 7806 27396
rect 9766 27344 9772 27396
rect 9824 27384 9830 27396
rect 13372 27384 13400 27415
rect 13446 27412 13452 27464
rect 13504 27412 13510 27464
rect 14292 27461 14320 27560
rect 15194 27548 15200 27560
rect 15252 27588 15258 27600
rect 16666 27588 16672 27600
rect 15252 27560 16672 27588
rect 15252 27548 15258 27560
rect 16666 27548 16672 27560
rect 16724 27588 16730 27600
rect 18325 27591 18383 27597
rect 18325 27588 18337 27591
rect 16724 27560 18337 27588
rect 16724 27548 16730 27560
rect 18325 27557 18337 27560
rect 18371 27557 18383 27591
rect 18325 27551 18383 27557
rect 15010 27520 15016 27532
rect 14384 27492 15016 27520
rect 14384 27461 14412 27492
rect 15010 27480 15016 27492
rect 15068 27480 15074 27532
rect 13725 27455 13783 27461
rect 13725 27421 13737 27455
rect 13771 27421 13783 27455
rect 13725 27415 13783 27421
rect 13909 27455 13967 27461
rect 13909 27421 13921 27455
rect 13955 27452 13967 27455
rect 14277 27455 14335 27461
rect 13955 27424 14228 27452
rect 13955 27421 13967 27424
rect 13909 27415 13967 27421
rect 9824 27356 13400 27384
rect 13740 27384 13768 27415
rect 14090 27384 14096 27396
rect 13740 27356 14096 27384
rect 9824 27344 9830 27356
rect 14090 27344 14096 27356
rect 14148 27344 14154 27396
rect 4338 27276 4344 27328
rect 4396 27316 4402 27328
rect 9107 27319 9165 27325
rect 9107 27316 9119 27319
rect 4396 27288 9119 27316
rect 4396 27276 4402 27288
rect 9107 27285 9119 27288
rect 9153 27285 9165 27319
rect 9107 27279 9165 27285
rect 9585 27319 9643 27325
rect 9585 27285 9597 27319
rect 9631 27316 9643 27319
rect 11146 27316 11152 27328
rect 9631 27288 11152 27316
rect 9631 27285 9643 27288
rect 9585 27279 9643 27285
rect 11146 27276 11152 27288
rect 11204 27276 11210 27328
rect 14200 27316 14228 27424
rect 14277 27421 14289 27455
rect 14323 27421 14335 27455
rect 14277 27415 14335 27421
rect 14369 27455 14427 27461
rect 14369 27421 14381 27455
rect 14415 27421 14427 27455
rect 14369 27415 14427 27421
rect 14550 27412 14556 27464
rect 14608 27412 14614 27464
rect 14642 27412 14648 27464
rect 14700 27412 14706 27464
rect 14734 27412 14740 27464
rect 14792 27412 14798 27464
rect 15212 27461 15240 27548
rect 15838 27520 15844 27532
rect 15580 27492 15844 27520
rect 15197 27455 15255 27461
rect 15197 27421 15209 27455
rect 15243 27421 15255 27455
rect 15197 27415 15255 27421
rect 15290 27455 15348 27461
rect 15290 27421 15302 27455
rect 15336 27421 15348 27455
rect 15290 27415 15348 27421
rect 14826 27344 14832 27396
rect 14884 27384 14890 27396
rect 15305 27384 15333 27415
rect 15470 27412 15476 27464
rect 15528 27412 15534 27464
rect 15580 27461 15608 27492
rect 15838 27480 15844 27492
rect 15896 27480 15902 27532
rect 15930 27480 15936 27532
rect 15988 27520 15994 27532
rect 18432 27520 18460 27628
rect 19886 27548 19892 27600
rect 19944 27588 19950 27600
rect 20898 27588 20904 27600
rect 19944 27560 20904 27588
rect 19944 27548 19950 27560
rect 20898 27548 20904 27560
rect 20956 27548 20962 27600
rect 24486 27548 24492 27600
rect 24544 27588 24550 27600
rect 28966 27588 28994 27628
rect 30374 27616 30380 27668
rect 30432 27656 30438 27668
rect 31202 27656 31208 27668
rect 30432 27628 31208 27656
rect 30432 27616 30438 27628
rect 31202 27616 31208 27628
rect 31260 27616 31266 27668
rect 36078 27616 36084 27668
rect 36136 27656 36142 27668
rect 36633 27659 36691 27665
rect 36633 27656 36645 27659
rect 36136 27628 36645 27656
rect 36136 27616 36142 27628
rect 36633 27625 36645 27628
rect 36679 27625 36691 27659
rect 36633 27619 36691 27625
rect 37090 27616 37096 27668
rect 37148 27656 37154 27668
rect 37277 27659 37335 27665
rect 37277 27656 37289 27659
rect 37148 27628 37289 27656
rect 37148 27616 37154 27628
rect 37277 27625 37289 27628
rect 37323 27625 37335 27659
rect 37277 27619 37335 27625
rect 30742 27588 30748 27600
rect 24544 27560 28304 27588
rect 28966 27560 30748 27588
rect 24544 27548 24550 27560
rect 20806 27520 20812 27532
rect 15988 27492 18460 27520
rect 18615 27492 18920 27520
rect 15988 27480 15994 27492
rect 15746 27461 15752 27464
rect 15565 27455 15623 27461
rect 15565 27421 15577 27455
rect 15611 27421 15623 27455
rect 15565 27415 15623 27421
rect 15703 27455 15752 27461
rect 15703 27421 15715 27455
rect 15749 27421 15752 27455
rect 15703 27415 15752 27421
rect 15746 27412 15752 27415
rect 15804 27412 15810 27464
rect 17313 27455 17371 27461
rect 17313 27421 17325 27455
rect 17359 27452 17371 27455
rect 17402 27452 17408 27464
rect 17359 27424 17408 27452
rect 17359 27421 17371 27424
rect 17313 27415 17371 27421
rect 17402 27412 17408 27424
rect 17460 27412 17466 27464
rect 17497 27455 17555 27461
rect 17497 27421 17509 27455
rect 17543 27452 17555 27455
rect 18506 27452 18512 27464
rect 17543 27424 18512 27452
rect 17543 27421 17555 27424
rect 17497 27415 17555 27421
rect 18506 27412 18512 27424
rect 18564 27412 18570 27464
rect 18615 27439 18643 27492
rect 18600 27433 18658 27439
rect 18600 27399 18612 27433
rect 18646 27399 18658 27433
rect 18690 27412 18696 27464
rect 18748 27412 18754 27464
rect 18782 27412 18788 27464
rect 18840 27412 18846 27464
rect 14884 27356 15333 27384
rect 14884 27344 14890 27356
rect 17770 27344 17776 27396
rect 17828 27393 17834 27396
rect 17828 27387 17877 27393
rect 17828 27353 17831 27387
rect 17865 27353 17877 27387
rect 17828 27347 17877 27353
rect 17828 27344 17834 27347
rect 18230 27344 18236 27396
rect 18288 27344 18294 27396
rect 18600 27393 18658 27399
rect 18892 27384 18920 27492
rect 19306 27492 20812 27520
rect 18966 27412 18972 27464
rect 19024 27452 19030 27464
rect 19306 27452 19334 27492
rect 20806 27480 20812 27492
rect 20864 27480 20870 27532
rect 22830 27480 22836 27532
rect 22888 27520 22894 27532
rect 23198 27520 23204 27532
rect 22888 27492 23204 27520
rect 22888 27480 22894 27492
rect 23198 27480 23204 27492
rect 23256 27480 23262 27532
rect 27890 27520 27896 27532
rect 25424 27492 27896 27520
rect 19024 27424 19334 27452
rect 19521 27455 19579 27461
rect 19024 27412 19030 27424
rect 19521 27421 19533 27455
rect 19567 27452 19579 27455
rect 19610 27452 19616 27464
rect 19567 27424 19616 27452
rect 19567 27421 19579 27424
rect 19521 27415 19579 27421
rect 19610 27412 19616 27424
rect 19668 27412 19674 27464
rect 19702 27412 19708 27464
rect 19760 27452 19766 27464
rect 20346 27452 20352 27464
rect 19760 27424 20352 27452
rect 19760 27412 19766 27424
rect 20346 27412 20352 27424
rect 20404 27452 20410 27464
rect 20441 27455 20499 27461
rect 20441 27452 20453 27455
rect 20404 27424 20453 27452
rect 20404 27412 20410 27424
rect 20441 27421 20453 27424
rect 20487 27421 20499 27455
rect 20441 27415 20499 27421
rect 20622 27412 20628 27464
rect 20680 27412 20686 27464
rect 25424 27461 25452 27492
rect 27890 27480 27896 27492
rect 27948 27520 27954 27532
rect 28166 27520 28172 27532
rect 27948 27492 28172 27520
rect 27948 27480 27954 27492
rect 28166 27480 28172 27492
rect 28224 27480 28230 27532
rect 25409 27455 25467 27461
rect 25409 27421 25421 27455
rect 25455 27421 25467 27455
rect 25409 27415 25467 27421
rect 25501 27455 25559 27461
rect 25501 27421 25513 27455
rect 25547 27452 25559 27455
rect 26510 27452 26516 27464
rect 25547 27424 26516 27452
rect 25547 27421 25559 27424
rect 25501 27415 25559 27421
rect 19426 27384 19432 27396
rect 18892 27356 19432 27384
rect 19426 27344 19432 27356
rect 19484 27344 19490 27396
rect 19628 27356 19840 27384
rect 14366 27316 14372 27328
rect 14200 27288 14372 27316
rect 14366 27276 14372 27288
rect 14424 27276 14430 27328
rect 14461 27319 14519 27325
rect 14461 27285 14473 27319
rect 14507 27316 14519 27319
rect 14918 27316 14924 27328
rect 14507 27288 14924 27316
rect 14507 27285 14519 27288
rect 14461 27279 14519 27285
rect 14918 27276 14924 27288
rect 14976 27276 14982 27328
rect 15841 27319 15899 27325
rect 15841 27285 15853 27319
rect 15887 27316 15899 27319
rect 16022 27316 16028 27328
rect 15887 27288 16028 27316
rect 15887 27285 15899 27288
rect 15841 27279 15899 27285
rect 16022 27276 16028 27288
rect 16080 27276 16086 27328
rect 16206 27276 16212 27328
rect 16264 27316 16270 27328
rect 17221 27319 17279 27325
rect 17221 27316 17233 27319
rect 16264 27288 17233 27316
rect 16264 27276 16270 27288
rect 17221 27285 17233 27288
rect 17267 27285 17279 27319
rect 17221 27279 17279 27285
rect 18046 27276 18052 27328
rect 18104 27316 18110 27328
rect 19628 27325 19656 27356
rect 19337 27319 19395 27325
rect 19337 27316 19349 27319
rect 18104 27288 19349 27316
rect 18104 27276 18110 27288
rect 19337 27285 19349 27288
rect 19383 27285 19395 27319
rect 19337 27279 19395 27285
rect 19613 27319 19671 27325
rect 19613 27285 19625 27319
rect 19659 27285 19671 27319
rect 19613 27279 19671 27285
rect 19702 27276 19708 27328
rect 19760 27276 19766 27328
rect 19812 27316 19840 27356
rect 19886 27344 19892 27396
rect 19944 27344 19950 27396
rect 24854 27344 24860 27396
rect 24912 27384 24918 27396
rect 25516 27384 25544 27415
rect 26510 27412 26516 27424
rect 26568 27452 26574 27464
rect 27338 27452 27344 27464
rect 26568 27424 27344 27452
rect 26568 27412 26574 27424
rect 27338 27412 27344 27424
rect 27396 27412 27402 27464
rect 27706 27412 27712 27464
rect 27764 27452 27770 27464
rect 28074 27452 28080 27464
rect 27764 27424 28080 27452
rect 27764 27412 27770 27424
rect 28074 27412 28080 27424
rect 28132 27412 28138 27464
rect 28276 27452 28304 27560
rect 30742 27548 30748 27560
rect 30800 27548 30806 27600
rect 30926 27548 30932 27600
rect 30984 27548 30990 27600
rect 31846 27588 31852 27600
rect 31726 27560 31852 27588
rect 29730 27480 29736 27532
rect 29788 27480 29794 27532
rect 30558 27480 30564 27532
rect 30616 27480 30622 27532
rect 31018 27480 31024 27532
rect 31076 27480 31082 27532
rect 28718 27452 28724 27464
rect 28276 27424 28724 27452
rect 28718 27412 28724 27424
rect 28776 27452 28782 27464
rect 29638 27452 29644 27464
rect 28776 27424 29644 27452
rect 28776 27412 28782 27424
rect 29638 27412 29644 27424
rect 29696 27452 29702 27464
rect 29917 27455 29975 27461
rect 29917 27452 29929 27455
rect 29696 27424 29929 27452
rect 29696 27412 29702 27424
rect 29917 27421 29929 27424
rect 29963 27421 29975 27455
rect 29917 27415 29975 27421
rect 30745 27455 30803 27461
rect 30745 27421 30757 27455
rect 30791 27452 30803 27455
rect 31726 27452 31754 27560
rect 31846 27548 31852 27560
rect 31904 27588 31910 27600
rect 32306 27588 32312 27600
rect 31904 27560 32312 27588
rect 31904 27548 31910 27560
rect 32306 27548 32312 27560
rect 32364 27548 32370 27600
rect 32582 27548 32588 27600
rect 32640 27588 32646 27600
rect 33505 27591 33563 27597
rect 32640 27560 33364 27588
rect 32640 27548 32646 27560
rect 32122 27480 32128 27532
rect 32180 27480 32186 27532
rect 32950 27520 32956 27532
rect 32298 27492 32956 27520
rect 32298 27461 32326 27492
rect 32950 27480 32956 27492
rect 33008 27480 33014 27532
rect 33336 27529 33364 27560
rect 33505 27557 33517 27591
rect 33551 27588 33563 27591
rect 38654 27588 38660 27600
rect 33551 27560 38660 27588
rect 33551 27557 33563 27560
rect 33505 27551 33563 27557
rect 38654 27548 38660 27560
rect 38712 27548 38718 27600
rect 33320 27523 33378 27529
rect 33320 27489 33332 27523
rect 33366 27489 33378 27523
rect 33320 27483 33378 27489
rect 34422 27480 34428 27532
rect 34480 27520 34486 27532
rect 37093 27523 37151 27529
rect 34480 27492 36768 27520
rect 34480 27480 34486 27492
rect 30791 27424 31754 27452
rect 32283 27455 32341 27461
rect 30791 27421 30803 27424
rect 30745 27415 30803 27421
rect 32283 27421 32295 27455
rect 32329 27421 32341 27455
rect 32283 27415 32341 27421
rect 32582 27412 32588 27464
rect 32640 27412 32646 27464
rect 32766 27412 32772 27464
rect 32824 27452 32830 27464
rect 33045 27455 33103 27461
rect 33045 27452 33057 27455
rect 32824 27424 33057 27452
rect 32824 27412 32830 27424
rect 33045 27421 33057 27424
rect 33091 27421 33103 27455
rect 33045 27415 33103 27421
rect 33134 27412 33140 27464
rect 33192 27412 33198 27464
rect 33229 27455 33287 27461
rect 33229 27421 33241 27455
rect 33275 27452 33287 27455
rect 33778 27452 33784 27464
rect 33275 27424 33784 27452
rect 33275 27421 33287 27424
rect 33229 27415 33287 27421
rect 24912 27356 25544 27384
rect 24912 27344 24918 27356
rect 25590 27344 25596 27396
rect 25648 27384 25654 27396
rect 25685 27387 25743 27393
rect 25685 27384 25697 27387
rect 25648 27356 25697 27384
rect 25648 27344 25654 27356
rect 25685 27353 25697 27356
rect 25731 27353 25743 27387
rect 25685 27347 25743 27353
rect 25774 27344 25780 27396
rect 25832 27384 25838 27396
rect 25832 27356 31156 27384
rect 25832 27344 25838 27356
rect 20254 27316 20260 27328
rect 19812 27288 20260 27316
rect 20254 27276 20260 27288
rect 20312 27276 20318 27328
rect 24302 27276 24308 27328
rect 24360 27316 24366 27328
rect 24578 27316 24584 27328
rect 24360 27288 24584 27316
rect 24360 27276 24366 27288
rect 24578 27276 24584 27288
rect 24636 27316 24642 27328
rect 25409 27319 25467 27325
rect 25409 27316 25421 27319
rect 24636 27288 25421 27316
rect 24636 27276 24642 27288
rect 25409 27285 25421 27288
rect 25455 27285 25467 27319
rect 31128 27316 31156 27356
rect 31202 27344 31208 27396
rect 31260 27344 31266 27396
rect 31386 27344 31392 27396
rect 31444 27384 31450 27396
rect 32122 27384 32128 27396
rect 31444 27356 32128 27384
rect 31444 27344 31450 27356
rect 32122 27344 32128 27356
rect 32180 27344 32186 27396
rect 32398 27344 32404 27396
rect 32456 27344 32462 27396
rect 32493 27387 32551 27393
rect 32493 27353 32505 27387
rect 32539 27384 32551 27387
rect 33244 27384 33272 27415
rect 33778 27412 33784 27424
rect 33836 27412 33842 27464
rect 36633 27455 36691 27461
rect 36633 27421 36645 27455
rect 36679 27421 36691 27455
rect 36633 27415 36691 27421
rect 36648 27384 36676 27415
rect 32539 27356 33272 27384
rect 36556 27356 36676 27384
rect 36740 27384 36768 27492
rect 37093 27489 37105 27523
rect 37139 27520 37151 27523
rect 37182 27520 37188 27532
rect 37139 27492 37188 27520
rect 37139 27489 37151 27492
rect 37093 27483 37151 27489
rect 37182 27480 37188 27492
rect 37240 27480 37246 27532
rect 38102 27480 38108 27532
rect 38160 27520 38166 27532
rect 39301 27523 39359 27529
rect 39301 27520 39313 27523
rect 38160 27492 39313 27520
rect 38160 27480 38166 27492
rect 39301 27489 39313 27492
rect 39347 27489 39359 27523
rect 39301 27483 39359 27489
rect 36814 27412 36820 27464
rect 36872 27412 36878 27464
rect 37366 27412 37372 27464
rect 37424 27452 37430 27464
rect 38010 27452 38016 27464
rect 37424 27424 38016 27452
rect 37424 27412 37430 27424
rect 38010 27412 38016 27424
rect 38068 27412 38074 27464
rect 38838 27384 38844 27396
rect 36740 27356 38844 27384
rect 32539 27353 32551 27356
rect 32493 27347 32551 27353
rect 32508 27316 32536 27347
rect 36556 27328 36584 27356
rect 38838 27344 38844 27356
rect 38896 27344 38902 27396
rect 39574 27344 39580 27396
rect 39632 27344 39638 27396
rect 31128 27288 32536 27316
rect 25409 27279 25467 27285
rect 32766 27276 32772 27328
rect 32824 27276 32830 27328
rect 32950 27276 32956 27328
rect 33008 27316 33014 27328
rect 35986 27316 35992 27328
rect 33008 27288 35992 27316
rect 33008 27276 33014 27288
rect 35986 27276 35992 27288
rect 36044 27276 36050 27328
rect 36538 27276 36544 27328
rect 36596 27276 36602 27328
rect 36906 27276 36912 27328
rect 36964 27316 36970 27328
rect 37001 27319 37059 27325
rect 37001 27316 37013 27319
rect 36964 27288 37013 27316
rect 36964 27276 36970 27288
rect 37001 27285 37013 27288
rect 37047 27285 37059 27319
rect 37001 27279 37059 27285
rect 37093 27319 37151 27325
rect 37093 27285 37105 27319
rect 37139 27316 37151 27319
rect 37458 27316 37464 27328
rect 37139 27288 37464 27316
rect 37139 27285 37151 27288
rect 37093 27279 37151 27285
rect 37458 27276 37464 27288
rect 37516 27276 37522 27328
rect 1104 27226 40572 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 40572 27226
rect 1104 27152 40572 27174
rect 3973 27115 4031 27121
rect 3973 27081 3985 27115
rect 4019 27112 4031 27115
rect 4062 27112 4068 27124
rect 4019 27084 4068 27112
rect 4019 27081 4031 27084
rect 3973 27075 4031 27081
rect 4062 27072 4068 27084
rect 4120 27072 4126 27124
rect 4338 27072 4344 27124
rect 4396 27072 4402 27124
rect 4433 27115 4491 27121
rect 4433 27081 4445 27115
rect 4479 27112 4491 27115
rect 5534 27112 5540 27124
rect 4479 27084 5540 27112
rect 4479 27081 4491 27084
rect 4433 27075 4491 27081
rect 5534 27072 5540 27084
rect 5592 27072 5598 27124
rect 5902 27072 5908 27124
rect 5960 27112 5966 27124
rect 6730 27112 6736 27124
rect 5960 27084 6736 27112
rect 5960 27072 5966 27084
rect 6730 27072 6736 27084
rect 6788 27072 6794 27124
rect 8386 27072 8392 27124
rect 8444 27072 8450 27124
rect 8757 27115 8815 27121
rect 8757 27081 8769 27115
rect 8803 27112 8815 27115
rect 9674 27112 9680 27124
rect 8803 27084 9680 27112
rect 8803 27081 8815 27084
rect 8757 27075 8815 27081
rect 9674 27072 9680 27084
rect 9732 27072 9738 27124
rect 9766 27072 9772 27124
rect 9824 27072 9830 27124
rect 10226 27072 10232 27124
rect 10284 27072 10290 27124
rect 11054 27112 11060 27124
rect 10428 27084 11060 27112
rect 3142 27004 3148 27056
rect 3200 27044 3206 27056
rect 4356 27044 4384 27072
rect 3200 27016 4384 27044
rect 3200 27004 3206 27016
rect 6086 27004 6092 27056
rect 6144 27044 6150 27056
rect 6457 27047 6515 27053
rect 6457 27044 6469 27047
rect 6144 27016 6469 27044
rect 6144 27004 6150 27016
rect 6457 27013 6469 27016
rect 6503 27013 6515 27047
rect 6457 27007 6515 27013
rect 6641 27047 6699 27053
rect 6641 27013 6653 27047
rect 6687 27044 6699 27047
rect 7282 27044 7288 27056
rect 6687 27016 7288 27044
rect 6687 27013 6699 27016
rect 6641 27007 6699 27013
rect 7282 27004 7288 27016
rect 7340 27004 7346 27056
rect 7926 27004 7932 27056
rect 7984 27044 7990 27056
rect 10428 27044 10456 27084
rect 11054 27072 11060 27084
rect 11112 27072 11118 27124
rect 11149 27115 11207 27121
rect 11149 27081 11161 27115
rect 11195 27112 11207 27115
rect 11238 27112 11244 27124
rect 11195 27084 11244 27112
rect 11195 27081 11207 27084
rect 11149 27075 11207 27081
rect 11238 27072 11244 27084
rect 11296 27072 11302 27124
rect 11701 27115 11759 27121
rect 11701 27081 11713 27115
rect 11747 27081 11759 27115
rect 11701 27075 11759 27081
rect 13541 27115 13599 27121
rect 13541 27081 13553 27115
rect 13587 27112 13599 27115
rect 13722 27112 13728 27124
rect 13587 27084 13728 27112
rect 13587 27081 13599 27084
rect 13541 27075 13599 27081
rect 7984 27016 9720 27044
rect 7984 27004 7990 27016
rect 5629 26979 5687 26985
rect 5629 26945 5641 26979
rect 5675 26976 5687 26979
rect 5675 26948 5764 26976
rect 5675 26945 5687 26948
rect 5629 26939 5687 26945
rect 4614 26868 4620 26920
rect 4672 26868 4678 26920
rect 5736 26840 5764 26948
rect 5810 26936 5816 26988
rect 5868 26936 5874 26988
rect 5902 26936 5908 26988
rect 5960 26936 5966 26988
rect 5997 26979 6055 26985
rect 5997 26945 6009 26979
rect 6043 26976 6055 26979
rect 6362 26976 6368 26988
rect 6043 26948 6368 26976
rect 6043 26945 6055 26948
rect 5997 26939 6055 26945
rect 6362 26936 6368 26948
rect 6420 26936 6426 26988
rect 6822 26936 6828 26988
rect 6880 26936 6886 26988
rect 9692 26985 9720 27016
rect 9876 27016 10456 27044
rect 9876 26985 9904 27016
rect 8849 26979 8907 26985
rect 8849 26945 8861 26979
rect 8895 26976 8907 26979
rect 9677 26979 9735 26985
rect 8895 26948 9628 26976
rect 8895 26945 8907 26948
rect 8849 26939 8907 26945
rect 8478 26868 8484 26920
rect 8536 26908 8542 26920
rect 8754 26908 8760 26920
rect 8536 26880 8760 26908
rect 8536 26868 8542 26880
rect 8754 26868 8760 26880
rect 8812 26908 8818 26920
rect 8941 26911 8999 26917
rect 8941 26908 8953 26911
rect 8812 26880 8953 26908
rect 8812 26868 8818 26880
rect 8941 26877 8953 26880
rect 8987 26877 8999 26911
rect 9600 26908 9628 26948
rect 9677 26945 9689 26979
rect 9723 26945 9735 26979
rect 9677 26939 9735 26945
rect 9861 26979 9919 26985
rect 9861 26945 9873 26979
rect 9907 26945 9919 26979
rect 9861 26939 9919 26945
rect 10137 26979 10195 26985
rect 10137 26945 10149 26979
rect 10183 26976 10195 26979
rect 10226 26976 10232 26988
rect 10183 26948 10232 26976
rect 10183 26945 10195 26948
rect 10137 26939 10195 26945
rect 10226 26936 10232 26948
rect 10284 26936 10290 26988
rect 10428 26985 10456 27016
rect 10686 27004 10692 27056
rect 10744 27004 10750 27056
rect 10962 27004 10968 27056
rect 11020 27044 11026 27056
rect 11716 27044 11744 27075
rect 13722 27072 13728 27084
rect 13780 27072 13786 27124
rect 14642 27072 14648 27124
rect 14700 27112 14706 27124
rect 15102 27112 15108 27124
rect 14700 27084 15108 27112
rect 14700 27072 14706 27084
rect 15102 27072 15108 27084
rect 15160 27072 15166 27124
rect 15286 27072 15292 27124
rect 15344 27112 15350 27124
rect 15838 27112 15844 27124
rect 15344 27084 15844 27112
rect 15344 27072 15350 27084
rect 15838 27072 15844 27084
rect 15896 27072 15902 27124
rect 16482 27072 16488 27124
rect 16540 27112 16546 27124
rect 16669 27115 16727 27121
rect 16669 27112 16681 27115
rect 16540 27084 16681 27112
rect 16540 27072 16546 27084
rect 16669 27081 16681 27084
rect 16715 27081 16727 27115
rect 16669 27075 16727 27081
rect 18432 27084 19564 27112
rect 11020 27016 11744 27044
rect 11020 27004 11026 27016
rect 12434 27004 12440 27056
rect 12492 27044 12498 27056
rect 17497 27047 17555 27053
rect 17497 27044 17509 27047
rect 12492 27016 17509 27044
rect 12492 27004 12498 27016
rect 17497 27013 17509 27016
rect 17543 27013 17555 27047
rect 18432 27044 18460 27084
rect 17497 27007 17555 27013
rect 17788 27016 18460 27044
rect 17788 26988 17816 27016
rect 10321 26979 10379 26985
rect 10321 26945 10333 26979
rect 10367 26945 10379 26979
rect 10321 26939 10379 26945
rect 10413 26979 10471 26985
rect 10413 26945 10425 26979
rect 10459 26945 10471 26979
rect 10413 26939 10471 26945
rect 9766 26908 9772 26920
rect 9600 26880 9772 26908
rect 8941 26871 8999 26877
rect 9766 26868 9772 26880
rect 9824 26868 9830 26920
rect 6270 26840 6276 26852
rect 5736 26812 6276 26840
rect 6270 26800 6276 26812
rect 6328 26840 6334 26852
rect 9490 26840 9496 26852
rect 6328 26812 9496 26840
rect 6328 26800 6334 26812
rect 9490 26800 9496 26812
rect 9548 26800 9554 26852
rect 9784 26840 9812 26868
rect 10134 26840 10140 26852
rect 9784 26812 10140 26840
rect 10134 26800 10140 26812
rect 10192 26800 10198 26852
rect 10336 26840 10364 26939
rect 10502 26936 10508 26988
rect 10560 26936 10566 26988
rect 10781 26979 10839 26985
rect 10781 26976 10793 26979
rect 10612 26948 10793 26976
rect 10612 26920 10640 26948
rect 10781 26945 10793 26948
rect 10827 26945 10839 26979
rect 10781 26939 10839 26945
rect 11514 26936 11520 26988
rect 11572 26936 11578 26988
rect 13354 26936 13360 26988
rect 13412 26936 13418 26988
rect 13633 26979 13691 26985
rect 13633 26945 13645 26979
rect 13679 26976 13691 26979
rect 13814 26976 13820 26988
rect 13679 26948 13820 26976
rect 13679 26945 13691 26948
rect 13633 26939 13691 26945
rect 13814 26936 13820 26948
rect 13872 26976 13878 26988
rect 14550 26976 14556 26988
rect 13872 26948 14556 26976
rect 13872 26936 13878 26948
rect 14550 26936 14556 26948
rect 14608 26936 14614 26988
rect 14918 26936 14924 26988
rect 14976 26936 14982 26988
rect 15286 26936 15292 26988
rect 15344 26936 15350 26988
rect 15473 26979 15531 26985
rect 15473 26945 15485 26979
rect 15519 26976 15531 26979
rect 16206 26976 16212 26988
rect 15519 26948 16212 26976
rect 15519 26945 15531 26948
rect 15473 26939 15531 26945
rect 10594 26908 10600 26920
rect 10652 26917 10658 26920
rect 10652 26911 10674 26917
rect 10526 26880 10600 26908
rect 10594 26868 10600 26880
rect 10662 26877 10674 26911
rect 10652 26871 10674 26877
rect 10873 26911 10931 26917
rect 10873 26877 10885 26911
rect 10919 26908 10931 26911
rect 11146 26908 11152 26920
rect 10919 26880 11152 26908
rect 10919 26877 10931 26880
rect 10873 26871 10931 26877
rect 10652 26868 10658 26871
rect 11146 26868 11152 26880
rect 11204 26908 11210 26920
rect 11330 26908 11336 26920
rect 11204 26880 11336 26908
rect 11204 26868 11210 26880
rect 11330 26868 11336 26880
rect 11388 26868 11394 26920
rect 11885 26911 11943 26917
rect 11885 26877 11897 26911
rect 11931 26908 11943 26911
rect 12526 26908 12532 26920
rect 11931 26880 12532 26908
rect 11931 26877 11943 26880
rect 11885 26871 11943 26877
rect 11900 26840 11928 26871
rect 12526 26868 12532 26880
rect 12584 26868 12590 26920
rect 13906 26868 13912 26920
rect 13964 26908 13970 26920
rect 14734 26908 14740 26920
rect 13964 26880 14740 26908
rect 13964 26868 13970 26880
rect 14734 26868 14740 26880
rect 14792 26868 14798 26920
rect 14826 26868 14832 26920
rect 14884 26868 14890 26920
rect 15013 26911 15071 26917
rect 15013 26877 15025 26911
rect 15059 26877 15071 26911
rect 15013 26871 15071 26877
rect 10336 26812 11928 26840
rect 11974 26800 11980 26852
rect 12032 26840 12038 26852
rect 12032 26812 12204 26840
rect 12032 26800 12038 26812
rect 5994 26732 6000 26784
rect 6052 26772 6058 26784
rect 6181 26775 6239 26781
rect 6181 26772 6193 26775
rect 6052 26744 6193 26772
rect 6052 26732 6058 26744
rect 6181 26741 6193 26744
rect 6227 26741 6239 26775
rect 6181 26735 6239 26741
rect 6454 26732 6460 26784
rect 6512 26772 6518 26784
rect 9766 26772 9772 26784
rect 6512 26744 9772 26772
rect 6512 26732 6518 26744
rect 9766 26732 9772 26744
rect 9824 26732 9830 26784
rect 10594 26732 10600 26784
rect 10652 26772 10658 26784
rect 10781 26775 10839 26781
rect 10781 26772 10793 26775
rect 10652 26744 10793 26772
rect 10652 26732 10658 26744
rect 10781 26741 10793 26744
rect 10827 26772 10839 26775
rect 11882 26772 11888 26784
rect 10827 26744 11888 26772
rect 10827 26741 10839 26744
rect 10781 26735 10839 26741
rect 11882 26732 11888 26744
rect 11940 26732 11946 26784
rect 12066 26732 12072 26784
rect 12124 26732 12130 26784
rect 12176 26772 12204 26812
rect 13262 26800 13268 26852
rect 13320 26840 13326 26852
rect 13357 26843 13415 26849
rect 13357 26840 13369 26843
rect 13320 26812 13369 26840
rect 13320 26800 13326 26812
rect 13357 26809 13369 26812
rect 13403 26809 13415 26843
rect 15028 26840 15056 26871
rect 15102 26868 15108 26920
rect 15160 26868 15166 26920
rect 15381 26843 15439 26849
rect 15381 26840 15393 26843
rect 13357 26803 13415 26809
rect 14108 26812 14964 26840
rect 15028 26812 15393 26840
rect 14108 26772 14136 26812
rect 14936 26784 14964 26812
rect 15381 26809 15393 26812
rect 15427 26809 15439 26843
rect 15381 26803 15439 26809
rect 12176 26744 14136 26772
rect 14182 26732 14188 26784
rect 14240 26772 14246 26784
rect 14645 26775 14703 26781
rect 14645 26772 14657 26775
rect 14240 26744 14657 26772
rect 14240 26732 14246 26744
rect 14645 26741 14657 26744
rect 14691 26741 14703 26775
rect 14645 26735 14703 26741
rect 14918 26732 14924 26784
rect 14976 26772 14982 26784
rect 15488 26772 15516 26939
rect 16206 26936 16212 26948
rect 16264 26936 16270 26988
rect 16758 26936 16764 26988
rect 16816 26985 16822 26988
rect 16816 26979 16865 26985
rect 16816 26945 16819 26979
rect 16853 26945 16865 26979
rect 16816 26939 16865 26945
rect 16816 26936 16822 26939
rect 16942 26936 16948 26988
rect 17000 26936 17006 26988
rect 17037 26979 17095 26985
rect 17037 26945 17049 26979
rect 17083 26945 17095 26979
rect 17218 26976 17224 26988
rect 17179 26948 17224 26976
rect 17037 26939 17095 26945
rect 16390 26868 16396 26920
rect 16448 26908 16454 26920
rect 17052 26908 17080 26939
rect 17218 26936 17224 26948
rect 17276 26936 17282 26988
rect 17310 26936 17316 26988
rect 17368 26936 17374 26988
rect 17681 26979 17739 26985
rect 17681 26945 17693 26979
rect 17727 26976 17739 26979
rect 17770 26976 17776 26988
rect 17727 26948 17776 26976
rect 17727 26945 17739 26948
rect 17681 26939 17739 26945
rect 17770 26936 17776 26948
rect 17828 26936 17834 26988
rect 17865 26979 17923 26985
rect 17865 26945 17877 26979
rect 17911 26976 17923 26979
rect 17911 26948 18276 26976
rect 17911 26945 17923 26948
rect 17865 26939 17923 26945
rect 18046 26908 18052 26920
rect 16448 26880 18052 26908
rect 16448 26868 16454 26880
rect 18046 26868 18052 26880
rect 18104 26868 18110 26920
rect 18248 26840 18276 26948
rect 18322 26936 18328 26988
rect 18380 26936 18386 26988
rect 18432 26985 18460 27016
rect 18690 27004 18696 27056
rect 18748 27044 18754 27056
rect 18969 27047 19027 27053
rect 18969 27044 18981 27047
rect 18748 27016 18981 27044
rect 18748 27004 18754 27016
rect 18969 27013 18981 27016
rect 19015 27013 19027 27047
rect 18969 27007 19027 27013
rect 18417 26979 18475 26985
rect 18417 26945 18429 26979
rect 18463 26945 18475 26979
rect 18417 26939 18475 26945
rect 18509 26979 18567 26985
rect 18509 26945 18521 26979
rect 18555 26945 18567 26979
rect 18509 26939 18567 26945
rect 18601 26979 18659 26985
rect 18601 26945 18613 26979
rect 18647 26976 18659 26979
rect 18647 26948 19104 26976
rect 18647 26945 18659 26948
rect 18601 26939 18659 26945
rect 18524 26908 18552 26939
rect 18690 26908 18696 26920
rect 18524 26880 18696 26908
rect 18690 26868 18696 26880
rect 18748 26868 18754 26920
rect 18782 26868 18788 26920
rect 18840 26868 18846 26920
rect 19076 26908 19104 26948
rect 19150 26936 19156 26988
rect 19208 26976 19214 26988
rect 19536 26976 19564 27084
rect 19702 27072 19708 27124
rect 19760 27112 19766 27124
rect 19797 27115 19855 27121
rect 19797 27112 19809 27115
rect 19760 27084 19809 27112
rect 19760 27072 19766 27084
rect 19797 27081 19809 27084
rect 19843 27081 19855 27115
rect 19797 27075 19855 27081
rect 19886 27072 19892 27124
rect 19944 27112 19950 27124
rect 20165 27115 20223 27121
rect 20165 27112 20177 27115
rect 19944 27084 20177 27112
rect 19944 27072 19950 27084
rect 20165 27081 20177 27084
rect 20211 27081 20223 27115
rect 20165 27075 20223 27081
rect 20806 27072 20812 27124
rect 20864 27072 20870 27124
rect 22557 27115 22615 27121
rect 22557 27081 22569 27115
rect 22603 27112 22615 27115
rect 24118 27112 24124 27124
rect 22603 27084 24124 27112
rect 22603 27081 22615 27084
rect 22557 27075 22615 27081
rect 24118 27072 24124 27084
rect 24176 27072 24182 27124
rect 25958 27112 25964 27124
rect 24780 27084 25964 27112
rect 19613 27047 19671 27053
rect 19613 27013 19625 27047
rect 19659 27044 19671 27047
rect 23201 27047 23259 27053
rect 19659 27016 20300 27044
rect 19659 27013 19671 27016
rect 19613 27007 19671 27013
rect 20272 26988 20300 27016
rect 20548 27016 23060 27044
rect 19797 26979 19855 26985
rect 19797 26976 19809 26979
rect 19208 26948 19380 26976
rect 19536 26948 19809 26976
rect 19208 26936 19214 26948
rect 19242 26908 19248 26920
rect 19076 26880 19248 26908
rect 19242 26868 19248 26880
rect 19300 26868 19306 26920
rect 19352 26908 19380 26948
rect 19797 26945 19809 26948
rect 19843 26976 19855 26979
rect 19886 26976 19892 26988
rect 19843 26948 19892 26976
rect 19843 26945 19855 26948
rect 19797 26939 19855 26945
rect 19886 26936 19892 26948
rect 19944 26936 19950 26988
rect 19981 26979 20039 26985
rect 19981 26945 19993 26979
rect 20027 26976 20039 26979
rect 20070 26976 20076 26988
rect 20027 26948 20076 26976
rect 20027 26945 20039 26948
rect 19981 26939 20039 26945
rect 20070 26936 20076 26948
rect 20128 26936 20134 26988
rect 20254 26936 20260 26988
rect 20312 26976 20318 26988
rect 20548 26985 20576 27016
rect 20349 26979 20407 26985
rect 20349 26976 20361 26979
rect 20312 26948 20361 26976
rect 20312 26936 20318 26948
rect 20349 26945 20361 26948
rect 20395 26945 20407 26979
rect 20349 26939 20407 26945
rect 20533 26979 20591 26985
rect 20533 26945 20545 26979
rect 20579 26945 20591 26979
rect 20533 26939 20591 26945
rect 20622 26936 20628 26988
rect 20680 26976 20686 26988
rect 21085 26979 21143 26985
rect 21085 26976 21097 26979
rect 20680 26948 21097 26976
rect 20680 26936 20686 26948
rect 21085 26945 21097 26948
rect 21131 26945 21143 26979
rect 21085 26939 21143 26945
rect 21818 26936 21824 26988
rect 21876 26976 21882 26988
rect 22005 26979 22063 26985
rect 22005 26976 22017 26979
rect 21876 26948 22017 26976
rect 21876 26936 21882 26948
rect 22005 26945 22017 26948
rect 22051 26945 22063 26979
rect 22005 26939 22063 26945
rect 22186 26936 22192 26988
rect 22244 26936 22250 26988
rect 22480 26985 22508 27016
rect 22465 26979 22523 26985
rect 22465 26945 22477 26979
rect 22511 26976 22523 26979
rect 22511 26948 22545 26976
rect 22511 26945 22523 26948
rect 22465 26939 22523 26945
rect 20901 26911 20959 26917
rect 20901 26908 20913 26911
rect 19352 26880 20913 26908
rect 20901 26877 20913 26880
rect 20947 26877 20959 26911
rect 20901 26871 20959 26877
rect 21361 26911 21419 26917
rect 21361 26877 21373 26911
rect 21407 26908 21419 26911
rect 21450 26908 21456 26920
rect 21407 26880 21456 26908
rect 21407 26877 21419 26880
rect 21361 26871 21419 26877
rect 21450 26868 21456 26880
rect 21508 26868 21514 26920
rect 18598 26840 18604 26852
rect 18248 26812 18604 26840
rect 18598 26800 18604 26812
rect 18656 26840 18662 26852
rect 21821 26843 21879 26849
rect 21821 26840 21833 26843
rect 18656 26812 21833 26840
rect 18656 26800 18662 26812
rect 21821 26809 21833 26812
rect 21867 26809 21879 26843
rect 22480 26840 22508 26939
rect 22646 26936 22652 26988
rect 22704 26936 22710 26988
rect 22738 26936 22744 26988
rect 22796 26976 22802 26988
rect 22925 26979 22983 26985
rect 22925 26976 22937 26979
rect 22796 26948 22937 26976
rect 22796 26936 22802 26948
rect 22925 26945 22937 26948
rect 22971 26945 22983 26979
rect 23032 26976 23060 27016
rect 23201 27013 23213 27047
rect 23247 27044 23259 27047
rect 24780 27044 24808 27084
rect 25958 27072 25964 27084
rect 26016 27072 26022 27124
rect 29825 27115 29883 27121
rect 29825 27081 29837 27115
rect 29871 27112 29883 27115
rect 30006 27112 30012 27124
rect 29871 27084 30012 27112
rect 29871 27081 29883 27084
rect 29825 27075 29883 27081
rect 30006 27072 30012 27084
rect 30064 27072 30070 27124
rect 30193 27115 30251 27121
rect 30193 27081 30205 27115
rect 30239 27112 30251 27115
rect 31018 27112 31024 27124
rect 30239 27084 31024 27112
rect 30239 27081 30251 27084
rect 30193 27075 30251 27081
rect 23247 27016 24808 27044
rect 24857 27047 24915 27053
rect 23247 27013 23259 27016
rect 23201 27007 23259 27013
rect 24857 27013 24869 27047
rect 24903 27044 24915 27047
rect 25222 27044 25228 27056
rect 24903 27016 25228 27044
rect 24903 27013 24915 27016
rect 24857 27007 24915 27013
rect 25222 27004 25228 27016
rect 25280 27004 25286 27056
rect 28626 27004 28632 27056
rect 28684 27044 28690 27056
rect 30208 27044 30236 27075
rect 31018 27072 31024 27084
rect 31076 27072 31082 27124
rect 31110 27072 31116 27124
rect 31168 27112 31174 27124
rect 31205 27115 31263 27121
rect 31205 27112 31217 27115
rect 31168 27084 31217 27112
rect 31168 27072 31174 27084
rect 31205 27081 31217 27084
rect 31251 27081 31263 27115
rect 31205 27075 31263 27081
rect 31389 27115 31447 27121
rect 31389 27081 31401 27115
rect 31435 27112 31447 27115
rect 31570 27112 31576 27124
rect 31435 27084 31576 27112
rect 31435 27081 31447 27084
rect 31389 27075 31447 27081
rect 31570 27072 31576 27084
rect 31628 27112 31634 27124
rect 36538 27112 36544 27124
rect 31628 27084 34652 27112
rect 31628 27072 31634 27084
rect 28684 27016 30236 27044
rect 31680 27016 31984 27044
rect 28684 27004 28690 27016
rect 23032 26948 23208 26976
rect 22925 26939 22983 26945
rect 22664 26908 22692 26936
rect 23017 26911 23075 26917
rect 23017 26908 23029 26911
rect 22664 26880 23029 26908
rect 23017 26877 23029 26880
rect 23063 26877 23075 26911
rect 23180 26908 23208 26948
rect 23290 26936 23296 26988
rect 23348 26936 23354 26988
rect 24118 26936 24124 26988
rect 24176 26976 24182 26988
rect 24489 26979 24547 26985
rect 24489 26976 24501 26979
rect 24176 26948 24501 26976
rect 24176 26936 24182 26948
rect 24489 26945 24501 26948
rect 24535 26945 24547 26979
rect 24489 26939 24547 26945
rect 24765 26979 24823 26985
rect 24765 26945 24777 26979
rect 24811 26976 24823 26979
rect 25314 26976 25320 26988
rect 24811 26948 25320 26976
rect 24811 26945 24823 26948
rect 24765 26939 24823 26945
rect 25314 26936 25320 26948
rect 25372 26936 25378 26988
rect 25593 26979 25651 26985
rect 25593 26945 25605 26979
rect 25639 26945 25651 26979
rect 25593 26939 25651 26945
rect 23385 26911 23443 26917
rect 23385 26908 23397 26911
rect 23180 26880 23397 26908
rect 23017 26871 23075 26877
rect 23385 26877 23397 26880
rect 23431 26908 23443 26911
rect 23474 26908 23480 26920
rect 23431 26880 23480 26908
rect 23431 26877 23443 26880
rect 23385 26871 23443 26877
rect 22480 26812 22876 26840
rect 21821 26803 21879 26809
rect 14976 26744 15516 26772
rect 20441 26775 20499 26781
rect 14976 26732 14982 26744
rect 20441 26741 20453 26775
rect 20487 26772 20499 26775
rect 20714 26772 20720 26784
rect 20487 26744 20720 26772
rect 20487 26741 20499 26744
rect 20441 26735 20499 26741
rect 20714 26732 20720 26744
rect 20772 26732 20778 26784
rect 21269 26775 21327 26781
rect 21269 26741 21281 26775
rect 21315 26772 21327 26775
rect 21358 26772 21364 26784
rect 21315 26744 21364 26772
rect 21315 26741 21327 26744
rect 21269 26735 21327 26741
rect 21358 26732 21364 26744
rect 21416 26732 21422 26784
rect 22738 26732 22744 26784
rect 22796 26732 22802 26784
rect 22848 26772 22876 26812
rect 22925 26775 22983 26781
rect 22925 26772 22937 26775
rect 22848 26744 22937 26772
rect 22925 26741 22937 26744
rect 22971 26741 22983 26775
rect 23032 26772 23060 26871
rect 23474 26868 23480 26880
rect 23532 26868 23538 26920
rect 24397 26911 24455 26917
rect 24397 26877 24409 26911
rect 24443 26908 24455 26911
rect 24578 26908 24584 26920
rect 24443 26880 24584 26908
rect 24443 26877 24455 26880
rect 24397 26871 24455 26877
rect 24578 26868 24584 26880
rect 24636 26868 24642 26920
rect 24670 26868 24676 26920
rect 24728 26908 24734 26920
rect 25409 26911 25467 26917
rect 25409 26908 25421 26911
rect 24728 26880 25421 26908
rect 24728 26868 24734 26880
rect 25409 26877 25421 26880
rect 25455 26877 25467 26911
rect 25409 26871 25467 26877
rect 23198 26800 23204 26852
rect 23256 26840 23262 26852
rect 23661 26843 23719 26849
rect 23661 26840 23673 26843
rect 23256 26812 23673 26840
rect 23256 26800 23262 26812
rect 23661 26809 23673 26812
rect 23707 26840 23719 26843
rect 25608 26840 25636 26939
rect 25774 26936 25780 26988
rect 25832 26936 25838 26988
rect 25869 26979 25927 26985
rect 25869 26945 25881 26979
rect 25915 26976 25927 26979
rect 26786 26976 26792 26988
rect 25915 26948 26792 26976
rect 25915 26945 25927 26948
rect 25869 26939 25927 26945
rect 26786 26936 26792 26948
rect 26844 26936 26850 26988
rect 30742 26936 30748 26988
rect 30800 26976 30806 26988
rect 31680 26985 31708 27016
rect 31956 26988 31984 27016
rect 32122 27004 32128 27056
rect 32180 27004 32186 27056
rect 32309 27047 32367 27053
rect 32309 27013 32321 27047
rect 32355 27013 32367 27047
rect 32309 27007 32367 27013
rect 30837 26979 30895 26985
rect 30837 26976 30849 26979
rect 30800 26948 30849 26976
rect 30800 26936 30806 26948
rect 30837 26945 30849 26948
rect 30883 26945 30895 26979
rect 30837 26939 30895 26945
rect 31665 26979 31723 26985
rect 31665 26945 31677 26979
rect 31711 26945 31723 26979
rect 31665 26939 31723 26945
rect 31754 26936 31760 26988
rect 31812 26936 31818 26988
rect 31938 26936 31944 26988
rect 31996 26936 32002 26988
rect 32324 26976 32352 27007
rect 32048 26948 32352 26976
rect 32048 26920 32076 26948
rect 34422 26936 34428 26988
rect 34480 26936 34486 26988
rect 34624 26985 34652 27084
rect 36372 27084 36544 27112
rect 34609 26979 34667 26985
rect 34609 26945 34621 26979
rect 34655 26976 34667 26979
rect 36173 26979 36231 26985
rect 36173 26976 36185 26979
rect 34655 26948 36185 26976
rect 34655 26945 34667 26948
rect 34609 26939 34667 26945
rect 36173 26945 36185 26948
rect 36219 26945 36231 26979
rect 36173 26939 36231 26945
rect 36265 26979 36323 26985
rect 36265 26945 36277 26979
rect 36311 26945 36323 26979
rect 36372 26976 36400 27084
rect 36538 27072 36544 27084
rect 36596 27112 36602 27124
rect 36596 27084 37596 27112
rect 36596 27072 36602 27084
rect 37568 27056 37596 27084
rect 37826 27072 37832 27124
rect 37884 27112 37890 27124
rect 38010 27112 38016 27124
rect 37884 27084 38016 27112
rect 37884 27072 37890 27084
rect 38010 27072 38016 27084
rect 38068 27112 38074 27124
rect 38105 27115 38163 27121
rect 38105 27112 38117 27115
rect 38068 27084 38117 27112
rect 38068 27072 38074 27084
rect 38105 27081 38117 27084
rect 38151 27081 38163 27115
rect 38105 27075 38163 27081
rect 38746 27072 38752 27124
rect 38804 27112 38810 27124
rect 40037 27115 40095 27121
rect 40037 27112 40049 27115
rect 38804 27084 40049 27112
rect 38804 27072 38810 27084
rect 40037 27081 40049 27084
rect 40083 27081 40095 27115
rect 40037 27075 40095 27081
rect 36449 27047 36507 27053
rect 36449 27013 36461 27047
rect 36495 27044 36507 27047
rect 36495 27016 37504 27044
rect 36495 27013 36507 27016
rect 36449 27007 36507 27013
rect 37476 26988 37504 27016
rect 37550 27004 37556 27056
rect 37608 27004 37614 27056
rect 39209 27047 39267 27053
rect 39209 27044 39221 27047
rect 37936 27016 38976 27044
rect 36541 26979 36599 26985
rect 36541 26976 36553 26979
rect 36372 26948 36553 26976
rect 36265 26939 36323 26945
rect 36541 26945 36553 26948
rect 36587 26945 36599 26979
rect 36541 26939 36599 26945
rect 36725 26979 36783 26985
rect 36725 26945 36737 26979
rect 36771 26945 36783 26979
rect 36725 26939 36783 26945
rect 30006 26868 30012 26920
rect 30064 26908 30070 26920
rect 30285 26911 30343 26917
rect 30285 26908 30297 26911
rect 30064 26880 30297 26908
rect 30064 26868 30070 26880
rect 30285 26877 30297 26880
rect 30331 26877 30343 26911
rect 30285 26871 30343 26877
rect 30377 26911 30435 26917
rect 30377 26877 30389 26911
rect 30423 26877 30435 26911
rect 32030 26908 32036 26920
rect 30377 26871 30435 26877
rect 31220 26880 32036 26908
rect 23707 26812 25636 26840
rect 23707 26809 23719 26812
rect 23661 26803 23719 26809
rect 29914 26800 29920 26852
rect 29972 26840 29978 26852
rect 30392 26840 30420 26871
rect 29972 26812 30420 26840
rect 29972 26800 29978 26812
rect 23293 26775 23351 26781
rect 23293 26772 23305 26775
rect 23032 26744 23305 26772
rect 22925 26735 22983 26741
rect 23293 26741 23305 26744
rect 23339 26741 23351 26775
rect 23293 26735 23351 26741
rect 24210 26732 24216 26784
rect 24268 26732 24274 26784
rect 31220 26781 31248 26880
rect 32030 26868 32036 26880
rect 32088 26868 32094 26920
rect 32582 26868 32588 26920
rect 32640 26908 32646 26920
rect 36280 26908 36308 26939
rect 36354 26908 36360 26920
rect 32640 26880 36360 26908
rect 32640 26868 32646 26880
rect 36354 26868 36360 26880
rect 36412 26868 36418 26920
rect 36740 26908 36768 26939
rect 36814 26936 36820 26988
rect 36872 26936 36878 26988
rect 36909 26979 36967 26985
rect 36909 26945 36921 26979
rect 36955 26976 36967 26979
rect 37090 26976 37096 26988
rect 36955 26948 37096 26976
rect 36955 26945 36967 26948
rect 36909 26939 36967 26945
rect 37090 26936 37096 26948
rect 37148 26936 37154 26988
rect 37458 26936 37464 26988
rect 37516 26936 37522 26988
rect 37642 26936 37648 26988
rect 37700 26936 37706 26988
rect 37734 26936 37740 26988
rect 37792 26985 37798 26988
rect 37936 26985 37964 27016
rect 38948 26988 38976 27016
rect 39040 27016 39221 27044
rect 37792 26979 37821 26985
rect 37809 26945 37821 26979
rect 37792 26939 37821 26945
rect 37921 26979 37979 26985
rect 37921 26945 37933 26979
rect 37967 26945 37979 26979
rect 37921 26939 37979 26945
rect 37792 26936 37798 26939
rect 36464 26880 36768 26908
rect 36832 26908 36860 26936
rect 37936 26908 37964 26939
rect 38378 26936 38384 26988
rect 38436 26936 38442 26988
rect 38654 26936 38660 26988
rect 38712 26936 38718 26988
rect 38930 26936 38936 26988
rect 38988 26936 38994 26988
rect 36832 26880 37964 26908
rect 31849 26843 31907 26849
rect 31849 26809 31861 26843
rect 31895 26840 31907 26843
rect 34054 26840 34060 26852
rect 31895 26812 34060 26840
rect 31895 26809 31907 26812
rect 31849 26803 31907 26809
rect 34054 26800 34060 26812
rect 34112 26840 34118 26852
rect 35526 26840 35532 26852
rect 34112 26812 35532 26840
rect 34112 26800 34118 26812
rect 35526 26800 35532 26812
rect 35584 26800 35590 26852
rect 36464 26849 36492 26880
rect 38746 26868 38752 26920
rect 38804 26868 38810 26920
rect 38838 26868 38844 26920
rect 38896 26868 38902 26920
rect 36449 26843 36507 26849
rect 36449 26809 36461 26843
rect 36495 26809 36507 26843
rect 36449 26803 36507 26809
rect 37093 26843 37151 26849
rect 37093 26809 37105 26843
rect 37139 26840 37151 26843
rect 38010 26840 38016 26852
rect 37139 26812 38016 26840
rect 37139 26809 37151 26812
rect 37093 26803 37151 26809
rect 38010 26800 38016 26812
rect 38068 26800 38074 26852
rect 38286 26800 38292 26852
rect 38344 26840 38350 26852
rect 39040 26840 39068 27016
rect 39209 27013 39221 27016
rect 39255 27013 39267 27047
rect 39209 27007 39267 27013
rect 39298 27004 39304 27056
rect 39356 27044 39362 27056
rect 39393 27047 39451 27053
rect 39393 27044 39405 27047
rect 39356 27016 39405 27044
rect 39356 27004 39362 27016
rect 39393 27013 39405 27016
rect 39439 27013 39451 27047
rect 39393 27007 39451 27013
rect 39669 26979 39727 26985
rect 39669 26945 39681 26979
rect 39715 26976 39727 26979
rect 39758 26976 39764 26988
rect 39715 26948 39764 26976
rect 39715 26945 39727 26948
rect 39669 26939 39727 26945
rect 39758 26936 39764 26948
rect 39816 26936 39822 26988
rect 40218 26936 40224 26988
rect 40276 26936 40282 26988
rect 38344 26812 39068 26840
rect 39117 26843 39175 26849
rect 38344 26800 38350 26812
rect 39117 26809 39129 26843
rect 39163 26840 39175 26843
rect 39850 26840 39856 26852
rect 39163 26812 39856 26840
rect 39163 26809 39175 26812
rect 39117 26803 39175 26809
rect 39850 26800 39856 26812
rect 39908 26800 39914 26852
rect 31205 26775 31263 26781
rect 31205 26741 31217 26775
rect 31251 26741 31263 26775
rect 31205 26735 31263 26741
rect 32306 26732 32312 26784
rect 32364 26732 32370 26784
rect 32493 26775 32551 26781
rect 32493 26741 32505 26775
rect 32539 26772 32551 26775
rect 34422 26772 34428 26784
rect 32539 26744 34428 26772
rect 32539 26741 32551 26744
rect 32493 26735 32551 26741
rect 34422 26732 34428 26744
rect 34480 26732 34486 26784
rect 34609 26775 34667 26781
rect 34609 26741 34621 26775
rect 34655 26772 34667 26775
rect 35342 26772 35348 26784
rect 34655 26744 35348 26772
rect 34655 26741 34667 26744
rect 34609 26735 34667 26741
rect 35342 26732 35348 26744
rect 35400 26732 35406 26784
rect 37277 26775 37335 26781
rect 37277 26741 37289 26775
rect 37323 26772 37335 26775
rect 37366 26772 37372 26784
rect 37323 26744 37372 26772
rect 37323 26741 37335 26744
rect 37277 26735 37335 26741
rect 37366 26732 37372 26744
rect 37424 26732 37430 26784
rect 38838 26732 38844 26784
rect 38896 26772 38902 26784
rect 39206 26772 39212 26784
rect 38896 26744 39212 26772
rect 38896 26732 38902 26744
rect 39206 26732 39212 26744
rect 39264 26772 39270 26784
rect 39393 26775 39451 26781
rect 39393 26772 39405 26775
rect 39264 26744 39405 26772
rect 39264 26732 39270 26744
rect 39393 26741 39405 26744
rect 39439 26741 39451 26775
rect 39393 26735 39451 26741
rect 1104 26682 40572 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 40572 26682
rect 1104 26608 40572 26630
rect 3050 26528 3056 26580
rect 3108 26568 3114 26580
rect 5258 26568 5264 26580
rect 3108 26540 5264 26568
rect 3108 26528 3114 26540
rect 5258 26528 5264 26540
rect 5316 26528 5322 26580
rect 5350 26528 5356 26580
rect 5408 26568 5414 26580
rect 6454 26568 6460 26580
rect 5408 26540 6460 26568
rect 5408 26528 5414 26540
rect 6454 26528 6460 26540
rect 6512 26528 6518 26580
rect 6641 26571 6699 26577
rect 6641 26537 6653 26571
rect 6687 26568 6699 26571
rect 6822 26568 6828 26580
rect 6687 26540 6828 26568
rect 6687 26537 6699 26540
rect 6641 26531 6699 26537
rect 6822 26528 6828 26540
rect 6880 26528 6886 26580
rect 8665 26571 8723 26577
rect 8665 26537 8677 26571
rect 8711 26568 8723 26571
rect 9306 26568 9312 26580
rect 8711 26540 9312 26568
rect 8711 26537 8723 26540
rect 8665 26531 8723 26537
rect 9306 26528 9312 26540
rect 9364 26528 9370 26580
rect 10502 26568 10508 26580
rect 9416 26540 10508 26568
rect 2774 26392 2780 26444
rect 2832 26432 2838 26444
rect 3142 26432 3148 26444
rect 2832 26404 3148 26432
rect 2832 26392 2838 26404
rect 3142 26392 3148 26404
rect 3200 26392 3206 26444
rect 3329 26435 3387 26441
rect 3329 26401 3341 26435
rect 3375 26432 3387 26435
rect 5258 26432 5264 26444
rect 3375 26404 5264 26432
rect 3375 26401 3387 26404
rect 3329 26395 3387 26401
rect 5258 26392 5264 26404
rect 5316 26392 5322 26444
rect 4338 26324 4344 26376
rect 4396 26324 4402 26376
rect 5368 26373 5396 26528
rect 5905 26503 5963 26509
rect 5905 26469 5917 26503
rect 5951 26500 5963 26503
rect 7006 26500 7012 26512
rect 5951 26472 7012 26500
rect 5951 26469 5963 26472
rect 5905 26463 5963 26469
rect 7006 26460 7012 26472
rect 7064 26460 7070 26512
rect 8938 26460 8944 26512
rect 8996 26460 9002 26512
rect 6362 26432 6368 26444
rect 5736 26404 6368 26432
rect 5736 26373 5764 26404
rect 6362 26392 6368 26404
rect 6420 26392 6426 26444
rect 6638 26392 6644 26444
rect 6696 26432 6702 26444
rect 6733 26435 6791 26441
rect 6733 26432 6745 26435
rect 6696 26404 6745 26432
rect 6696 26392 6702 26404
rect 6733 26401 6745 26404
rect 6779 26401 6791 26435
rect 9416 26432 9444 26540
rect 10502 26528 10508 26540
rect 10560 26528 10566 26580
rect 10594 26528 10600 26580
rect 10652 26528 10658 26580
rect 10778 26528 10784 26580
rect 10836 26568 10842 26580
rect 10965 26571 11023 26577
rect 10965 26568 10977 26571
rect 10836 26540 10977 26568
rect 10836 26528 10842 26540
rect 10965 26537 10977 26540
rect 11011 26537 11023 26571
rect 11241 26571 11299 26577
rect 11241 26568 11253 26571
rect 10965 26531 11023 26537
rect 11072 26540 11253 26568
rect 10137 26503 10195 26509
rect 10137 26469 10149 26503
rect 10183 26500 10195 26503
rect 10226 26500 10232 26512
rect 10183 26472 10232 26500
rect 10183 26469 10195 26472
rect 10137 26463 10195 26469
rect 10226 26460 10232 26472
rect 10284 26460 10290 26512
rect 10870 26460 10876 26512
rect 10928 26500 10934 26512
rect 11072 26500 11100 26540
rect 11241 26537 11253 26540
rect 11287 26537 11299 26571
rect 11241 26531 11299 26537
rect 12066 26528 12072 26580
rect 12124 26528 12130 26580
rect 12250 26528 12256 26580
rect 12308 26528 12314 26580
rect 12618 26528 12624 26580
rect 12676 26528 12682 26580
rect 14274 26568 14280 26580
rect 13372 26540 14280 26568
rect 11698 26500 11704 26512
rect 10928 26472 11100 26500
rect 11240 26472 11704 26500
rect 10928 26460 10934 26472
rect 6733 26395 6791 26401
rect 8312 26404 9444 26432
rect 5353 26367 5411 26373
rect 5353 26333 5365 26367
rect 5399 26333 5411 26367
rect 5353 26327 5411 26333
rect 5721 26367 5779 26373
rect 5721 26333 5733 26367
rect 5767 26333 5779 26367
rect 5721 26327 5779 26333
rect 5994 26324 6000 26376
rect 6052 26324 6058 26376
rect 6086 26324 6092 26376
rect 6144 26324 6150 26376
rect 6503 26367 6561 26373
rect 6503 26333 6515 26367
rect 6549 26364 6561 26367
rect 6822 26364 6828 26376
rect 6549 26336 6828 26364
rect 6549 26333 6561 26336
rect 6503 26327 6561 26333
rect 6822 26324 6828 26336
rect 6880 26324 6886 26376
rect 6917 26367 6975 26373
rect 6917 26333 6929 26367
rect 6963 26364 6975 26367
rect 7282 26364 7288 26376
rect 6963 26336 7288 26364
rect 6963 26333 6975 26336
rect 6917 26327 6975 26333
rect 7282 26324 7288 26336
rect 7340 26324 7346 26376
rect 8018 26324 8024 26376
rect 8076 26324 8082 26376
rect 8169 26367 8227 26373
rect 8169 26333 8181 26367
rect 8215 26364 8227 26367
rect 8312 26364 8340 26404
rect 9490 26392 9496 26444
rect 9548 26432 9554 26444
rect 10962 26432 10968 26444
rect 9548 26404 9996 26432
rect 9548 26392 9554 26404
rect 8215 26336 8340 26364
rect 8215 26333 8227 26336
rect 8169 26327 8227 26333
rect 8386 26324 8392 26376
rect 8444 26324 8450 26376
rect 8478 26324 8484 26376
rect 8536 26373 8542 26376
rect 8536 26367 8585 26373
rect 8536 26333 8539 26367
rect 8573 26364 8585 26367
rect 8573 26336 9260 26364
rect 8573 26333 8585 26336
rect 8536 26327 8585 26333
rect 8536 26324 8542 26327
rect 3053 26299 3111 26305
rect 3053 26265 3065 26299
rect 3099 26296 3111 26299
rect 3789 26299 3847 26305
rect 3789 26296 3801 26299
rect 3099 26268 3801 26296
rect 3099 26265 3111 26268
rect 3053 26259 3111 26265
rect 3789 26265 3801 26268
rect 3835 26265 3847 26299
rect 3789 26259 3847 26265
rect 5537 26299 5595 26305
rect 5537 26265 5549 26299
rect 5583 26265 5595 26299
rect 5537 26259 5595 26265
rect 1854 26188 1860 26240
rect 1912 26228 1918 26240
rect 2685 26231 2743 26237
rect 2685 26228 2697 26231
rect 1912 26200 2697 26228
rect 1912 26188 1918 26200
rect 2685 26197 2697 26200
rect 2731 26197 2743 26231
rect 5552 26228 5580 26259
rect 5626 26256 5632 26308
rect 5684 26256 5690 26308
rect 6270 26256 6276 26308
rect 6328 26256 6334 26308
rect 6365 26299 6423 26305
rect 6365 26265 6377 26299
rect 6411 26296 6423 26299
rect 6730 26296 6736 26308
rect 6411 26268 6736 26296
rect 6411 26265 6423 26268
rect 6365 26259 6423 26265
rect 6730 26256 6736 26268
rect 6788 26256 6794 26308
rect 7098 26256 7104 26308
rect 7156 26256 7162 26308
rect 8297 26299 8355 26305
rect 8297 26296 8309 26299
rect 8220 26268 8309 26296
rect 8220 26240 8248 26268
rect 8297 26265 8309 26268
rect 8343 26265 8355 26299
rect 8297 26259 8355 26265
rect 9030 26256 9036 26308
rect 9088 26296 9094 26308
rect 9125 26299 9183 26305
rect 9125 26296 9137 26299
rect 9088 26268 9137 26296
rect 9088 26256 9094 26268
rect 9125 26265 9137 26268
rect 9171 26265 9183 26299
rect 9232 26296 9260 26336
rect 9306 26324 9312 26376
rect 9364 26324 9370 26376
rect 9968 26373 9996 26404
rect 10152 26404 10968 26432
rect 10152 26373 10180 26404
rect 10962 26392 10968 26404
rect 11020 26392 11026 26444
rect 9861 26367 9919 26373
rect 9861 26333 9873 26367
rect 9907 26333 9919 26367
rect 9861 26327 9919 26333
rect 9953 26367 10011 26373
rect 9953 26333 9965 26367
rect 9999 26333 10011 26367
rect 9953 26327 10011 26333
rect 10137 26367 10195 26373
rect 10137 26333 10149 26367
rect 10183 26333 10195 26367
rect 10137 26327 10195 26333
rect 9490 26296 9496 26308
rect 9232 26268 9496 26296
rect 9125 26259 9183 26265
rect 9490 26256 9496 26268
rect 9548 26256 9554 26308
rect 9876 26296 9904 26327
rect 10318 26324 10324 26376
rect 10376 26364 10382 26376
rect 10597 26367 10655 26373
rect 10597 26364 10609 26367
rect 10376 26336 10609 26364
rect 10376 26324 10382 26336
rect 10597 26333 10609 26336
rect 10643 26333 10655 26367
rect 10597 26327 10655 26333
rect 10781 26367 10839 26373
rect 10781 26333 10793 26367
rect 10827 26364 10839 26367
rect 11146 26364 11152 26376
rect 10827 26336 11152 26364
rect 10827 26333 10839 26336
rect 10781 26327 10839 26333
rect 11146 26324 11152 26336
rect 11204 26324 11210 26376
rect 11240 26373 11268 26472
rect 11698 26460 11704 26472
rect 11756 26460 11762 26512
rect 11977 26503 12035 26509
rect 11977 26469 11989 26503
rect 12023 26500 12035 26503
rect 13372 26500 13400 26540
rect 14274 26528 14280 26540
rect 14332 26528 14338 26580
rect 14550 26528 14556 26580
rect 14608 26528 14614 26580
rect 14826 26528 14832 26580
rect 14884 26568 14890 26580
rect 16853 26571 16911 26577
rect 16853 26568 16865 26571
rect 14884 26540 16865 26568
rect 14884 26528 14890 26540
rect 16853 26537 16865 26540
rect 16899 26537 16911 26571
rect 16853 26531 16911 26537
rect 18322 26528 18328 26580
rect 18380 26568 18386 26580
rect 18601 26571 18659 26577
rect 18601 26568 18613 26571
rect 18380 26540 18613 26568
rect 18380 26528 18386 26540
rect 18601 26537 18613 26540
rect 18647 26537 18659 26571
rect 18601 26531 18659 26537
rect 18690 26528 18696 26580
rect 18748 26568 18754 26580
rect 19150 26568 19156 26580
rect 18748 26540 19156 26568
rect 18748 26528 18754 26540
rect 19150 26528 19156 26540
rect 19208 26528 19214 26580
rect 20070 26528 20076 26580
rect 20128 26568 20134 26580
rect 20257 26571 20315 26577
rect 20257 26568 20269 26571
rect 20128 26540 20269 26568
rect 20128 26528 20134 26540
rect 20257 26537 20269 26540
rect 20303 26537 20315 26571
rect 20257 26531 20315 26537
rect 22462 26528 22468 26580
rect 22520 26528 22526 26580
rect 22646 26528 22652 26580
rect 22704 26568 22710 26580
rect 22922 26568 22928 26580
rect 22704 26540 22928 26568
rect 22704 26528 22710 26540
rect 22922 26528 22928 26540
rect 22980 26568 22986 26580
rect 23477 26571 23535 26577
rect 23477 26568 23489 26571
rect 22980 26540 23489 26568
rect 22980 26528 22986 26540
rect 23477 26537 23489 26540
rect 23523 26537 23535 26571
rect 23477 26531 23535 26537
rect 24026 26528 24032 26580
rect 24084 26568 24090 26580
rect 24397 26571 24455 26577
rect 24397 26568 24409 26571
rect 24084 26540 24409 26568
rect 24084 26528 24090 26540
rect 24397 26537 24409 26540
rect 24443 26537 24455 26571
rect 24397 26531 24455 26537
rect 24581 26571 24639 26577
rect 24581 26537 24593 26571
rect 24627 26537 24639 26571
rect 24581 26531 24639 26537
rect 12023 26472 13400 26500
rect 12023 26469 12035 26472
rect 11977 26463 12035 26469
rect 14090 26460 14096 26512
rect 14148 26460 14154 26512
rect 14568 26500 14596 26528
rect 15470 26500 15476 26512
rect 14471 26472 15476 26500
rect 11330 26392 11336 26444
rect 11388 26432 11394 26444
rect 14366 26432 14372 26444
rect 11388 26404 12480 26432
rect 11388 26392 11394 26404
rect 11440 26373 11468 26404
rect 12452 26376 12480 26404
rect 14287 26404 14372 26432
rect 11240 26367 11299 26373
rect 11240 26333 11253 26367
rect 11287 26333 11299 26367
rect 11240 26330 11299 26333
rect 11241 26327 11299 26330
rect 11425 26367 11483 26373
rect 11425 26333 11437 26367
rect 11471 26333 11483 26367
rect 11425 26327 11483 26333
rect 12069 26367 12127 26373
rect 12069 26333 12081 26367
rect 12115 26333 12127 26367
rect 12069 26327 12127 26333
rect 10042 26296 10048 26308
rect 9876 26268 10048 26296
rect 10042 26256 10048 26268
rect 10100 26296 10106 26308
rect 11054 26296 11060 26308
rect 10100 26268 11060 26296
rect 10100 26256 10106 26268
rect 11054 26256 11060 26268
rect 11112 26296 11118 26308
rect 11701 26299 11759 26305
rect 11701 26296 11713 26299
rect 11112 26268 11713 26296
rect 11112 26256 11118 26268
rect 11701 26265 11713 26268
rect 11747 26296 11759 26299
rect 11974 26296 11980 26308
rect 11747 26268 11980 26296
rect 11747 26265 11759 26268
rect 11701 26259 11759 26265
rect 11974 26256 11980 26268
rect 12032 26256 12038 26308
rect 12084 26296 12112 26327
rect 12158 26324 12164 26376
rect 12216 26364 12222 26376
rect 12253 26367 12311 26373
rect 12253 26364 12265 26367
rect 12216 26336 12265 26364
rect 12216 26324 12222 26336
rect 12253 26333 12265 26336
rect 12299 26333 12311 26367
rect 12253 26327 12311 26333
rect 12434 26324 12440 26376
rect 12492 26324 12498 26376
rect 14287 26373 14315 26404
rect 14366 26392 14372 26404
rect 14424 26392 14430 26444
rect 14471 26373 14499 26472
rect 15470 26460 15476 26472
rect 15528 26460 15534 26512
rect 20533 26503 20591 26509
rect 20533 26500 20545 26503
rect 18708 26472 20545 26500
rect 15575 26404 16625 26432
rect 14272 26367 14330 26373
rect 14272 26333 14284 26367
rect 14318 26333 14330 26367
rect 14272 26327 14330 26333
rect 14461 26367 14519 26373
rect 14461 26333 14473 26367
rect 14507 26333 14519 26367
rect 14642 26364 14648 26376
rect 14603 26336 14648 26364
rect 14461 26327 14519 26333
rect 12618 26296 12624 26308
rect 12084 26268 12624 26296
rect 12618 26256 12624 26268
rect 12676 26256 12682 26308
rect 14287 26240 14315 26327
rect 14642 26324 14648 26336
rect 14700 26324 14706 26376
rect 14734 26324 14740 26376
rect 14792 26324 14798 26376
rect 15575 26373 15603 26404
rect 15560 26367 15618 26373
rect 15560 26333 15572 26367
rect 15606 26333 15618 26367
rect 15560 26327 15618 26333
rect 14369 26299 14427 26305
rect 14369 26265 14381 26299
rect 14415 26296 14427 26299
rect 14826 26296 14832 26308
rect 14415 26268 14832 26296
rect 14415 26265 14427 26268
rect 14369 26259 14427 26265
rect 14826 26256 14832 26268
rect 14884 26256 14890 26308
rect 15575 26296 15603 26327
rect 15838 26324 15844 26376
rect 15896 26373 15902 26376
rect 15896 26367 15935 26373
rect 15923 26333 15935 26367
rect 15896 26327 15935 26333
rect 15896 26324 15902 26327
rect 16022 26324 16028 26376
rect 16080 26324 16086 26376
rect 16114 26324 16120 26376
rect 16172 26324 16178 26376
rect 16298 26373 16304 26376
rect 16265 26367 16304 26373
rect 16265 26333 16277 26367
rect 16265 26327 16304 26333
rect 16298 26324 16304 26327
rect 16356 26324 16362 26376
rect 16390 26324 16396 26376
rect 16448 26324 16454 26376
rect 16597 26373 16625 26404
rect 17256 26404 18184 26432
rect 16582 26367 16640 26373
rect 16582 26333 16594 26367
rect 16628 26364 16640 26367
rect 16758 26364 16764 26376
rect 16628 26336 16764 26364
rect 16628 26333 16640 26336
rect 16582 26327 16640 26333
rect 16758 26324 16764 26336
rect 16816 26364 16822 26376
rect 17256 26373 17284 26404
rect 18156 26376 18184 26404
rect 17241 26367 17299 26373
rect 17241 26364 17253 26367
rect 16816 26336 17253 26364
rect 16816 26324 16822 26336
rect 17241 26333 17253 26336
rect 17287 26333 17299 26367
rect 17241 26327 17299 26333
rect 17773 26367 17831 26373
rect 17773 26333 17785 26367
rect 17819 26364 17831 26367
rect 18046 26364 18052 26376
rect 17819 26336 18052 26364
rect 17819 26333 17831 26336
rect 17773 26327 17831 26333
rect 14936 26268 15603 26296
rect 5810 26228 5816 26240
rect 5552 26200 5816 26228
rect 2685 26191 2743 26197
rect 5810 26188 5816 26200
rect 5868 26228 5874 26240
rect 8202 26228 8208 26240
rect 5868 26200 8208 26228
rect 5868 26188 5874 26200
rect 8202 26188 8208 26200
rect 8260 26188 8266 26240
rect 9766 26188 9772 26240
rect 9824 26228 9830 26240
rect 11793 26231 11851 26237
rect 11793 26228 11805 26231
rect 9824 26200 11805 26228
rect 9824 26188 9830 26200
rect 11793 26197 11805 26200
rect 11839 26197 11851 26231
rect 11793 26191 11851 26197
rect 14274 26188 14280 26240
rect 14332 26228 14338 26240
rect 14936 26228 14964 26268
rect 15654 26256 15660 26308
rect 15712 26256 15718 26308
rect 15749 26299 15807 26305
rect 15749 26265 15761 26299
rect 15795 26296 15807 26299
rect 16408 26296 16436 26324
rect 15795 26268 16436 26296
rect 16485 26299 16543 26305
rect 15795 26265 15807 26268
rect 15749 26259 15807 26265
rect 16485 26265 16497 26299
rect 16531 26265 16543 26299
rect 16485 26259 16543 26265
rect 14332 26200 14964 26228
rect 14332 26188 14338 26200
rect 15378 26188 15384 26240
rect 15436 26188 15442 26240
rect 15470 26188 15476 26240
rect 15528 26228 15534 26240
rect 15764 26228 15792 26259
rect 15528 26200 15792 26228
rect 15528 26188 15534 26200
rect 16206 26188 16212 26240
rect 16264 26228 16270 26240
rect 16500 26228 16528 26259
rect 16850 26256 16856 26308
rect 16908 26256 16914 26308
rect 17037 26299 17095 26305
rect 17037 26265 17049 26299
rect 17083 26265 17095 26299
rect 17037 26259 17095 26265
rect 16264 26200 16528 26228
rect 16264 26188 16270 26200
rect 16758 26188 16764 26240
rect 16816 26188 16822 26240
rect 17052 26228 17080 26259
rect 17126 26256 17132 26308
rect 17184 26256 17190 26308
rect 17788 26296 17816 26327
rect 18046 26324 18052 26336
rect 18104 26324 18110 26376
rect 18138 26324 18144 26376
rect 18196 26324 18202 26376
rect 18230 26324 18236 26376
rect 18288 26364 18294 26376
rect 18708 26373 18736 26472
rect 20533 26469 20545 26472
rect 20579 26500 20591 26503
rect 24596 26500 24624 26531
rect 24670 26528 24676 26580
rect 24728 26568 24734 26580
rect 24949 26571 25007 26577
rect 24949 26568 24961 26571
rect 24728 26540 24961 26568
rect 24728 26528 24734 26540
rect 24949 26537 24961 26540
rect 24995 26537 25007 26571
rect 24949 26531 25007 26537
rect 20579 26472 24624 26500
rect 20579 26469 20591 26472
rect 20533 26463 20591 26469
rect 18785 26435 18843 26441
rect 18785 26401 18797 26435
rect 18831 26432 18843 26435
rect 20438 26432 20444 26444
rect 18831 26404 20444 26432
rect 18831 26401 18843 26404
rect 18785 26395 18843 26401
rect 20438 26392 20444 26404
rect 20496 26432 20502 26444
rect 20625 26435 20683 26441
rect 20625 26432 20637 26435
rect 20496 26404 20637 26432
rect 20496 26392 20502 26404
rect 20625 26401 20637 26404
rect 20671 26401 20683 26435
rect 20625 26395 20683 26401
rect 20717 26435 20775 26441
rect 20717 26401 20729 26435
rect 20763 26432 20775 26435
rect 21177 26435 21235 26441
rect 21177 26432 21189 26435
rect 20763 26404 21189 26432
rect 20763 26401 20775 26404
rect 20717 26395 20775 26401
rect 21177 26401 21189 26404
rect 21223 26401 21235 26435
rect 21177 26395 21235 26401
rect 22281 26435 22339 26441
rect 22281 26401 22293 26435
rect 22327 26432 22339 26435
rect 22649 26435 22707 26441
rect 22649 26432 22661 26435
rect 22327 26404 22661 26432
rect 22327 26401 22339 26404
rect 22281 26395 22339 26401
rect 22649 26401 22661 26404
rect 22695 26401 22707 26435
rect 22649 26395 22707 26401
rect 22741 26435 22799 26441
rect 22741 26401 22753 26435
rect 22787 26432 22799 26435
rect 22830 26432 22836 26444
rect 22787 26404 22836 26432
rect 22787 26401 22799 26404
rect 22741 26395 22799 26401
rect 22830 26392 22836 26404
rect 22888 26392 22894 26444
rect 24688 26432 24716 26528
rect 24964 26500 24992 26531
rect 25038 26528 25044 26580
rect 25096 26568 25102 26580
rect 25409 26571 25467 26577
rect 25409 26568 25421 26571
rect 25096 26540 25421 26568
rect 25096 26528 25102 26540
rect 25409 26537 25421 26540
rect 25455 26537 25467 26571
rect 25409 26531 25467 26537
rect 25685 26571 25743 26577
rect 25685 26537 25697 26571
rect 25731 26568 25743 26571
rect 25866 26568 25872 26580
rect 25731 26540 25872 26568
rect 25731 26537 25743 26540
rect 25685 26531 25743 26537
rect 25130 26500 25136 26512
rect 24964 26472 25136 26500
rect 25130 26460 25136 26472
rect 25188 26460 25194 26512
rect 25222 26460 25228 26512
rect 25280 26460 25286 26512
rect 25498 26460 25504 26512
rect 25556 26460 25562 26512
rect 25700 26500 25728 26531
rect 25866 26528 25872 26540
rect 25924 26528 25930 26580
rect 26786 26528 26792 26580
rect 26844 26528 26850 26580
rect 28445 26571 28503 26577
rect 28445 26568 28457 26571
rect 27540 26540 28457 26568
rect 25684 26472 25728 26500
rect 22940 26404 24716 26432
rect 25240 26432 25268 26460
rect 25684 26432 25712 26472
rect 25240 26404 25712 26432
rect 18693 26367 18751 26373
rect 18693 26364 18705 26367
rect 18288 26336 18705 26364
rect 18288 26324 18294 26336
rect 18693 26333 18705 26336
rect 18739 26333 18751 26367
rect 18693 26327 18751 26333
rect 18969 26367 19027 26373
rect 18969 26333 18981 26367
rect 19015 26364 19027 26367
rect 19334 26364 19340 26376
rect 19015 26336 19340 26364
rect 19015 26333 19027 26336
rect 18969 26327 19027 26333
rect 19334 26324 19340 26336
rect 19392 26364 19398 26376
rect 20346 26364 20352 26376
rect 19392 26336 20352 26364
rect 19392 26324 19398 26336
rect 20346 26324 20352 26336
rect 20404 26364 20410 26376
rect 20809 26367 20867 26373
rect 20809 26364 20821 26367
rect 20404 26336 20821 26364
rect 20404 26324 20410 26336
rect 20809 26333 20821 26336
rect 20855 26333 20867 26367
rect 20809 26327 20867 26333
rect 20993 26367 21051 26373
rect 20993 26333 21005 26367
rect 21039 26333 21051 26367
rect 20993 26327 21051 26333
rect 21269 26367 21327 26373
rect 21269 26333 21281 26367
rect 21315 26364 21327 26367
rect 21358 26364 21364 26376
rect 21315 26336 21364 26364
rect 21315 26333 21327 26336
rect 21269 26327 21327 26333
rect 17235 26268 17816 26296
rect 17235 26228 17263 26268
rect 17862 26256 17868 26308
rect 17920 26256 17926 26308
rect 17957 26299 18015 26305
rect 17957 26265 17969 26299
rect 18003 26296 18015 26299
rect 19061 26299 19119 26305
rect 18003 26268 18736 26296
rect 18003 26265 18015 26268
rect 17957 26259 18015 26265
rect 18708 26240 18736 26268
rect 19061 26265 19073 26299
rect 19107 26296 19119 26299
rect 21008 26296 21036 26327
rect 21358 26324 21364 26336
rect 21416 26324 21422 26376
rect 22186 26324 22192 26376
rect 22244 26324 22250 26376
rect 22370 26324 22376 26376
rect 22428 26324 22434 26376
rect 22940 26296 22968 26404
rect 26694 26392 26700 26444
rect 26752 26392 26758 26444
rect 23109 26367 23167 26373
rect 23109 26333 23121 26367
rect 23155 26364 23167 26367
rect 23155 26336 23525 26364
rect 23155 26333 23167 26336
rect 23109 26327 23167 26333
rect 19107 26268 22968 26296
rect 23017 26299 23075 26305
rect 19107 26265 19119 26268
rect 19061 26259 19119 26265
rect 17052 26200 17263 26228
rect 17310 26188 17316 26240
rect 17368 26228 17374 26240
rect 17589 26231 17647 26237
rect 17589 26228 17601 26231
rect 17368 26200 17601 26228
rect 17368 26188 17374 26200
rect 17589 26197 17601 26200
rect 17635 26197 17647 26231
rect 17589 26191 17647 26197
rect 18690 26188 18696 26240
rect 18748 26188 18754 26240
rect 20806 26188 20812 26240
rect 20864 26228 20870 26240
rect 21008 26228 21036 26268
rect 23017 26265 23029 26299
rect 23063 26296 23075 26299
rect 23382 26296 23388 26308
rect 23063 26268 23388 26296
rect 23063 26265 23075 26268
rect 23017 26259 23075 26265
rect 23382 26256 23388 26268
rect 23440 26256 23446 26308
rect 23497 26296 23525 26336
rect 23566 26324 23572 26376
rect 23624 26324 23630 26376
rect 23661 26367 23719 26373
rect 23661 26333 23673 26367
rect 23707 26364 23719 26367
rect 24210 26364 24216 26376
rect 23707 26336 24216 26364
rect 23707 26333 23719 26336
rect 23661 26327 23719 26333
rect 24210 26324 24216 26336
rect 24268 26324 24274 26376
rect 24486 26324 24492 26376
rect 24544 26364 24550 26376
rect 24581 26367 24639 26373
rect 24581 26364 24593 26367
rect 24544 26336 24593 26364
rect 24544 26324 24550 26336
rect 24581 26333 24593 26336
rect 24627 26333 24639 26367
rect 24581 26327 24639 26333
rect 24670 26324 24676 26376
rect 24728 26324 24734 26376
rect 24762 26324 24768 26376
rect 24820 26364 24826 26376
rect 25133 26367 25191 26373
rect 25133 26364 25145 26367
rect 24820 26336 25145 26364
rect 24820 26324 24826 26336
rect 25133 26333 25145 26336
rect 25179 26333 25191 26367
rect 25133 26327 25191 26333
rect 25225 26367 25283 26373
rect 25225 26333 25237 26367
rect 25271 26364 25283 26367
rect 25498 26364 25504 26376
rect 25271 26336 25504 26364
rect 25271 26333 25283 26336
rect 25225 26327 25283 26333
rect 25498 26324 25504 26336
rect 25556 26324 25562 26376
rect 26881 26367 26939 26373
rect 26881 26333 26893 26367
rect 26927 26333 26939 26367
rect 26881 26327 26939 26333
rect 26973 26367 27031 26373
rect 26973 26333 26985 26367
rect 27019 26364 27031 26367
rect 27062 26364 27068 26376
rect 27019 26336 27068 26364
rect 27019 26333 27031 26336
rect 26973 26327 27031 26333
rect 24857 26299 24915 26305
rect 23497 26268 24624 26296
rect 24596 26240 24624 26268
rect 24857 26265 24869 26299
rect 24903 26296 24915 26299
rect 24949 26299 25007 26305
rect 24949 26296 24961 26299
rect 24903 26268 24961 26296
rect 24903 26265 24915 26268
rect 24857 26259 24915 26265
rect 24949 26265 24961 26268
rect 24995 26296 25007 26299
rect 25038 26296 25044 26308
rect 24995 26268 25044 26296
rect 24995 26265 25007 26268
rect 24949 26259 25007 26265
rect 25038 26256 25044 26268
rect 25096 26256 25102 26308
rect 25682 26305 25688 26308
rect 25669 26299 25688 26305
rect 25669 26265 25681 26299
rect 25669 26259 25688 26265
rect 25682 26256 25688 26259
rect 25740 26256 25746 26308
rect 25869 26299 25927 26305
rect 25869 26265 25881 26299
rect 25915 26296 25927 26299
rect 26050 26296 26056 26308
rect 25915 26268 26056 26296
rect 25915 26265 25927 26268
rect 25869 26259 25927 26265
rect 26050 26256 26056 26268
rect 26108 26256 26114 26308
rect 26896 26296 26924 26327
rect 27062 26324 27068 26336
rect 27120 26364 27126 26376
rect 27540 26364 27568 26540
rect 28445 26537 28457 26540
rect 28491 26537 28503 26571
rect 28445 26531 28503 26537
rect 29730 26528 29736 26580
rect 29788 26528 29794 26580
rect 31481 26571 31539 26577
rect 31481 26537 31493 26571
rect 31527 26568 31539 26571
rect 31754 26568 31760 26580
rect 31527 26540 31760 26568
rect 31527 26537 31539 26540
rect 31481 26531 31539 26537
rect 27982 26460 27988 26512
rect 28040 26460 28046 26512
rect 28534 26460 28540 26512
rect 28592 26500 28598 26512
rect 28997 26503 29055 26509
rect 28997 26500 29009 26503
rect 28592 26472 29009 26500
rect 28592 26460 28598 26472
rect 28997 26469 29009 26472
rect 29043 26469 29055 26503
rect 28997 26463 29055 26469
rect 27614 26392 27620 26444
rect 27672 26392 27678 26444
rect 28000 26432 28028 26460
rect 28077 26435 28135 26441
rect 28077 26432 28089 26435
rect 28000 26404 28089 26432
rect 28077 26401 28089 26404
rect 28123 26401 28135 26435
rect 28077 26395 28135 26401
rect 28166 26392 28172 26444
rect 28224 26432 28230 26444
rect 28721 26435 28779 26441
rect 28721 26432 28733 26435
rect 28224 26404 28733 26432
rect 28224 26392 28230 26404
rect 28721 26401 28733 26404
rect 28767 26401 28779 26435
rect 28721 26395 28779 26401
rect 29270 26392 29276 26444
rect 29328 26432 29334 26444
rect 29748 26432 29776 26528
rect 31496 26500 31524 26531
rect 31754 26528 31760 26540
rect 31812 26528 31818 26580
rect 34514 26528 34520 26580
rect 34572 26528 34578 26580
rect 34977 26571 35035 26577
rect 34624 26540 34928 26568
rect 29328 26404 29776 26432
rect 31220 26472 31524 26500
rect 32401 26503 32459 26509
rect 29328 26392 29334 26404
rect 27120 26336 27568 26364
rect 27120 26324 27126 26336
rect 27706 26324 27712 26376
rect 27764 26324 27770 26376
rect 27798 26324 27804 26376
rect 27856 26324 27862 26376
rect 27890 26324 27896 26376
rect 27948 26324 27954 26376
rect 27982 26324 27988 26376
rect 28040 26324 28046 26376
rect 28261 26367 28319 26373
rect 28261 26333 28273 26367
rect 28307 26364 28319 26367
rect 28307 26336 28396 26364
rect 28307 26333 28319 26336
rect 28261 26327 28319 26333
rect 27724 26296 27752 26324
rect 26896 26268 27752 26296
rect 20864 26200 21036 26228
rect 20864 26188 20870 26200
rect 22830 26188 22836 26240
rect 22888 26188 22894 26240
rect 23106 26188 23112 26240
rect 23164 26228 23170 26240
rect 23293 26231 23351 26237
rect 23293 26228 23305 26231
rect 23164 26200 23305 26228
rect 23164 26188 23170 26200
rect 23293 26197 23305 26200
rect 23339 26197 23351 26231
rect 23293 26191 23351 26197
rect 24026 26188 24032 26240
rect 24084 26228 24090 26240
rect 24394 26228 24400 26240
rect 24084 26200 24400 26228
rect 24084 26188 24090 26200
rect 24394 26188 24400 26200
rect 24452 26188 24458 26240
rect 24578 26188 24584 26240
rect 24636 26188 24642 26240
rect 28258 26188 28264 26240
rect 28316 26228 28322 26240
rect 28368 26228 28396 26336
rect 28442 26324 28448 26376
rect 28500 26324 28506 26376
rect 28810 26324 28816 26376
rect 28868 26324 28874 26376
rect 29914 26324 29920 26376
rect 29972 26324 29978 26376
rect 30742 26324 30748 26376
rect 30800 26364 30806 26376
rect 31113 26367 31171 26373
rect 31113 26364 31125 26367
rect 30800 26336 31125 26364
rect 30800 26324 30806 26336
rect 31113 26333 31125 26336
rect 31159 26333 31171 26367
rect 31220 26364 31248 26472
rect 32401 26469 32413 26503
rect 32447 26500 32459 26503
rect 32490 26500 32496 26512
rect 32447 26472 32496 26500
rect 32447 26469 32459 26472
rect 32401 26463 32459 26469
rect 32490 26460 32496 26472
rect 32548 26460 32554 26512
rect 33594 26460 33600 26512
rect 33652 26500 33658 26512
rect 33870 26500 33876 26512
rect 33652 26472 33876 26500
rect 33652 26460 33658 26472
rect 33870 26460 33876 26472
rect 33928 26460 33934 26512
rect 31938 26392 31944 26444
rect 31996 26432 32002 26444
rect 34624 26432 34652 26540
rect 34701 26503 34759 26509
rect 34701 26469 34713 26503
rect 34747 26469 34759 26503
rect 34701 26463 34759 26469
rect 31996 26404 34652 26432
rect 31996 26392 32002 26404
rect 31297 26367 31355 26373
rect 31297 26364 31309 26367
rect 31220 26336 31309 26364
rect 31113 26327 31171 26333
rect 31297 26333 31309 26336
rect 31343 26333 31355 26367
rect 31297 26327 31355 26333
rect 31386 26324 31392 26376
rect 31444 26324 31450 26376
rect 31570 26324 31576 26376
rect 31628 26364 31634 26376
rect 31665 26367 31723 26373
rect 31665 26364 31677 26367
rect 31628 26336 31677 26364
rect 31628 26324 31634 26336
rect 31665 26333 31677 26336
rect 31711 26333 31723 26367
rect 31665 26327 31723 26333
rect 31846 26324 31852 26376
rect 31904 26324 31910 26376
rect 32030 26324 32036 26376
rect 32088 26364 32094 26376
rect 32309 26367 32367 26373
rect 32309 26364 32321 26367
rect 32088 26336 32321 26364
rect 32088 26324 32094 26336
rect 32309 26333 32321 26336
rect 32355 26364 32367 26367
rect 32398 26364 32404 26376
rect 32355 26336 32404 26364
rect 32355 26333 32367 26336
rect 32309 26327 32367 26333
rect 32398 26324 32404 26336
rect 32456 26324 32462 26376
rect 32490 26324 32496 26376
rect 32548 26324 32554 26376
rect 32582 26324 32588 26376
rect 32640 26324 32646 26376
rect 33502 26324 33508 26376
rect 33560 26364 33566 26376
rect 33870 26364 33876 26376
rect 33560 26336 33876 26364
rect 33560 26324 33566 26336
rect 33870 26324 33876 26336
rect 33928 26364 33934 26376
rect 34333 26367 34391 26373
rect 34333 26364 34345 26367
rect 33928 26336 34345 26364
rect 33928 26324 33934 26336
rect 34333 26333 34345 26336
rect 34379 26333 34391 26367
rect 34333 26327 34391 26333
rect 34422 26324 34428 26376
rect 34480 26364 34486 26376
rect 34517 26367 34575 26373
rect 34517 26364 34529 26367
rect 34480 26336 34529 26364
rect 34480 26324 34486 26336
rect 34517 26333 34529 26336
rect 34563 26364 34575 26367
rect 34716 26364 34744 26463
rect 34900 26373 34928 26540
rect 34977 26537 34989 26571
rect 35023 26568 35035 26571
rect 35023 26540 36308 26568
rect 35023 26537 35035 26540
rect 34977 26531 35035 26537
rect 35342 26460 35348 26512
rect 35400 26460 35406 26512
rect 36280 26500 36308 26540
rect 36354 26528 36360 26580
rect 36412 26568 36418 26580
rect 38378 26568 38384 26580
rect 36412 26540 38384 26568
rect 36412 26528 36418 26540
rect 38378 26528 38384 26540
rect 38436 26568 38442 26580
rect 40037 26571 40095 26577
rect 40037 26568 40049 26571
rect 38436 26540 40049 26568
rect 38436 26528 38442 26540
rect 40037 26537 40049 26540
rect 40083 26537 40095 26571
rect 40037 26531 40095 26537
rect 37550 26500 37556 26512
rect 36280 26472 37556 26500
rect 37550 26460 37556 26472
rect 37608 26500 37614 26512
rect 37737 26503 37795 26509
rect 37737 26500 37749 26503
rect 37608 26472 37749 26500
rect 37608 26460 37614 26472
rect 37737 26469 37749 26472
rect 37783 26500 37795 26503
rect 38470 26500 38476 26512
rect 37783 26472 38476 26500
rect 37783 26469 37795 26472
rect 37737 26463 37795 26469
rect 38470 26460 38476 26472
rect 38528 26460 38534 26512
rect 38930 26460 38936 26512
rect 38988 26500 38994 26512
rect 39298 26500 39304 26512
rect 38988 26472 39304 26500
rect 38988 26460 38994 26472
rect 39298 26460 39304 26472
rect 39356 26460 39362 26512
rect 35360 26432 35388 26460
rect 37090 26432 37096 26444
rect 35268 26404 37096 26432
rect 35268 26373 35296 26404
rect 37090 26392 37096 26404
rect 37148 26392 37154 26444
rect 37274 26392 37280 26444
rect 37332 26432 37338 26444
rect 38013 26435 38071 26441
rect 38013 26432 38025 26435
rect 37332 26404 38025 26432
rect 37332 26392 37338 26404
rect 38013 26401 38025 26404
rect 38059 26401 38071 26435
rect 38013 26395 38071 26401
rect 38102 26392 38108 26444
rect 38160 26392 38166 26444
rect 34563 26336 34744 26364
rect 34885 26367 34943 26373
rect 34563 26333 34575 26336
rect 34517 26327 34575 26333
rect 34885 26333 34897 26367
rect 34931 26333 34943 26367
rect 34885 26327 34943 26333
rect 35253 26367 35311 26373
rect 35253 26333 35265 26367
rect 35299 26333 35311 26367
rect 35253 26327 35311 26333
rect 35345 26367 35403 26373
rect 35345 26333 35357 26367
rect 35391 26333 35403 26367
rect 35345 26327 35403 26333
rect 28626 26256 28632 26308
rect 28684 26296 28690 26308
rect 29730 26296 29736 26308
rect 28684 26268 29736 26296
rect 28684 26256 28690 26268
rect 29730 26256 29736 26268
rect 29788 26256 29794 26308
rect 31202 26256 31208 26308
rect 31260 26256 31266 26308
rect 32508 26296 32536 26324
rect 31726 26268 32536 26296
rect 28316 26200 28396 26228
rect 28316 26188 28322 26200
rect 31110 26188 31116 26240
rect 31168 26228 31174 26240
rect 31726 26228 31754 26268
rect 32766 26256 32772 26308
rect 32824 26296 32830 26308
rect 35360 26296 35388 26327
rect 35526 26324 35532 26376
rect 35584 26364 35590 26376
rect 37734 26364 37740 26376
rect 35584 26336 37740 26364
rect 35584 26324 35590 26336
rect 37734 26324 37740 26336
rect 37792 26324 37798 26376
rect 37826 26324 37832 26376
rect 37884 26364 37890 26376
rect 37921 26367 37979 26373
rect 37921 26364 37933 26367
rect 37884 26336 37933 26364
rect 37884 26324 37890 26336
rect 37921 26333 37933 26336
rect 37967 26333 37979 26367
rect 39758 26364 39764 26376
rect 37921 26327 37979 26333
rect 38028 26336 39764 26364
rect 32824 26268 35388 26296
rect 32824 26256 32830 26268
rect 35618 26256 35624 26308
rect 35676 26256 35682 26308
rect 35986 26256 35992 26308
rect 36044 26296 36050 26308
rect 38028 26296 38056 26336
rect 39758 26324 39764 26336
rect 39816 26324 39822 26376
rect 39942 26324 39948 26376
rect 40000 26364 40006 26376
rect 40221 26367 40279 26373
rect 40221 26364 40233 26367
rect 40000 26336 40233 26364
rect 40000 26324 40006 26336
rect 40221 26333 40233 26336
rect 40267 26333 40279 26367
rect 40221 26327 40279 26333
rect 36044 26268 38056 26296
rect 36044 26256 36050 26268
rect 38378 26256 38384 26308
rect 38436 26256 38442 26308
rect 31168 26200 31754 26228
rect 31168 26188 31174 26200
rect 31846 26188 31852 26240
rect 31904 26188 31910 26240
rect 33134 26188 33140 26240
rect 33192 26228 33198 26240
rect 34882 26228 34888 26240
rect 33192 26200 34888 26228
rect 33192 26188 33198 26200
rect 34882 26188 34888 26200
rect 34940 26188 34946 26240
rect 35066 26188 35072 26240
rect 35124 26228 35130 26240
rect 35713 26231 35771 26237
rect 35713 26228 35725 26231
rect 35124 26200 35725 26228
rect 35124 26188 35130 26200
rect 35713 26197 35725 26200
rect 35759 26228 35771 26231
rect 36538 26228 36544 26240
rect 35759 26200 36544 26228
rect 35759 26197 35771 26200
rect 35713 26191 35771 26197
rect 36538 26188 36544 26200
rect 36596 26188 36602 26240
rect 1104 26138 40572 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 40572 26138
rect 1104 26064 40572 26086
rect 3329 26027 3387 26033
rect 3329 25993 3341 26027
rect 3375 26024 3387 26027
rect 4338 26024 4344 26036
rect 3375 25996 4344 26024
rect 3375 25993 3387 25996
rect 3329 25987 3387 25993
rect 4338 25984 4344 25996
rect 4396 26024 4402 26036
rect 5350 26024 5356 26036
rect 4396 25996 5356 26024
rect 4396 25984 4402 25996
rect 5350 25984 5356 25996
rect 5408 25984 5414 26036
rect 5445 26027 5503 26033
rect 5445 25993 5457 26027
rect 5491 26024 5503 26027
rect 5626 26024 5632 26036
rect 5491 25996 5632 26024
rect 5491 25993 5503 25996
rect 5445 25987 5503 25993
rect 5626 25984 5632 25996
rect 5684 25984 5690 26036
rect 7098 25984 7104 26036
rect 7156 26024 7162 26036
rect 7745 26027 7803 26033
rect 7745 26024 7757 26027
rect 7156 25996 7757 26024
rect 7156 25984 7162 25996
rect 7745 25993 7757 25996
rect 7791 25993 7803 26027
rect 7745 25987 7803 25993
rect 9214 25984 9220 26036
rect 9272 26024 9278 26036
rect 10137 26027 10195 26033
rect 10137 26024 10149 26027
rect 9272 25996 10149 26024
rect 9272 25984 9278 25996
rect 10137 25993 10149 25996
rect 10183 25993 10195 26027
rect 10137 25987 10195 25993
rect 11882 25984 11888 26036
rect 11940 26024 11946 26036
rect 12250 26024 12256 26036
rect 11940 25996 12256 26024
rect 11940 25984 11946 25996
rect 12250 25984 12256 25996
rect 12308 25984 12314 26036
rect 16758 26024 16764 26036
rect 12406 25996 16764 26024
rect 1854 25916 1860 25968
rect 1912 25916 1918 25968
rect 3142 25956 3148 25968
rect 3082 25928 3148 25956
rect 3142 25916 3148 25928
rect 3200 25956 3206 25968
rect 3970 25956 3976 25968
rect 3200 25928 3976 25956
rect 3200 25916 3206 25928
rect 3970 25916 3976 25928
rect 4028 25956 4034 25968
rect 4430 25956 4436 25968
rect 4028 25928 4436 25956
rect 4028 25916 4034 25928
rect 4430 25916 4436 25928
rect 4488 25916 4494 25968
rect 3694 25848 3700 25900
rect 3752 25848 3758 25900
rect 5644 25888 5672 25984
rect 6270 25916 6276 25968
rect 6328 25956 6334 25968
rect 6641 25959 6699 25965
rect 6641 25956 6653 25959
rect 6328 25928 6653 25956
rect 6328 25916 6334 25928
rect 6641 25925 6653 25928
rect 6687 25956 6699 25959
rect 7377 25959 7435 25965
rect 7377 25956 7389 25959
rect 6687 25928 7389 25956
rect 6687 25925 6699 25928
rect 6641 25919 6699 25925
rect 7377 25925 7389 25928
rect 7423 25925 7435 25959
rect 7377 25919 7435 25925
rect 10321 25959 10379 25965
rect 10321 25925 10333 25959
rect 10367 25956 10379 25959
rect 12406 25956 12434 25996
rect 16758 25984 16764 25996
rect 16816 25984 16822 26036
rect 18417 26027 18475 26033
rect 18417 25993 18429 26027
rect 18463 26024 18475 26027
rect 18874 26024 18880 26036
rect 18463 25996 18880 26024
rect 18463 25993 18475 25996
rect 18417 25987 18475 25993
rect 18874 25984 18880 25996
rect 18932 25984 18938 26036
rect 24210 25984 24216 26036
rect 24268 26024 24274 26036
rect 25590 26024 25596 26036
rect 24268 25996 25596 26024
rect 24268 25984 24274 25996
rect 25590 25984 25596 25996
rect 25648 25984 25654 26036
rect 25774 25984 25780 26036
rect 25832 26024 25838 26036
rect 26053 26027 26111 26033
rect 26053 26024 26065 26027
rect 25832 25996 26065 26024
rect 25832 25984 25838 25996
rect 26053 25993 26065 25996
rect 26099 25993 26111 26027
rect 26053 25987 26111 25993
rect 28258 25984 28264 26036
rect 28316 26024 28322 26036
rect 28353 26027 28411 26033
rect 28353 26024 28365 26027
rect 28316 25996 28365 26024
rect 28316 25984 28322 25996
rect 28353 25993 28365 25996
rect 28399 25993 28411 26027
rect 28353 25987 28411 25993
rect 29362 25984 29368 26036
rect 29420 26024 29426 26036
rect 29457 26027 29515 26033
rect 29457 26024 29469 26027
rect 29420 25996 29469 26024
rect 29420 25984 29426 25996
rect 29457 25993 29469 25996
rect 29503 25993 29515 26027
rect 29457 25987 29515 25993
rect 30561 26027 30619 26033
rect 30561 25993 30573 26027
rect 30607 26024 30619 26027
rect 30834 26024 30840 26036
rect 30607 25996 30840 26024
rect 30607 25993 30619 25996
rect 30561 25987 30619 25993
rect 30834 25984 30840 25996
rect 30892 25984 30898 26036
rect 33962 26024 33968 26036
rect 30944 25996 33968 26024
rect 10367 25928 12434 25956
rect 12621 25959 12679 25965
rect 10367 25925 10379 25928
rect 10321 25919 10379 25925
rect 12621 25925 12633 25959
rect 12667 25956 12679 25959
rect 15378 25956 15384 25968
rect 12667 25928 15384 25956
rect 12667 25925 12679 25928
rect 12621 25919 12679 25925
rect 6089 25891 6147 25897
rect 6089 25888 6101 25891
rect 5644 25860 6101 25888
rect 6089 25857 6101 25860
rect 6135 25857 6147 25891
rect 6089 25851 6147 25857
rect 6362 25848 6368 25900
rect 6420 25848 6426 25900
rect 6546 25897 6552 25900
rect 6513 25891 6552 25897
rect 6513 25857 6525 25891
rect 6513 25851 6552 25857
rect 6546 25848 6552 25851
rect 6604 25848 6610 25900
rect 1578 25780 1584 25832
rect 1636 25780 1642 25832
rect 3970 25780 3976 25832
rect 4028 25780 4034 25832
rect 6546 25712 6552 25764
rect 6604 25752 6610 25764
rect 6656 25752 6684 25919
rect 15378 25916 15384 25928
rect 15436 25916 15442 25968
rect 19245 25959 19303 25965
rect 18708 25928 19196 25956
rect 6733 25891 6791 25897
rect 6733 25857 6745 25891
rect 6779 25857 6791 25891
rect 6733 25851 6791 25857
rect 6604 25724 6684 25752
rect 6748 25752 6776 25851
rect 6822 25848 6828 25900
rect 6880 25897 6886 25900
rect 6880 25891 6929 25897
rect 6880 25857 6883 25891
rect 6917 25857 6929 25891
rect 6880 25851 6929 25857
rect 6880 25848 6914 25851
rect 7006 25848 7012 25900
rect 7064 25888 7070 25900
rect 7101 25891 7159 25897
rect 7101 25888 7113 25891
rect 7064 25860 7113 25888
rect 7064 25848 7070 25860
rect 7101 25857 7113 25860
rect 7147 25857 7159 25891
rect 7101 25851 7159 25857
rect 7190 25848 7196 25900
rect 7248 25848 7254 25900
rect 7466 25848 7472 25900
rect 7524 25848 7530 25900
rect 7607 25891 7665 25897
rect 7607 25857 7619 25891
rect 7653 25888 7665 25891
rect 8478 25888 8484 25900
rect 7653 25860 8484 25888
rect 7653 25857 7665 25860
rect 7607 25851 7665 25857
rect 6886 25820 6914 25848
rect 7622 25820 7650 25851
rect 8478 25848 8484 25860
rect 8536 25848 8542 25900
rect 10042 25848 10048 25900
rect 10100 25848 10106 25900
rect 11517 25891 11575 25897
rect 11517 25857 11529 25891
rect 11563 25857 11575 25891
rect 11517 25851 11575 25857
rect 6886 25792 7650 25820
rect 11532 25820 11560 25851
rect 11698 25848 11704 25900
rect 11756 25848 11762 25900
rect 11882 25848 11888 25900
rect 11940 25848 11946 25900
rect 11974 25848 11980 25900
rect 12032 25888 12038 25900
rect 12345 25891 12403 25897
rect 12345 25888 12357 25891
rect 12032 25860 12357 25888
rect 12032 25848 12038 25860
rect 12345 25857 12357 25860
rect 12391 25857 12403 25891
rect 12345 25851 12403 25857
rect 12434 25848 12440 25900
rect 12492 25888 12498 25900
rect 13078 25888 13084 25900
rect 12492 25860 13084 25888
rect 12492 25848 12498 25860
rect 13078 25848 13084 25860
rect 13136 25848 13142 25900
rect 13354 25848 13360 25900
rect 13412 25848 13418 25900
rect 13541 25891 13599 25897
rect 13541 25857 13553 25891
rect 13587 25857 13599 25891
rect 13541 25851 13599 25857
rect 12526 25820 12532 25832
rect 11532 25792 12532 25820
rect 12526 25780 12532 25792
rect 12584 25820 12590 25832
rect 13372 25820 13400 25848
rect 12584 25792 13400 25820
rect 13556 25820 13584 25851
rect 13630 25848 13636 25900
rect 13688 25848 13694 25900
rect 13814 25848 13820 25900
rect 13872 25848 13878 25900
rect 13906 25848 13912 25900
rect 13964 25848 13970 25900
rect 13998 25848 14004 25900
rect 14056 25848 14062 25900
rect 14090 25848 14096 25900
rect 14148 25888 14154 25900
rect 14461 25891 14519 25897
rect 14461 25888 14473 25891
rect 14148 25860 14473 25888
rect 14148 25848 14154 25860
rect 14461 25857 14473 25860
rect 14507 25857 14519 25891
rect 14461 25851 14519 25857
rect 14550 25848 14556 25900
rect 14608 25848 14614 25900
rect 14737 25891 14795 25897
rect 14737 25857 14749 25891
rect 14783 25888 14795 25891
rect 14918 25888 14924 25900
rect 14783 25860 14924 25888
rect 14783 25857 14795 25860
rect 14737 25851 14795 25857
rect 14918 25848 14924 25860
rect 14976 25848 14982 25900
rect 18141 25891 18199 25897
rect 18141 25857 18153 25891
rect 18187 25888 18199 25891
rect 18230 25888 18236 25900
rect 18187 25860 18236 25888
rect 18187 25857 18199 25860
rect 18141 25851 18199 25857
rect 18230 25848 18236 25860
rect 18288 25848 18294 25900
rect 18322 25848 18328 25900
rect 18380 25888 18386 25900
rect 18417 25891 18475 25897
rect 18417 25888 18429 25891
rect 18380 25860 18429 25888
rect 18380 25848 18386 25860
rect 18417 25857 18429 25860
rect 18463 25888 18475 25891
rect 18708 25888 18736 25928
rect 18463 25860 18736 25888
rect 18463 25857 18475 25860
rect 18417 25851 18475 25857
rect 19058 25848 19064 25900
rect 19116 25848 19122 25900
rect 19168 25888 19196 25928
rect 19245 25925 19257 25959
rect 19291 25956 19303 25959
rect 19334 25956 19340 25968
rect 19291 25928 19340 25956
rect 19291 25925 19303 25928
rect 19245 25919 19303 25925
rect 19334 25916 19340 25928
rect 19392 25916 19398 25968
rect 25608 25956 25636 25984
rect 28534 25956 28540 25968
rect 25608 25928 28540 25956
rect 24670 25888 24676 25900
rect 19168 25860 24676 25888
rect 24670 25848 24676 25860
rect 24728 25848 24734 25900
rect 25961 25891 26019 25897
rect 25961 25857 25973 25891
rect 26007 25857 26019 25891
rect 25961 25851 26019 25857
rect 14277 25823 14335 25829
rect 14277 25820 14289 25823
rect 13556 25792 13860 25820
rect 12584 25780 12590 25792
rect 13722 25752 13728 25764
rect 6748 25724 13728 25752
rect 6604 25712 6610 25724
rect 13722 25712 13728 25724
rect 13780 25712 13786 25764
rect 13832 25752 13860 25792
rect 14108 25792 14289 25820
rect 14108 25752 14136 25792
rect 14277 25789 14289 25792
rect 14323 25789 14335 25823
rect 14277 25783 14335 25789
rect 14369 25823 14427 25829
rect 14369 25789 14381 25823
rect 14415 25789 14427 25823
rect 14369 25783 14427 25789
rect 13832 25724 14136 25752
rect 14185 25755 14243 25761
rect 14185 25721 14197 25755
rect 14231 25752 14243 25755
rect 14384 25752 14412 25783
rect 15102 25780 15108 25832
rect 15160 25820 15166 25832
rect 15473 25823 15531 25829
rect 15473 25820 15485 25823
rect 15160 25792 15485 25820
rect 15160 25780 15166 25792
rect 15473 25789 15485 25792
rect 15519 25789 15531 25823
rect 15473 25783 15531 25789
rect 15933 25823 15991 25829
rect 15933 25789 15945 25823
rect 15979 25820 15991 25823
rect 16022 25820 16028 25832
rect 15979 25792 16028 25820
rect 15979 25789 15991 25792
rect 15933 25783 15991 25789
rect 16022 25780 16028 25792
rect 16080 25780 16086 25832
rect 17678 25780 17684 25832
rect 17736 25820 17742 25832
rect 23198 25820 23204 25832
rect 17736 25792 23204 25820
rect 17736 25780 17742 25792
rect 23198 25780 23204 25792
rect 23256 25780 23262 25832
rect 25976 25820 26004 25851
rect 26050 25848 26056 25900
rect 26108 25888 26114 25900
rect 28460 25897 28488 25928
rect 28534 25916 28540 25928
rect 28592 25916 28598 25968
rect 29181 25959 29239 25965
rect 29181 25925 29193 25959
rect 29227 25956 29239 25959
rect 30377 25959 30435 25965
rect 30377 25956 30389 25959
rect 29227 25928 30389 25956
rect 29227 25925 29239 25928
rect 29181 25919 29239 25925
rect 29380 25900 29408 25928
rect 30377 25925 30389 25928
rect 30423 25925 30435 25959
rect 30944 25956 30972 25996
rect 33962 25984 33968 25996
rect 34020 25984 34026 26036
rect 36078 26024 36084 26036
rect 34624 25996 36084 26024
rect 30377 25919 30435 25925
rect 30852 25928 30972 25956
rect 26145 25891 26203 25897
rect 26145 25888 26157 25891
rect 26108 25860 26157 25888
rect 26108 25848 26114 25860
rect 26145 25857 26157 25860
rect 26191 25857 26203 25891
rect 26145 25851 26203 25857
rect 28445 25891 28503 25897
rect 28445 25857 28457 25891
rect 28491 25857 28503 25891
rect 28445 25851 28503 25857
rect 28997 25891 29055 25897
rect 28997 25857 29009 25891
rect 29043 25857 29055 25891
rect 28997 25851 29055 25857
rect 29012 25820 29040 25851
rect 29270 25848 29276 25900
rect 29328 25848 29334 25900
rect 29362 25848 29368 25900
rect 29420 25848 29426 25900
rect 29546 25848 29552 25900
rect 29604 25888 29610 25900
rect 29825 25891 29883 25897
rect 29825 25888 29837 25891
rect 29604 25860 29837 25888
rect 29604 25848 29610 25860
rect 29825 25857 29837 25860
rect 29871 25888 29883 25891
rect 30193 25891 30251 25897
rect 30193 25888 30205 25891
rect 29871 25860 30205 25888
rect 29871 25857 29883 25860
rect 29825 25851 29883 25857
rect 30193 25857 30205 25860
rect 30239 25888 30251 25891
rect 30852 25888 30880 25928
rect 31110 25916 31116 25968
rect 31168 25956 31174 25968
rect 31205 25959 31263 25965
rect 31205 25956 31217 25959
rect 31168 25928 31217 25956
rect 31168 25916 31174 25928
rect 31205 25925 31217 25928
rect 31251 25925 31263 25959
rect 31205 25919 31263 25925
rect 31294 25916 31300 25968
rect 31352 25916 31358 25968
rect 31386 25916 31392 25968
rect 31444 25956 31450 25968
rect 34624 25956 34652 25996
rect 34782 25965 34810 25996
rect 36078 25984 36084 25996
rect 36136 25984 36142 26036
rect 38010 25984 38016 26036
rect 38068 26024 38074 26036
rect 38105 26027 38163 26033
rect 38105 26024 38117 26027
rect 38068 25996 38117 26024
rect 38068 25984 38074 25996
rect 38105 25993 38117 25996
rect 38151 25993 38163 26027
rect 38105 25987 38163 25993
rect 31444 25928 34652 25956
rect 34767 25959 34825 25965
rect 31444 25916 31450 25928
rect 34767 25925 34779 25959
rect 34813 25925 34825 25959
rect 34767 25919 34825 25925
rect 34977 25959 35035 25965
rect 34977 25925 34989 25959
rect 35023 25956 35035 25959
rect 35342 25956 35348 25968
rect 35023 25928 35348 25956
rect 35023 25925 35035 25928
rect 34977 25919 35035 25925
rect 30239 25860 30880 25888
rect 30239 25857 30251 25860
rect 30193 25851 30251 25857
rect 30926 25848 30932 25900
rect 30984 25848 30990 25900
rect 31312 25888 31340 25916
rect 31570 25888 31576 25900
rect 31312 25860 31576 25888
rect 31570 25848 31576 25860
rect 31628 25888 31634 25900
rect 31665 25891 31723 25897
rect 31665 25888 31677 25891
rect 31628 25860 31677 25888
rect 31628 25848 31634 25860
rect 31665 25857 31677 25860
rect 31711 25857 31723 25891
rect 31665 25851 31723 25857
rect 32490 25848 32496 25900
rect 32548 25848 32554 25900
rect 33870 25848 33876 25900
rect 33928 25848 33934 25900
rect 34057 25891 34115 25897
rect 34057 25857 34069 25891
rect 34103 25888 34115 25891
rect 34149 25891 34207 25897
rect 34149 25888 34161 25891
rect 34103 25860 34161 25888
rect 34103 25857 34115 25860
rect 34057 25851 34115 25857
rect 34149 25857 34161 25860
rect 34195 25888 34207 25891
rect 34330 25888 34336 25900
rect 34195 25860 34336 25888
rect 34195 25857 34207 25860
rect 34149 25851 34207 25857
rect 29564 25820 29592 25848
rect 25976 25792 26188 25820
rect 29012 25792 29592 25820
rect 31297 25823 31355 25829
rect 26160 25764 26188 25792
rect 31297 25789 31309 25823
rect 31343 25820 31355 25823
rect 34072 25820 34100 25851
rect 34330 25848 34336 25860
rect 34388 25848 34394 25900
rect 34422 25848 34428 25900
rect 34480 25848 34486 25900
rect 34514 25848 34520 25900
rect 34572 25888 34578 25900
rect 34609 25891 34667 25897
rect 34609 25888 34621 25891
rect 34572 25860 34621 25888
rect 34572 25848 34578 25860
rect 34609 25857 34621 25860
rect 34655 25857 34667 25891
rect 34609 25851 34667 25857
rect 34882 25848 34888 25900
rect 34940 25848 34946 25900
rect 34992 25820 35020 25919
rect 35342 25916 35348 25928
rect 35400 25916 35406 25968
rect 36170 25916 36176 25968
rect 36228 25956 36234 25968
rect 36722 25956 36728 25968
rect 36228 25928 36728 25956
rect 36228 25916 36234 25928
rect 36722 25916 36728 25928
rect 36780 25916 36786 25968
rect 35066 25848 35072 25900
rect 35124 25848 35130 25900
rect 37642 25848 37648 25900
rect 37700 25888 37706 25900
rect 37988 25891 38046 25897
rect 37988 25888 38000 25891
rect 37700 25860 38000 25888
rect 37700 25848 37706 25860
rect 37988 25857 38000 25860
rect 38034 25888 38046 25891
rect 38034 25860 38332 25888
rect 38034 25857 38046 25860
rect 37988 25851 38046 25857
rect 31343 25792 34100 25820
rect 34128 25792 35020 25820
rect 31343 25789 31355 25792
rect 31297 25783 31355 25789
rect 14231 25724 14412 25752
rect 14231 25721 14243 25724
rect 14185 25715 14243 25721
rect 15194 25712 15200 25764
rect 15252 25752 15258 25764
rect 15565 25755 15623 25761
rect 15565 25752 15577 25755
rect 15252 25724 15577 25752
rect 15252 25712 15258 25724
rect 15565 25721 15577 25724
rect 15611 25721 15623 25755
rect 15565 25715 15623 25721
rect 18138 25712 18144 25764
rect 18196 25752 18202 25764
rect 18325 25755 18383 25761
rect 18325 25752 18337 25755
rect 18196 25724 18337 25752
rect 18196 25712 18202 25724
rect 18325 25721 18337 25724
rect 18371 25721 18383 25755
rect 18325 25715 18383 25721
rect 26142 25712 26148 25764
rect 26200 25712 26206 25764
rect 27982 25712 27988 25764
rect 28040 25752 28046 25764
rect 34128 25752 34156 25792
rect 35158 25780 35164 25832
rect 35216 25820 35222 25832
rect 35437 25823 35495 25829
rect 35437 25820 35449 25823
rect 35216 25792 35449 25820
rect 35216 25780 35222 25792
rect 35437 25789 35449 25792
rect 35483 25789 35495 25823
rect 35437 25783 35495 25789
rect 35986 25780 35992 25832
rect 36044 25820 36050 25832
rect 36998 25820 37004 25832
rect 36044 25792 37004 25820
rect 36044 25780 36050 25792
rect 36998 25780 37004 25792
rect 37056 25780 37062 25832
rect 38197 25823 38255 25829
rect 38197 25789 38209 25823
rect 38243 25789 38255 25823
rect 38304 25820 38332 25860
rect 38470 25848 38476 25900
rect 38528 25848 38534 25900
rect 38746 25820 38752 25832
rect 38304 25792 38752 25820
rect 38197 25783 38255 25789
rect 28040 25724 34156 25752
rect 28040 25712 28046 25724
rect 34422 25712 34428 25764
rect 34480 25712 34486 25764
rect 35713 25755 35771 25761
rect 35713 25752 35725 25755
rect 34716 25724 35725 25752
rect 34716 25696 34744 25724
rect 35713 25721 35725 25724
rect 35759 25752 35771 25755
rect 38212 25752 38240 25783
rect 38746 25780 38752 25792
rect 38804 25780 38810 25832
rect 35759 25724 38240 25752
rect 35759 25721 35771 25724
rect 35713 25715 35771 25721
rect 5534 25644 5540 25696
rect 5592 25644 5598 25696
rect 7006 25644 7012 25696
rect 7064 25644 7070 25696
rect 10318 25644 10324 25696
rect 10376 25644 10382 25696
rect 12158 25644 12164 25696
rect 12216 25684 12222 25696
rect 12621 25687 12679 25693
rect 12621 25684 12633 25687
rect 12216 25656 12633 25684
rect 12216 25644 12222 25656
rect 12621 25653 12633 25656
rect 12667 25653 12679 25687
rect 12621 25647 12679 25653
rect 13541 25687 13599 25693
rect 13541 25653 13553 25687
rect 13587 25684 13599 25687
rect 14458 25684 14464 25696
rect 13587 25656 14464 25684
rect 13587 25653 13599 25656
rect 13541 25647 13599 25653
rect 14458 25644 14464 25656
rect 14516 25644 14522 25696
rect 16850 25644 16856 25696
rect 16908 25684 16914 25696
rect 18969 25687 19027 25693
rect 18969 25684 18981 25687
rect 16908 25656 18981 25684
rect 16908 25644 16914 25656
rect 18969 25653 18981 25656
rect 19015 25684 19027 25687
rect 23566 25684 23572 25696
rect 19015 25656 23572 25684
rect 19015 25653 19027 25656
rect 18969 25647 19027 25653
rect 23566 25644 23572 25656
rect 23624 25644 23630 25696
rect 28994 25644 29000 25696
rect 29052 25644 29058 25696
rect 30742 25644 30748 25696
rect 30800 25644 30806 25696
rect 31938 25644 31944 25696
rect 31996 25684 32002 25696
rect 32122 25684 32128 25696
rect 31996 25656 32128 25684
rect 31996 25644 32002 25656
rect 32122 25644 32128 25656
rect 32180 25684 32186 25696
rect 32309 25687 32367 25693
rect 32309 25684 32321 25687
rect 32180 25656 32321 25684
rect 32180 25644 32186 25656
rect 32309 25653 32321 25656
rect 32355 25653 32367 25687
rect 32309 25647 32367 25653
rect 34057 25687 34115 25693
rect 34057 25653 34069 25687
rect 34103 25684 34115 25687
rect 34698 25684 34704 25696
rect 34103 25656 34704 25684
rect 34103 25653 34115 25656
rect 34057 25647 34115 25653
rect 34698 25644 34704 25656
rect 34756 25644 34762 25696
rect 35253 25687 35311 25693
rect 35253 25653 35265 25687
rect 35299 25684 35311 25687
rect 35802 25684 35808 25696
rect 35299 25656 35808 25684
rect 35299 25653 35311 25656
rect 35253 25647 35311 25653
rect 35802 25644 35808 25656
rect 35860 25644 35866 25696
rect 35897 25687 35955 25693
rect 35897 25653 35909 25687
rect 35943 25684 35955 25687
rect 36354 25684 36360 25696
rect 35943 25656 36360 25684
rect 35943 25653 35955 25656
rect 35897 25647 35955 25653
rect 36354 25644 36360 25656
rect 36412 25644 36418 25696
rect 37829 25687 37887 25693
rect 37829 25653 37841 25687
rect 37875 25684 37887 25687
rect 38010 25684 38016 25696
rect 37875 25656 38016 25684
rect 37875 25653 37887 25656
rect 37829 25647 37887 25653
rect 38010 25644 38016 25656
rect 38068 25644 38074 25696
rect 1104 25594 40572 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 40572 25594
rect 1104 25520 40572 25542
rect 3970 25440 3976 25492
rect 4028 25480 4034 25492
rect 4525 25483 4583 25489
rect 4525 25480 4537 25483
rect 4028 25452 4537 25480
rect 4028 25440 4034 25452
rect 4525 25449 4537 25452
rect 4571 25449 4583 25483
rect 4525 25443 4583 25449
rect 6362 25440 6368 25492
rect 6420 25440 6426 25492
rect 6914 25440 6920 25492
rect 6972 25480 6978 25492
rect 7285 25483 7343 25489
rect 7285 25480 7297 25483
rect 6972 25452 7297 25480
rect 6972 25440 6978 25452
rect 7285 25449 7297 25452
rect 7331 25480 7343 25483
rect 8110 25480 8116 25492
rect 7331 25452 8116 25480
rect 7331 25449 7343 25452
rect 7285 25443 7343 25449
rect 8110 25440 8116 25452
rect 8168 25440 8174 25492
rect 11241 25483 11299 25489
rect 11241 25449 11253 25483
rect 11287 25480 11299 25483
rect 11330 25480 11336 25492
rect 11287 25452 11336 25480
rect 11287 25449 11299 25452
rect 11241 25443 11299 25449
rect 11330 25440 11336 25452
rect 11388 25440 11394 25492
rect 13354 25440 13360 25492
rect 13412 25480 13418 25492
rect 15102 25480 15108 25492
rect 13412 25452 15108 25480
rect 13412 25440 13418 25452
rect 15102 25440 15108 25452
rect 15160 25440 15166 25492
rect 15473 25483 15531 25489
rect 15473 25449 15485 25483
rect 15519 25480 15531 25483
rect 15654 25480 15660 25492
rect 15519 25452 15660 25480
rect 15519 25449 15531 25452
rect 15473 25443 15531 25449
rect 15654 25440 15660 25452
rect 15712 25480 15718 25492
rect 16209 25483 16267 25489
rect 16209 25480 16221 25483
rect 15712 25452 16221 25480
rect 15712 25440 15718 25452
rect 16209 25449 16221 25452
rect 16255 25449 16267 25483
rect 17862 25480 17868 25492
rect 16209 25443 16267 25449
rect 16868 25452 17868 25480
rect 7466 25372 7472 25424
rect 7524 25412 7530 25424
rect 16868 25412 16896 25452
rect 17862 25440 17868 25452
rect 17920 25440 17926 25492
rect 20349 25483 20407 25489
rect 20349 25449 20361 25483
rect 20395 25480 20407 25483
rect 20622 25480 20628 25492
rect 20395 25452 20628 25480
rect 20395 25449 20407 25452
rect 20349 25443 20407 25449
rect 20622 25440 20628 25452
rect 20680 25440 20686 25492
rect 22278 25440 22284 25492
rect 22336 25480 22342 25492
rect 23753 25483 23811 25489
rect 23753 25480 23765 25483
rect 22336 25452 23765 25480
rect 22336 25440 22342 25452
rect 23753 25449 23765 25452
rect 23799 25480 23811 25483
rect 24762 25480 24768 25492
rect 23799 25452 24768 25480
rect 23799 25449 23811 25452
rect 23753 25443 23811 25449
rect 24762 25440 24768 25452
rect 24820 25440 24826 25492
rect 24854 25440 24860 25492
rect 24912 25440 24918 25492
rect 25222 25440 25228 25492
rect 25280 25480 25286 25492
rect 30377 25483 30435 25489
rect 25280 25452 28580 25480
rect 25280 25440 25286 25452
rect 7524 25384 16896 25412
rect 7524 25372 7530 25384
rect 17402 25372 17408 25424
rect 17460 25412 17466 25424
rect 25961 25415 26019 25421
rect 25961 25412 25973 25415
rect 17460 25384 25973 25412
rect 17460 25372 17466 25384
rect 25961 25381 25973 25384
rect 26007 25381 26019 25415
rect 28442 25412 28448 25424
rect 25961 25375 26019 25381
rect 26436 25384 28448 25412
rect 1578 25304 1584 25356
rect 1636 25344 1642 25356
rect 2866 25344 2872 25356
rect 1636 25316 2872 25344
rect 1636 25304 1642 25316
rect 2866 25304 2872 25316
rect 2924 25344 2930 25356
rect 3694 25344 3700 25356
rect 2924 25316 3700 25344
rect 2924 25304 2930 25316
rect 3694 25304 3700 25316
rect 3752 25304 3758 25356
rect 4798 25304 4804 25356
rect 4856 25344 4862 25356
rect 4985 25347 5043 25353
rect 4985 25344 4997 25347
rect 4856 25316 4997 25344
rect 4856 25304 4862 25316
rect 4985 25313 4997 25316
rect 5031 25313 5043 25347
rect 4985 25307 5043 25313
rect 5169 25347 5227 25353
rect 5169 25313 5181 25347
rect 5215 25344 5227 25347
rect 5258 25344 5264 25356
rect 5215 25316 5264 25344
rect 5215 25313 5227 25316
rect 5169 25307 5227 25313
rect 5258 25304 5264 25316
rect 5316 25304 5322 25356
rect 5350 25304 5356 25356
rect 5408 25344 5414 25356
rect 7926 25344 7932 25356
rect 5408 25316 6684 25344
rect 5408 25304 5414 25316
rect 4433 25279 4491 25285
rect 4433 25245 4445 25279
rect 4479 25245 4491 25279
rect 4433 25239 4491 25245
rect 4893 25279 4951 25285
rect 4893 25245 4905 25279
rect 4939 25276 4951 25279
rect 5534 25276 5540 25288
rect 4939 25248 5540 25276
rect 4939 25245 4951 25248
rect 4893 25239 4951 25245
rect 1854 25168 1860 25220
rect 1912 25168 1918 25220
rect 3142 25208 3148 25220
rect 3082 25180 3148 25208
rect 3142 25168 3148 25180
rect 3200 25168 3206 25220
rect 4448 25208 4476 25239
rect 5534 25236 5540 25248
rect 5592 25236 5598 25288
rect 5626 25236 5632 25288
rect 5684 25276 5690 25288
rect 5721 25279 5779 25285
rect 5721 25276 5733 25279
rect 5684 25248 5733 25276
rect 5684 25236 5690 25248
rect 5721 25245 5733 25248
rect 5767 25245 5779 25279
rect 5721 25239 5779 25245
rect 6089 25279 6147 25285
rect 6089 25245 6101 25279
rect 6135 25276 6147 25279
rect 6178 25276 6184 25288
rect 6135 25248 6184 25276
rect 6135 25245 6147 25248
rect 6089 25239 6147 25245
rect 6178 25236 6184 25248
rect 6236 25236 6242 25288
rect 6270 25236 6276 25288
rect 6328 25236 6334 25288
rect 6454 25236 6460 25288
rect 6512 25276 6518 25288
rect 6656 25285 6684 25316
rect 6932 25316 7932 25344
rect 6932 25285 6960 25316
rect 7926 25304 7932 25316
rect 7984 25304 7990 25356
rect 8478 25304 8484 25356
rect 8536 25304 8542 25356
rect 9122 25304 9128 25356
rect 9180 25344 9186 25356
rect 13722 25344 13728 25356
rect 9180 25316 13728 25344
rect 9180 25304 9186 25316
rect 13722 25304 13728 25316
rect 13780 25304 13786 25356
rect 15838 25344 15844 25356
rect 15580 25316 15844 25344
rect 6549 25279 6607 25285
rect 6549 25276 6561 25279
rect 6512 25248 6561 25276
rect 6512 25236 6518 25248
rect 6549 25245 6561 25248
rect 6595 25245 6607 25279
rect 6549 25239 6607 25245
rect 6641 25279 6699 25285
rect 6641 25245 6653 25279
rect 6687 25245 6699 25279
rect 6641 25239 6699 25245
rect 6917 25279 6975 25285
rect 6917 25245 6929 25279
rect 6963 25245 6975 25279
rect 6917 25239 6975 25245
rect 7006 25236 7012 25288
rect 7064 25236 7070 25288
rect 7282 25276 7288 25288
rect 7208 25248 7288 25276
rect 5810 25208 5816 25220
rect 3344 25180 5816 25208
rect 3344 25149 3372 25180
rect 5810 25168 5816 25180
rect 5868 25168 5874 25220
rect 5905 25211 5963 25217
rect 5905 25177 5917 25211
rect 5951 25177 5963 25211
rect 5905 25171 5963 25177
rect 5997 25211 6055 25217
rect 5997 25177 6009 25211
rect 6043 25208 6055 25211
rect 6288 25208 6316 25236
rect 6043 25180 6316 25208
rect 6733 25211 6791 25217
rect 6043 25177 6055 25180
rect 5997 25171 6055 25177
rect 6733 25177 6745 25211
rect 6779 25208 6791 25211
rect 7098 25208 7104 25220
rect 6779 25180 7104 25208
rect 6779 25177 6791 25180
rect 6733 25171 6791 25177
rect 3329 25143 3387 25149
rect 3329 25109 3341 25143
rect 3375 25109 3387 25143
rect 3329 25103 3387 25109
rect 3786 25100 3792 25152
rect 3844 25100 3850 25152
rect 5534 25100 5540 25152
rect 5592 25140 5598 25152
rect 5920 25140 5948 25171
rect 7098 25168 7104 25180
rect 7156 25168 7162 25220
rect 7208 25217 7236 25248
rect 7282 25236 7288 25248
rect 7340 25276 7346 25288
rect 8294 25276 8300 25288
rect 7340 25248 8300 25276
rect 7340 25236 7346 25248
rect 8294 25236 8300 25248
rect 8352 25276 8358 25288
rect 9030 25276 9036 25288
rect 8352 25248 9036 25276
rect 8352 25236 8358 25248
rect 9030 25236 9036 25248
rect 9088 25236 9094 25288
rect 9398 25236 9404 25288
rect 9456 25276 9462 25288
rect 9493 25279 9551 25285
rect 9493 25276 9505 25279
rect 9456 25248 9505 25276
rect 9456 25236 9462 25248
rect 9493 25245 9505 25248
rect 9539 25245 9551 25279
rect 9493 25239 9551 25245
rect 11054 25236 11060 25288
rect 11112 25236 11118 25288
rect 11238 25236 11244 25288
rect 11296 25276 11302 25288
rect 11296 25248 11468 25276
rect 11296 25236 11302 25248
rect 7193 25211 7251 25217
rect 7193 25177 7205 25211
rect 7239 25177 7251 25211
rect 8941 25211 8999 25217
rect 8941 25208 8953 25211
rect 7193 25171 7251 25177
rect 8312 25180 8953 25208
rect 5592 25112 5948 25140
rect 6273 25143 6331 25149
rect 5592 25100 5598 25112
rect 6273 25109 6285 25143
rect 6319 25140 6331 25143
rect 6454 25140 6460 25152
rect 6319 25112 6460 25140
rect 6319 25109 6331 25112
rect 6273 25103 6331 25109
rect 6454 25100 6460 25112
rect 6512 25100 6518 25152
rect 7558 25100 7564 25152
rect 7616 25140 7622 25152
rect 8312 25149 8340 25180
rect 8941 25177 8953 25180
rect 8987 25177 8999 25211
rect 11072 25208 11100 25236
rect 11440 25217 11468 25248
rect 11974 25236 11980 25288
rect 12032 25276 12038 25288
rect 15580 25276 15608 25316
rect 15838 25304 15844 25316
rect 15896 25304 15902 25356
rect 18693 25347 18751 25353
rect 18693 25313 18705 25347
rect 18739 25344 18751 25347
rect 19058 25344 19064 25356
rect 18739 25316 19064 25344
rect 18739 25313 18751 25316
rect 18693 25307 18751 25313
rect 19058 25304 19064 25316
rect 19116 25304 19122 25356
rect 20806 25344 20812 25356
rect 19306 25316 20812 25344
rect 16298 25276 16304 25288
rect 12032 25248 15608 25276
rect 15672 25248 16304 25276
rect 12032 25236 12038 25248
rect 11425 25211 11483 25217
rect 11072 25180 11376 25208
rect 8941 25171 8999 25177
rect 7929 25143 7987 25149
rect 7929 25140 7941 25143
rect 7616 25112 7941 25140
rect 7616 25100 7622 25112
rect 7929 25109 7941 25112
rect 7975 25109 7987 25143
rect 7929 25103 7987 25109
rect 8297 25143 8355 25149
rect 8297 25109 8309 25143
rect 8343 25109 8355 25143
rect 8297 25103 8355 25109
rect 8386 25100 8392 25152
rect 8444 25100 8450 25152
rect 9766 25100 9772 25152
rect 9824 25140 9830 25152
rect 11238 25149 11244 25152
rect 11057 25143 11115 25149
rect 11057 25140 11069 25143
rect 9824 25112 11069 25140
rect 9824 25100 9830 25112
rect 11057 25109 11069 25112
rect 11103 25109 11115 25143
rect 11057 25103 11115 25109
rect 11225 25143 11244 25149
rect 11225 25109 11237 25143
rect 11225 25103 11244 25109
rect 11238 25100 11244 25103
rect 11296 25100 11302 25152
rect 11348 25140 11376 25180
rect 11425 25177 11437 25211
rect 11471 25208 11483 25211
rect 14550 25208 14556 25220
rect 11471 25180 14556 25208
rect 11471 25177 11483 25180
rect 11425 25171 11483 25177
rect 14550 25168 14556 25180
rect 14608 25168 14614 25220
rect 15672 25217 15700 25248
rect 16298 25236 16304 25248
rect 16356 25236 16362 25288
rect 16390 25236 16396 25288
rect 16448 25276 16454 25288
rect 16485 25279 16543 25285
rect 16485 25276 16497 25279
rect 16448 25248 16497 25276
rect 16448 25236 16454 25248
rect 16485 25245 16497 25248
rect 16531 25276 16543 25279
rect 18509 25279 18567 25285
rect 16531 25248 18460 25276
rect 16531 25245 16543 25248
rect 16485 25239 16543 25245
rect 15657 25211 15715 25217
rect 15657 25177 15669 25211
rect 15703 25177 15715 25211
rect 15657 25171 15715 25177
rect 16209 25211 16267 25217
rect 16209 25177 16221 25211
rect 16255 25208 16267 25211
rect 17310 25208 17316 25220
rect 16255 25180 17316 25208
rect 16255 25177 16267 25180
rect 16209 25171 16267 25177
rect 17310 25168 17316 25180
rect 17368 25168 17374 25220
rect 15470 25149 15476 25152
rect 15289 25143 15347 25149
rect 15289 25140 15301 25143
rect 11348 25112 15301 25140
rect 15289 25109 15301 25112
rect 15335 25109 15347 25143
rect 15289 25103 15347 25109
rect 15457 25143 15476 25149
rect 15457 25109 15469 25143
rect 15457 25103 15476 25109
rect 15470 25100 15476 25103
rect 15528 25100 15534 25152
rect 16298 25100 16304 25152
rect 16356 25140 16362 25152
rect 16393 25143 16451 25149
rect 16393 25140 16405 25143
rect 16356 25112 16405 25140
rect 16356 25100 16362 25112
rect 16393 25109 16405 25112
rect 16439 25140 16451 25143
rect 17126 25140 17132 25152
rect 16439 25112 17132 25140
rect 16439 25109 16451 25112
rect 16393 25103 16451 25109
rect 17126 25100 17132 25112
rect 17184 25100 17190 25152
rect 18138 25100 18144 25152
rect 18196 25140 18202 25152
rect 18325 25143 18383 25149
rect 18325 25140 18337 25143
rect 18196 25112 18337 25140
rect 18196 25100 18202 25112
rect 18325 25109 18337 25112
rect 18371 25109 18383 25143
rect 18432 25140 18460 25248
rect 18509 25245 18521 25279
rect 18555 25276 18567 25279
rect 19306 25276 19334 25316
rect 20806 25304 20812 25316
rect 20864 25304 20870 25356
rect 21450 25304 21456 25356
rect 21508 25344 21514 25356
rect 23014 25344 23020 25356
rect 21508 25316 23020 25344
rect 21508 25304 21514 25316
rect 23014 25304 23020 25316
rect 23072 25344 23078 25356
rect 23293 25347 23351 25353
rect 23293 25344 23305 25347
rect 23072 25316 23305 25344
rect 23072 25304 23078 25316
rect 23293 25313 23305 25316
rect 23339 25313 23351 25347
rect 23293 25307 23351 25313
rect 23477 25347 23535 25353
rect 23477 25313 23489 25347
rect 23523 25344 23535 25347
rect 23658 25344 23664 25356
rect 23523 25316 23664 25344
rect 23523 25313 23535 25316
rect 23477 25307 23535 25313
rect 23658 25304 23664 25316
rect 23716 25304 23722 25356
rect 24394 25304 24400 25356
rect 24452 25344 24458 25356
rect 25225 25347 25283 25353
rect 25225 25344 25237 25347
rect 24452 25316 25237 25344
rect 24452 25304 24458 25316
rect 25225 25313 25237 25316
rect 25271 25313 25283 25347
rect 25225 25307 25283 25313
rect 25317 25347 25375 25353
rect 25317 25313 25329 25347
rect 25363 25344 25375 25347
rect 25406 25344 25412 25356
rect 25363 25316 25412 25344
rect 25363 25313 25375 25316
rect 25317 25307 25375 25313
rect 25406 25304 25412 25316
rect 25464 25304 25470 25356
rect 26436 25344 26464 25384
rect 28442 25372 28448 25384
rect 28500 25372 28506 25424
rect 25992 25316 26464 25344
rect 26513 25347 26571 25353
rect 18555 25248 19334 25276
rect 18555 25245 18567 25248
rect 18509 25239 18567 25245
rect 20254 25236 20260 25288
rect 20312 25236 20318 25288
rect 20441 25279 20499 25285
rect 20441 25245 20453 25279
rect 20487 25276 20499 25279
rect 21082 25276 21088 25288
rect 20487 25248 21088 25276
rect 20487 25245 20499 25248
rect 20441 25239 20499 25245
rect 21082 25236 21088 25248
rect 21140 25236 21146 25288
rect 23385 25279 23443 25285
rect 23385 25245 23397 25279
rect 23431 25245 23443 25279
rect 23385 25239 23443 25245
rect 18598 25168 18604 25220
rect 18656 25208 18662 25220
rect 23106 25208 23112 25220
rect 18656 25180 23112 25208
rect 18656 25168 18662 25180
rect 23106 25168 23112 25180
rect 23164 25168 23170 25220
rect 23400 25208 23428 25239
rect 23566 25236 23572 25288
rect 23624 25276 23630 25288
rect 23624 25248 24348 25276
rect 23624 25236 23630 25248
rect 24210 25208 24216 25220
rect 23400 25180 24216 25208
rect 24210 25168 24216 25180
rect 24268 25168 24274 25220
rect 22738 25140 22744 25152
rect 18432 25112 22744 25140
rect 18325 25103 18383 25109
rect 22738 25100 22744 25112
rect 22796 25100 22802 25152
rect 24320 25140 24348 25248
rect 24578 25236 24584 25288
rect 24636 25276 24642 25288
rect 25041 25279 25099 25285
rect 25041 25276 25053 25279
rect 24636 25248 25053 25276
rect 24636 25236 24642 25248
rect 25041 25245 25053 25248
rect 25087 25245 25099 25279
rect 25041 25239 25099 25245
rect 25593 25279 25651 25285
rect 25593 25245 25605 25279
rect 25639 25276 25651 25279
rect 25682 25276 25688 25288
rect 25639 25248 25688 25276
rect 25639 25245 25651 25248
rect 25593 25239 25651 25245
rect 25682 25236 25688 25248
rect 25740 25236 25746 25288
rect 25866 25236 25872 25288
rect 25924 25236 25930 25288
rect 24486 25168 24492 25220
rect 24544 25208 24550 25220
rect 25409 25211 25467 25217
rect 25409 25208 25421 25211
rect 24544 25180 25421 25208
rect 24544 25168 24550 25180
rect 25409 25177 25421 25180
rect 25455 25177 25467 25211
rect 25409 25171 25467 25177
rect 25777 25143 25835 25149
rect 25777 25140 25789 25143
rect 24320 25112 25789 25140
rect 25777 25109 25789 25112
rect 25823 25140 25835 25143
rect 25992 25140 26020 25316
rect 26513 25313 26525 25347
rect 26559 25344 26571 25347
rect 26970 25344 26976 25356
rect 26559 25316 26976 25344
rect 26559 25313 26571 25316
rect 26513 25307 26571 25313
rect 26970 25304 26976 25316
rect 27028 25304 27034 25356
rect 26050 25236 26056 25288
rect 26108 25276 26114 25288
rect 26145 25279 26203 25285
rect 26145 25276 26157 25279
rect 26108 25248 26157 25276
rect 26108 25236 26114 25248
rect 26145 25245 26157 25248
rect 26191 25245 26203 25279
rect 26145 25239 26203 25245
rect 26234 25236 26240 25288
rect 26292 25236 26298 25288
rect 26329 25279 26387 25285
rect 26329 25245 26341 25279
rect 26375 25245 26387 25279
rect 26329 25239 26387 25245
rect 26344 25208 26372 25239
rect 26694 25236 26700 25288
rect 26752 25236 26758 25288
rect 26789 25279 26847 25285
rect 26789 25245 26801 25279
rect 26835 25276 26847 25279
rect 26878 25276 26884 25288
rect 26835 25248 26884 25276
rect 26835 25245 26847 25248
rect 26789 25239 26847 25245
rect 26878 25236 26884 25248
rect 26936 25236 26942 25288
rect 28552 25276 28580 25452
rect 30377 25449 30389 25483
rect 30423 25480 30435 25483
rect 30650 25480 30656 25492
rect 30423 25452 30656 25480
rect 30423 25449 30435 25452
rect 30377 25443 30435 25449
rect 30650 25440 30656 25452
rect 30708 25440 30714 25492
rect 31849 25483 31907 25489
rect 31849 25449 31861 25483
rect 31895 25480 31907 25483
rect 31938 25480 31944 25492
rect 31895 25452 31944 25480
rect 31895 25449 31907 25452
rect 31849 25443 31907 25449
rect 31938 25440 31944 25452
rect 31996 25440 32002 25492
rect 32585 25483 32643 25489
rect 32585 25449 32597 25483
rect 32631 25480 32643 25483
rect 32631 25452 33548 25480
rect 32631 25449 32643 25452
rect 32585 25443 32643 25449
rect 30561 25415 30619 25421
rect 30561 25381 30573 25415
rect 30607 25412 30619 25415
rect 33520 25412 33548 25452
rect 35802 25440 35808 25492
rect 35860 25480 35866 25492
rect 38013 25483 38071 25489
rect 38013 25480 38025 25483
rect 35860 25452 38025 25480
rect 35860 25440 35866 25452
rect 38013 25449 38025 25452
rect 38059 25449 38071 25483
rect 38013 25443 38071 25449
rect 33594 25412 33600 25424
rect 30607 25384 32260 25412
rect 30607 25381 30619 25384
rect 30561 25375 30619 25381
rect 28994 25304 29000 25356
rect 29052 25344 29058 25356
rect 30653 25347 30711 25353
rect 30653 25344 30665 25347
rect 29052 25316 30665 25344
rect 29052 25304 29058 25316
rect 30653 25313 30665 25316
rect 30699 25313 30711 25347
rect 30653 25307 30711 25313
rect 30926 25304 30932 25356
rect 30984 25304 30990 25356
rect 30742 25276 30748 25288
rect 28552 25248 30236 25276
rect 30438 25251 30748 25276
rect 30208 25217 30236 25248
rect 30423 25248 30748 25251
rect 30423 25245 30481 25248
rect 26513 25211 26571 25217
rect 26513 25208 26525 25211
rect 26344 25180 26525 25208
rect 26436 25152 26464 25180
rect 26513 25177 26525 25180
rect 26559 25177 26571 25211
rect 26513 25171 26571 25177
rect 30193 25211 30251 25217
rect 30193 25177 30205 25211
rect 30239 25177 30251 25211
rect 30423 25211 30435 25245
rect 30469 25211 30481 25245
rect 30742 25236 30748 25248
rect 30800 25276 30806 25288
rect 31665 25279 31723 25285
rect 31665 25276 31677 25279
rect 30800 25248 31677 25276
rect 30800 25236 30806 25248
rect 31665 25245 31677 25248
rect 31711 25276 31723 25279
rect 31754 25276 31760 25288
rect 31711 25248 31760 25276
rect 31711 25245 31723 25248
rect 31665 25239 31723 25245
rect 31754 25236 31760 25248
rect 31812 25236 31818 25288
rect 31846 25236 31852 25288
rect 31904 25276 31910 25288
rect 31941 25279 31999 25285
rect 31941 25276 31953 25279
rect 31904 25248 31953 25276
rect 31904 25236 31910 25248
rect 31941 25245 31953 25248
rect 31987 25245 31999 25279
rect 31941 25239 31999 25245
rect 32122 25236 32128 25288
rect 32180 25236 32186 25288
rect 32232 25276 32260 25384
rect 32692 25384 33180 25412
rect 33520 25384 33600 25412
rect 32692 25276 32720 25384
rect 32858 25304 32864 25356
rect 32916 25344 32922 25356
rect 32953 25347 33011 25353
rect 32953 25344 32965 25347
rect 32916 25316 32965 25344
rect 32916 25304 32922 25316
rect 32953 25313 32965 25316
rect 32999 25313 33011 25347
rect 32953 25307 33011 25313
rect 32232 25248 32720 25276
rect 33042 25236 33048 25288
rect 33100 25236 33106 25288
rect 33152 25285 33180 25384
rect 33594 25372 33600 25384
rect 33652 25412 33658 25424
rect 37090 25412 37096 25424
rect 33652 25384 37096 25412
rect 33652 25372 33658 25384
rect 37090 25372 37096 25384
rect 37148 25372 37154 25424
rect 34330 25304 34336 25356
rect 34388 25344 34394 25356
rect 35989 25347 36047 25353
rect 35989 25344 36001 25347
rect 34388 25316 36001 25344
rect 34388 25304 34394 25316
rect 35989 25313 36001 25316
rect 36035 25313 36047 25347
rect 36814 25344 36820 25356
rect 35989 25307 36047 25313
rect 36464 25316 36820 25344
rect 33137 25279 33195 25285
rect 33137 25245 33149 25279
rect 33183 25245 33195 25279
rect 33137 25239 33195 25245
rect 33318 25236 33324 25288
rect 33376 25236 33382 25288
rect 33413 25279 33471 25285
rect 33413 25245 33425 25279
rect 33459 25245 33471 25279
rect 33413 25239 33471 25245
rect 30423 25205 30481 25211
rect 33428 25208 33456 25239
rect 33686 25236 33692 25288
rect 33744 25236 33750 25288
rect 35526 25236 35532 25288
rect 35584 25236 35590 25288
rect 35621 25279 35679 25285
rect 35621 25245 35633 25279
rect 35667 25276 35679 25279
rect 35667 25248 36032 25276
rect 35667 25245 35679 25248
rect 35621 25239 35679 25245
rect 36004 25220 36032 25248
rect 36078 25236 36084 25288
rect 36136 25236 36142 25288
rect 36229 25279 36287 25285
rect 36229 25245 36241 25279
rect 36275 25245 36287 25279
rect 36229 25239 36287 25245
rect 30193 25171 30251 25177
rect 32140 25180 33456 25208
rect 33520 25180 33916 25208
rect 25823 25112 26020 25140
rect 25823 25109 25835 25112
rect 25777 25103 25835 25109
rect 26418 25100 26424 25152
rect 26476 25100 26482 25152
rect 30208 25140 30236 25171
rect 32140 25152 32168 25180
rect 31018 25140 31024 25152
rect 30208 25112 31024 25140
rect 31018 25100 31024 25112
rect 31076 25100 31082 25152
rect 32033 25143 32091 25149
rect 32033 25109 32045 25143
rect 32079 25140 32091 25143
rect 32122 25140 32128 25152
rect 32079 25112 32128 25140
rect 32079 25109 32091 25112
rect 32033 25103 32091 25109
rect 32122 25100 32128 25112
rect 32180 25100 32186 25152
rect 32398 25100 32404 25152
rect 32456 25100 32462 25152
rect 32582 25100 32588 25152
rect 32640 25140 32646 25152
rect 33520 25140 33548 25180
rect 32640 25112 33548 25140
rect 32640 25100 32646 25112
rect 33594 25100 33600 25152
rect 33652 25100 33658 25152
rect 33888 25149 33916 25180
rect 34790 25168 34796 25220
rect 34848 25208 34854 25220
rect 35897 25211 35955 25217
rect 35897 25208 35909 25211
rect 34848 25180 35909 25208
rect 34848 25168 34854 25180
rect 35897 25177 35909 25180
rect 35943 25177 35955 25211
rect 35897 25171 35955 25177
rect 35986 25168 35992 25220
rect 36044 25168 36050 25220
rect 36244 25208 36272 25239
rect 36354 25236 36360 25288
rect 36412 25236 36418 25288
rect 36464 25285 36492 25316
rect 36814 25304 36820 25316
rect 36872 25304 36878 25356
rect 37458 25304 37464 25356
rect 37516 25344 37522 25356
rect 38105 25347 38163 25353
rect 38105 25344 38117 25347
rect 37516 25316 38117 25344
rect 37516 25304 37522 25316
rect 38105 25313 38117 25316
rect 38151 25313 38163 25347
rect 38105 25307 38163 25313
rect 36449 25279 36507 25285
rect 36449 25245 36461 25279
rect 36495 25245 36507 25279
rect 36449 25239 36507 25245
rect 36587 25279 36645 25285
rect 36587 25245 36599 25279
rect 36633 25276 36645 25279
rect 36906 25276 36912 25288
rect 36633 25248 36912 25276
rect 36633 25245 36645 25248
rect 36587 25239 36645 25245
rect 36906 25236 36912 25248
rect 36964 25236 36970 25288
rect 38010 25236 38016 25288
rect 38068 25236 38074 25288
rect 36244 25180 36492 25208
rect 36464 25152 36492 25180
rect 33873 25143 33931 25149
rect 33873 25109 33885 25143
rect 33919 25109 33931 25143
rect 33873 25103 33931 25109
rect 35342 25100 35348 25152
rect 35400 25100 35406 25152
rect 35805 25143 35863 25149
rect 35805 25109 35817 25143
rect 35851 25140 35863 25143
rect 36170 25140 36176 25152
rect 35851 25112 36176 25140
rect 35851 25109 35863 25112
rect 35805 25103 35863 25109
rect 36170 25100 36176 25112
rect 36228 25100 36234 25152
rect 36446 25100 36452 25152
rect 36504 25100 36510 25152
rect 36725 25143 36783 25149
rect 36725 25109 36737 25143
rect 36771 25140 36783 25143
rect 37734 25140 37740 25152
rect 36771 25112 37740 25140
rect 36771 25109 36783 25112
rect 36725 25103 36783 25109
rect 37734 25100 37740 25112
rect 37792 25100 37798 25152
rect 38381 25143 38439 25149
rect 38381 25109 38393 25143
rect 38427 25140 38439 25143
rect 38470 25140 38476 25152
rect 38427 25112 38476 25140
rect 38427 25109 38439 25112
rect 38381 25103 38439 25109
rect 38470 25100 38476 25112
rect 38528 25100 38534 25152
rect 1104 25050 40572 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 40572 25050
rect 1104 24976 40572 24998
rect 1854 24896 1860 24948
rect 1912 24936 1918 24948
rect 2593 24939 2651 24945
rect 2593 24936 2605 24939
rect 1912 24908 2605 24936
rect 1912 24896 1918 24908
rect 2593 24905 2605 24908
rect 2639 24905 2651 24939
rect 2593 24899 2651 24905
rect 2961 24939 3019 24945
rect 2961 24905 2973 24939
rect 3007 24936 3019 24939
rect 3786 24936 3792 24948
rect 3007 24908 3792 24936
rect 3007 24905 3019 24908
rect 2961 24899 3019 24905
rect 3786 24896 3792 24908
rect 3844 24896 3850 24948
rect 5258 24896 5264 24948
rect 5316 24936 5322 24948
rect 8478 24936 8484 24948
rect 5316 24908 8484 24936
rect 5316 24896 5322 24908
rect 8478 24896 8484 24908
rect 8536 24896 8542 24948
rect 9033 24939 9091 24945
rect 9033 24905 9045 24939
rect 9079 24905 9091 24939
rect 9033 24899 9091 24905
rect 11057 24939 11115 24945
rect 11057 24905 11069 24939
rect 11103 24905 11115 24939
rect 11974 24936 11980 24948
rect 11057 24899 11115 24905
rect 11900 24908 11980 24936
rect 3053 24871 3111 24877
rect 3053 24837 3065 24871
rect 3099 24868 3111 24871
rect 3510 24868 3516 24880
rect 3099 24840 3516 24868
rect 3099 24837 3111 24840
rect 3053 24831 3111 24837
rect 3510 24828 3516 24840
rect 3568 24868 3574 24880
rect 4706 24868 4712 24880
rect 3568 24840 4712 24868
rect 3568 24828 3574 24840
rect 4706 24828 4712 24840
rect 4764 24828 4770 24880
rect 7558 24828 7564 24880
rect 7616 24828 7622 24880
rect 9048 24868 9076 24899
rect 9398 24868 9404 24880
rect 9048 24840 9404 24868
rect 9398 24828 9404 24840
rect 9456 24828 9462 24880
rect 10781 24871 10839 24877
rect 10781 24837 10793 24871
rect 10827 24868 10839 24871
rect 10962 24868 10968 24880
rect 10827 24840 10968 24868
rect 10827 24837 10839 24840
rect 10781 24831 10839 24837
rect 10962 24828 10968 24840
rect 11020 24828 11026 24880
rect 5258 24800 5264 24812
rect 3252 24772 5264 24800
rect 3252 24741 3280 24772
rect 5258 24760 5264 24772
rect 5316 24760 5322 24812
rect 5350 24760 5356 24812
rect 5408 24800 5414 24812
rect 5445 24803 5503 24809
rect 5445 24800 5457 24803
rect 5408 24772 5457 24800
rect 5408 24760 5414 24772
rect 5445 24769 5457 24772
rect 5491 24769 5503 24803
rect 5445 24763 5503 24769
rect 5534 24760 5540 24812
rect 5592 24800 5598 24812
rect 5629 24803 5687 24809
rect 5629 24800 5641 24803
rect 5592 24772 5641 24800
rect 5592 24760 5598 24772
rect 5629 24769 5641 24772
rect 5675 24769 5687 24803
rect 5629 24763 5687 24769
rect 5718 24760 5724 24812
rect 5776 24760 5782 24812
rect 5813 24803 5871 24809
rect 5813 24769 5825 24803
rect 5859 24800 5871 24803
rect 6086 24800 6092 24812
rect 5859 24772 6092 24800
rect 5859 24769 5871 24772
rect 5813 24763 5871 24769
rect 6086 24760 6092 24772
rect 6144 24760 6150 24812
rect 9306 24809 9312 24812
rect 9304 24800 9312 24809
rect 3237 24735 3295 24741
rect 3237 24701 3249 24735
rect 3283 24701 3295 24735
rect 3237 24695 3295 24701
rect 3878 24692 3884 24744
rect 3936 24732 3942 24744
rect 3973 24735 4031 24741
rect 3973 24732 3985 24735
rect 3936 24704 3985 24732
rect 3936 24692 3942 24704
rect 3973 24701 3985 24704
rect 4019 24701 4031 24735
rect 3973 24695 4031 24701
rect 7285 24735 7343 24741
rect 7285 24701 7297 24735
rect 7331 24701 7343 24735
rect 8680 24732 8708 24786
rect 9267 24772 9312 24800
rect 9304 24763 9312 24772
rect 9306 24760 9312 24763
rect 9364 24760 9370 24812
rect 9490 24760 9496 24812
rect 9548 24760 9554 24812
rect 9674 24760 9680 24812
rect 9732 24760 9738 24812
rect 9766 24760 9772 24812
rect 9824 24760 9830 24812
rect 10410 24760 10416 24812
rect 10468 24760 10474 24812
rect 10505 24803 10563 24809
rect 10505 24769 10517 24803
rect 10551 24769 10563 24803
rect 10505 24763 10563 24769
rect 9508 24732 9536 24760
rect 10428 24732 10456 24760
rect 8680 24704 9260 24732
rect 9508 24704 10456 24732
rect 10520 24732 10548 24763
rect 10594 24760 10600 24812
rect 10652 24800 10658 24812
rect 10689 24803 10747 24809
rect 10689 24800 10701 24803
rect 10652 24772 10701 24800
rect 10652 24760 10658 24772
rect 10689 24769 10701 24772
rect 10735 24769 10747 24803
rect 10689 24763 10747 24769
rect 10870 24760 10876 24812
rect 10928 24760 10934 24812
rect 11072 24800 11100 24899
rect 11900 24877 11928 24908
rect 11974 24896 11980 24908
rect 12032 24896 12038 24948
rect 12161 24939 12219 24945
rect 12161 24905 12173 24939
rect 12207 24905 12219 24939
rect 12161 24899 12219 24905
rect 11885 24871 11943 24877
rect 11885 24837 11897 24871
rect 11931 24837 11943 24871
rect 11885 24831 11943 24837
rect 11517 24803 11575 24809
rect 11517 24800 11529 24803
rect 11072 24772 11529 24800
rect 11517 24769 11529 24772
rect 11563 24769 11575 24803
rect 11517 24763 11575 24769
rect 11610 24803 11668 24809
rect 11610 24769 11622 24803
rect 11656 24769 11668 24803
rect 11610 24763 11668 24769
rect 10520 24704 10640 24732
rect 7285 24695 7343 24701
rect 3694 24624 3700 24676
rect 3752 24664 3758 24676
rect 7300 24664 7328 24695
rect 3752 24636 7328 24664
rect 9232 24664 9260 24704
rect 9490 24664 9496 24676
rect 9232 24636 9496 24664
rect 3752 24624 3758 24636
rect 9490 24624 9496 24636
rect 9548 24624 9554 24676
rect 2958 24556 2964 24608
rect 3016 24596 3022 24608
rect 3421 24599 3479 24605
rect 3421 24596 3433 24599
rect 3016 24568 3433 24596
rect 3016 24556 3022 24568
rect 3421 24565 3433 24568
rect 3467 24565 3479 24599
rect 3421 24559 3479 24565
rect 5902 24556 5908 24608
rect 5960 24596 5966 24608
rect 5997 24599 6055 24605
rect 5997 24596 6009 24599
rect 5960 24568 6009 24596
rect 5960 24556 5966 24568
rect 5997 24565 6009 24568
rect 6043 24565 6055 24599
rect 5997 24559 6055 24565
rect 6730 24556 6736 24608
rect 6788 24596 6794 24608
rect 7282 24596 7288 24608
rect 6788 24568 7288 24596
rect 6788 24556 6794 24568
rect 7282 24556 7288 24568
rect 7340 24556 7346 24608
rect 7374 24556 7380 24608
rect 7432 24596 7438 24608
rect 8110 24596 8116 24608
rect 7432 24568 8116 24596
rect 7432 24556 7438 24568
rect 8110 24556 8116 24568
rect 8168 24556 8174 24608
rect 9122 24556 9128 24608
rect 9180 24556 9186 24608
rect 10612 24596 10640 24704
rect 10778 24624 10784 24676
rect 10836 24664 10842 24676
rect 11624 24664 11652 24763
rect 11790 24760 11796 24812
rect 11848 24760 11854 24812
rect 11974 24760 11980 24812
rect 12032 24809 12038 24812
rect 12032 24800 12040 24809
rect 12176 24800 12204 24899
rect 12250 24896 12256 24948
rect 12308 24936 12314 24948
rect 15746 24936 15752 24948
rect 12308 24908 15752 24936
rect 12308 24896 12314 24908
rect 12452 24809 12480 24908
rect 15746 24896 15752 24908
rect 15804 24896 15810 24948
rect 16500 24908 17080 24936
rect 14384 24840 14596 24868
rect 12253 24803 12311 24809
rect 12253 24800 12265 24803
rect 12032 24772 12077 24800
rect 12176 24772 12265 24800
rect 12032 24763 12040 24772
rect 12253 24769 12265 24772
rect 12299 24769 12311 24803
rect 12253 24763 12311 24769
rect 12437 24803 12495 24809
rect 12437 24769 12449 24803
rect 12483 24769 12495 24803
rect 12437 24763 12495 24769
rect 12032 24760 12038 24763
rect 14090 24760 14096 24812
rect 14148 24800 14154 24812
rect 14384 24800 14412 24840
rect 14148 24772 14412 24800
rect 14148 24760 14154 24772
rect 14458 24760 14464 24812
rect 14516 24760 14522 24812
rect 14568 24809 14596 24840
rect 14660 24840 14872 24868
rect 14660 24812 14688 24840
rect 14553 24803 14611 24809
rect 14553 24769 14565 24803
rect 14599 24769 14611 24803
rect 14553 24763 14611 24769
rect 14642 24760 14648 24812
rect 14700 24760 14706 24812
rect 14734 24760 14740 24812
rect 14792 24760 14798 24812
rect 14844 24809 14872 24840
rect 14829 24803 14887 24809
rect 14829 24769 14841 24803
rect 14875 24769 14887 24803
rect 14829 24763 14887 24769
rect 14921 24803 14979 24809
rect 14921 24769 14933 24803
rect 14967 24800 14979 24803
rect 15289 24803 15347 24809
rect 15289 24800 15301 24803
rect 14967 24772 15301 24800
rect 14967 24769 14979 24772
rect 14921 24763 14979 24769
rect 15289 24769 15301 24772
rect 15335 24769 15347 24803
rect 15289 24763 15347 24769
rect 11997 24732 12025 24760
rect 14936 24732 14964 24763
rect 15470 24760 15476 24812
rect 15528 24800 15534 24812
rect 16025 24803 16083 24809
rect 16025 24800 16037 24803
rect 15528 24772 16037 24800
rect 15528 24760 15534 24772
rect 16025 24769 16037 24772
rect 16071 24769 16083 24803
rect 16025 24763 16083 24769
rect 16209 24803 16267 24809
rect 16209 24769 16221 24803
rect 16255 24800 16267 24803
rect 16298 24800 16304 24812
rect 16255 24772 16304 24800
rect 16255 24769 16267 24772
rect 16209 24763 16267 24769
rect 16298 24760 16304 24772
rect 16356 24760 16362 24812
rect 16500 24809 16528 24908
rect 16959 24815 16987 24908
rect 17052 24868 17080 24908
rect 17126 24896 17132 24948
rect 17184 24936 17190 24948
rect 18598 24936 18604 24948
rect 17184 24908 18604 24936
rect 17184 24896 17190 24908
rect 18598 24896 18604 24908
rect 18656 24896 18662 24948
rect 20254 24896 20260 24948
rect 20312 24936 20318 24948
rect 20349 24939 20407 24945
rect 20349 24936 20361 24939
rect 20312 24908 20361 24936
rect 20312 24896 20318 24908
rect 20349 24905 20361 24908
rect 20395 24905 20407 24939
rect 20349 24899 20407 24905
rect 21266 24896 21272 24948
rect 21324 24896 21330 24948
rect 22005 24939 22063 24945
rect 22005 24905 22017 24939
rect 22051 24936 22063 24939
rect 22186 24936 22192 24948
rect 22051 24908 22192 24936
rect 22051 24905 22063 24908
rect 22005 24899 22063 24905
rect 22186 24896 22192 24908
rect 22244 24936 22250 24948
rect 22554 24936 22560 24948
rect 22244 24908 22560 24936
rect 22244 24896 22250 24908
rect 22554 24896 22560 24908
rect 22612 24896 22618 24948
rect 23934 24896 23940 24948
rect 23992 24936 23998 24948
rect 24765 24939 24823 24945
rect 23992 24908 24624 24936
rect 23992 24896 23998 24908
rect 17678 24868 17684 24880
rect 17052 24840 17684 24868
rect 17678 24828 17684 24840
rect 17736 24828 17742 24880
rect 18984 24840 19840 24868
rect 16944 24809 17002 24815
rect 16485 24803 16543 24809
rect 16485 24769 16497 24803
rect 16531 24769 16543 24803
rect 16944 24775 16956 24809
rect 16990 24775 17002 24809
rect 16944 24769 17002 24775
rect 17037 24803 17095 24809
rect 17037 24769 17049 24803
rect 17083 24769 17095 24803
rect 16485 24763 16543 24769
rect 17037 24763 17095 24769
rect 11997 24704 14964 24732
rect 15013 24735 15071 24741
rect 15013 24701 15025 24735
rect 15059 24732 15071 24735
rect 15194 24732 15200 24744
rect 15059 24704 15200 24732
rect 15059 24701 15071 24704
rect 15013 24695 15071 24701
rect 15194 24692 15200 24704
rect 15252 24692 15258 24744
rect 15654 24692 15660 24744
rect 15712 24692 15718 24744
rect 16393 24735 16451 24741
rect 16393 24701 16405 24735
rect 16439 24732 16451 24735
rect 17052 24732 17080 24763
rect 17126 24760 17132 24812
rect 17184 24760 17190 24812
rect 17310 24760 17316 24812
rect 17368 24760 17374 24812
rect 17402 24760 17408 24812
rect 17460 24800 17466 24812
rect 17460 24772 17632 24800
rect 17460 24760 17466 24772
rect 17328 24732 17356 24760
rect 17497 24735 17555 24741
rect 17497 24732 17509 24735
rect 16439 24704 17172 24732
rect 17328 24704 17509 24732
rect 16439 24701 16451 24704
rect 16393 24695 16451 24701
rect 10836 24636 11652 24664
rect 10836 24624 10842 24636
rect 15930 24624 15936 24676
rect 15988 24664 15994 24676
rect 16669 24667 16727 24673
rect 16669 24664 16681 24667
rect 15988 24636 16681 24664
rect 15988 24624 15994 24636
rect 16669 24633 16681 24636
rect 16715 24633 16727 24667
rect 17144 24664 17172 24704
rect 17497 24701 17509 24704
rect 17543 24701 17555 24735
rect 17497 24695 17555 24701
rect 17604 24664 17632 24772
rect 18506 24760 18512 24812
rect 18564 24800 18570 24812
rect 18984 24800 19012 24840
rect 18564 24772 19012 24800
rect 18564 24760 18570 24772
rect 19058 24760 19064 24812
rect 19116 24760 19122 24812
rect 18414 24692 18420 24744
rect 18472 24732 18478 24744
rect 18874 24732 18880 24744
rect 18472 24704 18880 24732
rect 18472 24692 18478 24704
rect 18874 24692 18880 24704
rect 18932 24732 18938 24744
rect 18969 24735 19027 24741
rect 18969 24732 18981 24735
rect 18932 24704 18981 24732
rect 18932 24692 18938 24704
rect 18969 24701 18981 24704
rect 19015 24701 19027 24735
rect 18969 24695 19027 24701
rect 17144 24636 17632 24664
rect 16669 24627 16727 24633
rect 12434 24596 12440 24608
rect 10612 24568 12440 24596
rect 12434 24556 12440 24568
rect 12492 24556 12498 24608
rect 12526 24556 12532 24608
rect 12584 24556 12590 24608
rect 12618 24556 12624 24608
rect 12676 24596 12682 24608
rect 14550 24596 14556 24608
rect 12676 24568 14556 24596
rect 12676 24556 12682 24568
rect 14550 24556 14556 24568
rect 14608 24596 14614 24608
rect 16114 24596 16120 24608
rect 14608 24568 16120 24596
rect 14608 24556 14614 24568
rect 16114 24556 16120 24568
rect 16172 24596 16178 24608
rect 17405 24599 17463 24605
rect 17405 24596 17417 24599
rect 16172 24568 17417 24596
rect 16172 24556 16178 24568
rect 17405 24565 17417 24568
rect 17451 24565 17463 24599
rect 19168 24596 19196 24840
rect 19812 24809 19840 24840
rect 19886 24828 19892 24880
rect 19944 24868 19950 24880
rect 19981 24871 20039 24877
rect 19981 24868 19993 24871
rect 19944 24840 19993 24868
rect 19944 24828 19950 24840
rect 19981 24837 19993 24840
rect 20027 24868 20039 24871
rect 20622 24868 20628 24880
rect 20027 24840 20628 24868
rect 20027 24837 20039 24840
rect 19981 24831 20039 24837
rect 20622 24828 20628 24840
rect 20680 24828 20686 24880
rect 21284 24868 21312 24896
rect 21100 24840 21312 24868
rect 19245 24803 19303 24809
rect 19245 24769 19257 24803
rect 19291 24769 19303 24803
rect 19245 24763 19303 24769
rect 19797 24803 19855 24809
rect 19797 24769 19809 24803
rect 19843 24769 19855 24803
rect 19797 24763 19855 24769
rect 19260 24664 19288 24763
rect 20070 24760 20076 24812
rect 20128 24760 20134 24812
rect 20165 24803 20223 24809
rect 20165 24769 20177 24803
rect 20211 24769 20223 24803
rect 20165 24763 20223 24769
rect 19334 24692 19340 24744
rect 19392 24732 19398 24744
rect 20180 24732 20208 24763
rect 20714 24760 20720 24812
rect 20772 24760 20778 24812
rect 21100 24809 21128 24840
rect 21818 24828 21824 24880
rect 21876 24868 21882 24880
rect 23952 24868 23980 24896
rect 21876 24840 23980 24868
rect 21876 24828 21882 24840
rect 24394 24828 24400 24880
rect 24452 24828 24458 24880
rect 21085 24803 21143 24809
rect 21085 24769 21097 24803
rect 21131 24769 21143 24803
rect 21085 24763 21143 24769
rect 21269 24803 21327 24809
rect 21269 24769 21281 24803
rect 21315 24769 21327 24803
rect 21269 24763 21327 24769
rect 21545 24803 21603 24809
rect 21545 24769 21557 24803
rect 21591 24769 21603 24803
rect 21545 24763 21603 24769
rect 21284 24732 21312 24763
rect 19392 24704 21312 24732
rect 19392 24692 19398 24704
rect 21082 24664 21088 24676
rect 19260 24636 21088 24664
rect 21082 24624 21088 24636
rect 21140 24624 21146 24676
rect 21284 24664 21312 24704
rect 21358 24692 21364 24744
rect 21416 24692 21422 24744
rect 21450 24692 21456 24744
rect 21508 24732 21514 24744
rect 21560 24732 21588 24763
rect 21910 24760 21916 24812
rect 21968 24809 21974 24812
rect 21968 24803 22004 24809
rect 21992 24769 22004 24803
rect 21968 24763 22004 24769
rect 21968 24760 21974 24763
rect 22278 24760 22284 24812
rect 22336 24800 22342 24812
rect 22465 24803 22523 24809
rect 22465 24800 22477 24803
rect 22336 24772 22477 24800
rect 22336 24760 22342 24772
rect 22465 24769 22477 24772
rect 22511 24769 22523 24803
rect 24305 24803 24363 24809
rect 24305 24800 24317 24803
rect 22465 24763 22523 24769
rect 24228 24772 24317 24800
rect 23658 24732 23664 24744
rect 21508 24704 23664 24732
rect 21508 24692 21514 24704
rect 23658 24692 23664 24704
rect 23716 24692 23722 24744
rect 22094 24664 22100 24676
rect 21284 24636 22100 24664
rect 22094 24624 22100 24636
rect 22152 24624 22158 24676
rect 21450 24596 21456 24608
rect 19168 24568 21456 24596
rect 17405 24559 17463 24565
rect 21450 24556 21456 24568
rect 21508 24556 21514 24608
rect 21818 24556 21824 24608
rect 21876 24556 21882 24608
rect 22370 24556 22376 24608
rect 22428 24556 22434 24608
rect 24228 24596 24256 24772
rect 24305 24769 24317 24772
rect 24351 24769 24363 24803
rect 24305 24763 24363 24769
rect 24486 24760 24492 24812
rect 24544 24760 24550 24812
rect 24596 24809 24624 24908
rect 24765 24905 24777 24939
rect 24811 24936 24823 24939
rect 25133 24939 25191 24945
rect 25133 24936 25145 24939
rect 24811 24908 25145 24936
rect 24811 24905 24823 24908
rect 24765 24899 24823 24905
rect 25133 24905 25145 24908
rect 25179 24936 25191 24939
rect 25682 24936 25688 24948
rect 25179 24908 25688 24936
rect 25179 24905 25191 24908
rect 25133 24899 25191 24905
rect 25682 24896 25688 24908
rect 25740 24896 25746 24948
rect 25958 24896 25964 24948
rect 26016 24945 26022 24948
rect 26016 24939 26035 24945
rect 26023 24905 26035 24939
rect 26970 24936 26976 24948
rect 26016 24899 26035 24905
rect 26344 24908 26976 24936
rect 26016 24896 26022 24899
rect 25593 24871 25651 24877
rect 25593 24837 25605 24871
rect 25639 24868 25651 24871
rect 25639 24840 25712 24868
rect 25639 24837 25651 24840
rect 25593 24831 25651 24837
rect 24581 24803 24639 24809
rect 24581 24769 24593 24803
rect 24627 24769 24639 24803
rect 24581 24763 24639 24769
rect 24762 24760 24768 24812
rect 24820 24760 24826 24812
rect 24857 24803 24915 24809
rect 24857 24769 24869 24803
rect 24903 24800 24915 24803
rect 24946 24800 24952 24812
rect 24903 24772 24952 24800
rect 24903 24769 24915 24772
rect 24857 24763 24915 24769
rect 24946 24760 24952 24772
rect 25004 24760 25010 24812
rect 25684 24790 25712 24840
rect 25774 24828 25780 24880
rect 25832 24828 25838 24880
rect 26344 24868 26372 24908
rect 26970 24896 26976 24908
rect 27028 24896 27034 24948
rect 31312 24908 31708 24936
rect 25992 24840 26372 24868
rect 26421 24871 26479 24877
rect 25992 24800 26020 24840
rect 26421 24837 26433 24871
rect 26467 24837 26479 24871
rect 26421 24831 26479 24837
rect 27816 24840 28120 24868
rect 26436 24800 26464 24831
rect 25792 24790 26020 24800
rect 25684 24772 26020 24790
rect 26068 24772 26464 24800
rect 25684 24762 25820 24772
rect 25041 24735 25099 24741
rect 25041 24701 25053 24735
rect 25087 24732 25099 24735
rect 25406 24732 25412 24744
rect 25087 24704 25412 24732
rect 25087 24701 25099 24704
rect 25041 24695 25099 24701
rect 25406 24692 25412 24704
rect 25464 24732 25470 24744
rect 26068 24732 26096 24772
rect 26510 24760 26516 24812
rect 26568 24800 26574 24812
rect 26568 24772 27200 24800
rect 26568 24760 26574 24772
rect 26878 24732 26884 24744
rect 25464 24704 26096 24732
rect 26160 24704 26884 24732
rect 25464 24692 25470 24704
rect 24670 24624 24676 24676
rect 24728 24664 24734 24676
rect 26160 24673 26188 24704
rect 26878 24692 26884 24704
rect 26936 24732 26942 24744
rect 26973 24735 27031 24741
rect 26973 24732 26985 24735
rect 26936 24704 26985 24732
rect 26936 24692 26942 24704
rect 26973 24701 26985 24704
rect 27019 24701 27031 24735
rect 26973 24695 27031 24701
rect 27062 24692 27068 24744
rect 27120 24692 27126 24744
rect 27172 24732 27200 24772
rect 27246 24760 27252 24812
rect 27304 24760 27310 24812
rect 27430 24760 27436 24812
rect 27488 24800 27494 24812
rect 27709 24803 27767 24809
rect 27709 24800 27721 24803
rect 27488 24772 27721 24800
rect 27488 24760 27494 24772
rect 27709 24769 27721 24772
rect 27755 24769 27767 24803
rect 27709 24763 27767 24769
rect 27816 24732 27844 24840
rect 27893 24803 27951 24809
rect 27893 24769 27905 24803
rect 27939 24800 27951 24803
rect 28092 24800 28120 24840
rect 28169 24803 28227 24809
rect 28169 24800 28181 24803
rect 27939 24772 28028 24800
rect 28092 24772 28181 24800
rect 27939 24769 27951 24772
rect 27893 24763 27951 24769
rect 27172 24704 27844 24732
rect 25593 24667 25651 24673
rect 25593 24664 25605 24667
rect 24728 24636 25605 24664
rect 24728 24624 24734 24636
rect 25593 24633 25605 24636
rect 25639 24633 25651 24667
rect 25593 24627 25651 24633
rect 26145 24667 26203 24673
rect 26145 24633 26157 24667
rect 26191 24633 26203 24667
rect 26145 24627 26203 24633
rect 26237 24667 26295 24673
rect 26237 24633 26249 24667
rect 26283 24664 26295 24667
rect 26326 24664 26332 24676
rect 26283 24636 26332 24664
rect 26283 24633 26295 24636
rect 26237 24627 26295 24633
rect 26326 24624 26332 24636
rect 26384 24624 26390 24676
rect 26789 24667 26847 24673
rect 26789 24633 26801 24667
rect 26835 24633 26847 24667
rect 26789 24627 26847 24633
rect 25682 24596 25688 24608
rect 24228 24568 25688 24596
rect 25682 24556 25688 24568
rect 25740 24556 25746 24608
rect 25774 24556 25780 24608
rect 25832 24596 25838 24608
rect 25961 24599 26019 24605
rect 25961 24596 25973 24599
rect 25832 24568 25973 24596
rect 25832 24556 25838 24568
rect 25961 24565 25973 24568
rect 26007 24565 26019 24599
rect 25961 24559 26019 24565
rect 26418 24556 26424 24608
rect 26476 24556 26482 24608
rect 26804 24596 26832 24627
rect 27154 24624 27160 24676
rect 27212 24664 27218 24676
rect 27433 24667 27491 24673
rect 27433 24664 27445 24667
rect 27212 24636 27445 24664
rect 27212 24624 27218 24636
rect 27433 24633 27445 24636
rect 27479 24633 27491 24667
rect 27433 24627 27491 24633
rect 28000 24608 28028 24772
rect 28169 24769 28181 24772
rect 28215 24769 28227 24803
rect 28169 24763 28227 24769
rect 28353 24803 28411 24809
rect 28353 24769 28365 24803
rect 28399 24769 28411 24803
rect 28353 24763 28411 24769
rect 28368 24732 28396 24763
rect 28534 24760 28540 24812
rect 28592 24760 28598 24812
rect 30469 24803 30527 24809
rect 30469 24769 30481 24803
rect 30515 24800 30527 24803
rect 30650 24800 30656 24812
rect 30515 24772 30656 24800
rect 30515 24769 30527 24772
rect 30469 24763 30527 24769
rect 30650 24760 30656 24772
rect 30708 24760 30714 24812
rect 30834 24760 30840 24812
rect 30892 24800 30898 24812
rect 31312 24809 31340 24908
rect 31680 24868 31708 24908
rect 33318 24896 33324 24948
rect 33376 24936 33382 24948
rect 36722 24936 36728 24948
rect 33376 24908 36728 24936
rect 33376 24896 33382 24908
rect 36722 24896 36728 24908
rect 36780 24896 36786 24948
rect 40034 24896 40040 24948
rect 40092 24896 40098 24948
rect 34146 24868 34152 24880
rect 31404 24840 31616 24868
rect 31680 24840 34152 24868
rect 31297 24803 31355 24809
rect 31297 24800 31309 24803
rect 30892 24772 31309 24800
rect 30892 24760 30898 24772
rect 31297 24769 31309 24772
rect 31343 24769 31355 24803
rect 31297 24763 31355 24769
rect 28902 24732 28908 24744
rect 28368 24704 28908 24732
rect 28902 24692 28908 24704
rect 28960 24692 28966 24744
rect 30282 24692 30288 24744
rect 30340 24692 30346 24744
rect 30653 24667 30711 24673
rect 30653 24633 30665 24667
rect 30699 24664 30711 24667
rect 31404 24664 31432 24840
rect 31588 24809 31616 24840
rect 34146 24828 34152 24840
rect 34204 24828 34210 24880
rect 38838 24828 38844 24880
rect 38896 24828 38902 24880
rect 39071 24837 39129 24843
rect 39071 24834 39083 24837
rect 38948 24812 39083 24834
rect 31481 24803 31539 24809
rect 31481 24769 31493 24803
rect 31527 24769 31539 24803
rect 31481 24763 31539 24769
rect 31573 24803 31631 24809
rect 31573 24769 31585 24803
rect 31619 24769 31631 24803
rect 31573 24763 31631 24769
rect 31665 24803 31723 24809
rect 31665 24769 31677 24803
rect 31711 24800 31723 24803
rect 31754 24800 31760 24812
rect 31711 24772 31760 24800
rect 31711 24769 31723 24772
rect 31665 24763 31723 24769
rect 31496 24732 31524 24763
rect 31754 24760 31760 24772
rect 31812 24760 31818 24812
rect 35161 24803 35219 24809
rect 35161 24769 35173 24803
rect 35207 24769 35219 24803
rect 35161 24763 35219 24769
rect 31846 24732 31852 24744
rect 31496 24704 31852 24732
rect 31846 24692 31852 24704
rect 31904 24732 31910 24744
rect 32950 24732 32956 24744
rect 31904 24704 32956 24732
rect 31904 24692 31910 24704
rect 32950 24692 32956 24704
rect 33008 24692 33014 24744
rect 35176 24732 35204 24763
rect 35250 24760 35256 24812
rect 35308 24760 35314 24812
rect 35342 24760 35348 24812
rect 35400 24800 35406 24812
rect 35437 24803 35495 24809
rect 35437 24800 35449 24803
rect 35400 24772 35449 24800
rect 35400 24760 35406 24772
rect 35437 24769 35449 24772
rect 35483 24769 35495 24803
rect 35437 24763 35495 24769
rect 35621 24803 35679 24809
rect 35621 24769 35633 24803
rect 35667 24800 35679 24803
rect 37458 24800 37464 24812
rect 35667 24772 37464 24800
rect 35667 24769 35679 24772
rect 35621 24763 35679 24769
rect 37458 24760 37464 24772
rect 37516 24760 37522 24812
rect 37734 24760 37740 24812
rect 37792 24760 37798 24812
rect 38010 24760 38016 24812
rect 38068 24800 38074 24812
rect 38286 24800 38292 24812
rect 38068 24772 38292 24800
rect 38068 24760 38074 24772
rect 38286 24760 38292 24772
rect 38344 24800 38350 24812
rect 38381 24803 38439 24809
rect 38381 24800 38393 24803
rect 38344 24772 38393 24800
rect 38344 24760 38350 24772
rect 38381 24769 38393 24772
rect 38427 24769 38439 24803
rect 38381 24763 38439 24769
rect 38565 24803 38623 24809
rect 38565 24769 38577 24803
rect 38611 24769 38623 24803
rect 38565 24763 38623 24769
rect 35176 24704 35388 24732
rect 35360 24676 35388 24704
rect 36630 24692 36636 24744
rect 36688 24732 36694 24744
rect 36814 24732 36820 24744
rect 36688 24704 36820 24732
rect 36688 24692 36694 24704
rect 36814 24692 36820 24704
rect 36872 24692 36878 24744
rect 37645 24735 37703 24741
rect 37645 24701 37657 24735
rect 37691 24732 37703 24735
rect 37918 24732 37924 24744
rect 37691 24704 37924 24732
rect 37691 24701 37703 24704
rect 37645 24695 37703 24701
rect 37918 24692 37924 24704
rect 37976 24692 37982 24744
rect 38194 24692 38200 24744
rect 38252 24732 38258 24744
rect 38580 24732 38608 24763
rect 38930 24760 38936 24812
rect 38988 24806 39083 24812
rect 38988 24760 38994 24806
rect 39071 24803 39083 24806
rect 39117 24803 39129 24837
rect 39071 24797 39129 24803
rect 40218 24760 40224 24812
rect 40276 24760 40282 24812
rect 38252 24704 38608 24732
rect 38252 24692 38258 24704
rect 31938 24664 31944 24676
rect 30699 24636 31944 24664
rect 30699 24633 30711 24636
rect 30653 24627 30711 24633
rect 31938 24624 31944 24636
rect 31996 24624 32002 24676
rect 35342 24624 35348 24676
rect 35400 24624 35406 24676
rect 36998 24624 37004 24676
rect 37056 24664 37062 24676
rect 37056 24636 37504 24664
rect 37056 24624 37062 24636
rect 27338 24596 27344 24608
rect 26804 24568 27344 24596
rect 27338 24556 27344 24568
rect 27396 24556 27402 24608
rect 27522 24556 27528 24608
rect 27580 24556 27586 24608
rect 27982 24556 27988 24608
rect 28040 24556 28046 24608
rect 28166 24556 28172 24608
rect 28224 24556 28230 24608
rect 28442 24556 28448 24608
rect 28500 24596 28506 24608
rect 28721 24599 28779 24605
rect 28721 24596 28733 24599
rect 28500 24568 28733 24596
rect 28500 24556 28506 24568
rect 28721 24565 28733 24568
rect 28767 24565 28779 24599
rect 28721 24559 28779 24565
rect 31849 24599 31907 24605
rect 31849 24565 31861 24599
rect 31895 24596 31907 24599
rect 33134 24596 33140 24608
rect 31895 24568 33140 24596
rect 31895 24565 31907 24568
rect 31849 24559 31907 24565
rect 33134 24556 33140 24568
rect 33192 24556 33198 24608
rect 37274 24556 37280 24608
rect 37332 24556 37338 24608
rect 37476 24605 37504 24636
rect 37461 24599 37519 24605
rect 37461 24565 37473 24599
rect 37507 24565 37519 24599
rect 38580 24596 38608 24704
rect 38749 24735 38807 24741
rect 38749 24701 38761 24735
rect 38795 24732 38807 24735
rect 39114 24732 39120 24744
rect 38795 24704 39120 24732
rect 38795 24701 38807 24704
rect 38749 24695 38807 24701
rect 39114 24692 39120 24704
rect 39172 24692 39178 24744
rect 39025 24599 39083 24605
rect 39025 24596 39037 24599
rect 38580 24568 39037 24596
rect 37461 24559 37519 24565
rect 39025 24565 39037 24568
rect 39071 24565 39083 24599
rect 39025 24559 39083 24565
rect 39209 24599 39267 24605
rect 39209 24565 39221 24599
rect 39255 24596 39267 24599
rect 39390 24596 39396 24608
rect 39255 24568 39396 24596
rect 39255 24565 39267 24568
rect 39209 24559 39267 24565
rect 39390 24556 39396 24568
rect 39448 24556 39454 24608
rect 1104 24506 40572 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 40572 24506
rect 1104 24432 40572 24454
rect 3145 24395 3203 24401
rect 3145 24361 3157 24395
rect 3191 24392 3203 24395
rect 3878 24392 3884 24404
rect 3191 24364 3884 24392
rect 3191 24361 3203 24364
rect 3145 24355 3203 24361
rect 3878 24352 3884 24364
rect 3936 24352 3942 24404
rect 6917 24395 6975 24401
rect 6288 24364 6868 24392
rect 1397 24259 1455 24265
rect 1397 24225 1409 24259
rect 1443 24256 1455 24259
rect 2866 24256 2872 24268
rect 1443 24228 2872 24256
rect 1443 24225 1455 24228
rect 1397 24219 1455 24225
rect 2866 24216 2872 24228
rect 2924 24256 2930 24268
rect 3694 24256 3700 24268
rect 2924 24228 3700 24256
rect 2924 24216 2930 24228
rect 3694 24216 3700 24228
rect 3752 24256 3758 24268
rect 3789 24259 3847 24265
rect 3789 24256 3801 24259
rect 3752 24228 3801 24256
rect 3752 24216 3758 24228
rect 3789 24225 3801 24228
rect 3835 24225 3847 24259
rect 3789 24219 3847 24225
rect 5537 24259 5595 24265
rect 5537 24225 5549 24259
rect 5583 24256 5595 24259
rect 5718 24256 5724 24268
rect 5583 24228 5724 24256
rect 5583 24225 5595 24228
rect 5537 24219 5595 24225
rect 5718 24216 5724 24228
rect 5776 24256 5782 24268
rect 6181 24259 6239 24265
rect 6181 24256 6193 24259
rect 5776 24228 6193 24256
rect 5776 24216 5782 24228
rect 6181 24225 6193 24228
rect 6227 24256 6239 24259
rect 6288 24256 6316 24364
rect 6840 24336 6868 24364
rect 6917 24361 6929 24395
rect 6963 24392 6975 24395
rect 8018 24392 8024 24404
rect 6963 24364 8024 24392
rect 6963 24361 6975 24364
rect 6917 24355 6975 24361
rect 8018 24352 8024 24364
rect 8076 24352 8082 24404
rect 8110 24352 8116 24404
rect 8168 24392 8174 24404
rect 9585 24395 9643 24401
rect 9585 24392 9597 24395
rect 8168 24364 9597 24392
rect 8168 24352 8174 24364
rect 9585 24361 9597 24364
rect 9631 24361 9643 24395
rect 9585 24355 9643 24361
rect 9674 24352 9680 24404
rect 9732 24392 9738 24404
rect 13630 24392 13636 24404
rect 9732 24364 13636 24392
rect 9732 24352 9738 24364
rect 13630 24352 13636 24364
rect 13688 24352 13694 24404
rect 14458 24352 14464 24404
rect 14516 24392 14522 24404
rect 14737 24395 14795 24401
rect 14737 24392 14749 24395
rect 14516 24364 14749 24392
rect 14516 24352 14522 24364
rect 14737 24361 14749 24364
rect 14783 24361 14795 24395
rect 15654 24392 15660 24404
rect 14737 24355 14795 24361
rect 15304 24364 15660 24392
rect 6362 24284 6368 24336
rect 6420 24324 6426 24336
rect 6420 24296 6776 24324
rect 6420 24284 6426 24296
rect 6227 24228 6316 24256
rect 6472 24228 6684 24256
rect 6227 24225 6239 24228
rect 6181 24219 6239 24225
rect 3142 24188 3148 24200
rect 2806 24160 3148 24188
rect 3142 24148 3148 24160
rect 3200 24148 3206 24200
rect 6270 24148 6276 24200
rect 6328 24188 6334 24200
rect 6365 24191 6423 24197
rect 6365 24188 6377 24191
rect 6328 24160 6377 24188
rect 6328 24148 6334 24160
rect 6365 24157 6377 24160
rect 6411 24157 6423 24191
rect 6365 24151 6423 24157
rect 1670 24080 1676 24132
rect 1728 24080 1734 24132
rect 4062 24080 4068 24132
rect 4120 24080 4126 24132
rect 4614 24080 4620 24132
rect 4672 24080 4678 24132
rect 5994 24080 6000 24132
rect 6052 24120 6058 24132
rect 6472 24120 6500 24228
rect 6546 24148 6552 24200
rect 6604 24148 6610 24200
rect 6656 24197 6684 24228
rect 6748 24197 6776 24296
rect 6822 24284 6828 24336
rect 6880 24284 6886 24336
rect 7650 24284 7656 24336
rect 7708 24324 7714 24336
rect 7834 24324 7840 24336
rect 7708 24296 7840 24324
rect 7708 24284 7714 24296
rect 7834 24284 7840 24296
rect 7892 24284 7898 24336
rect 8294 24284 8300 24336
rect 8352 24324 8358 24336
rect 8352 24296 8616 24324
rect 8352 24284 8358 24296
rect 6641 24191 6699 24197
rect 6641 24157 6653 24191
rect 6687 24157 6699 24191
rect 6641 24151 6699 24157
rect 6733 24191 6791 24197
rect 6733 24157 6745 24191
rect 6779 24157 6791 24191
rect 6733 24151 6791 24157
rect 7834 24148 7840 24200
rect 7892 24188 7898 24200
rect 8501 24197 8529 24296
rect 8588 24256 8616 24296
rect 9030 24284 9036 24336
rect 9088 24324 9094 24336
rect 9088 24296 9260 24324
rect 9088 24284 9094 24296
rect 9232 24256 9260 24296
rect 9306 24284 9312 24336
rect 9364 24324 9370 24336
rect 14918 24324 14924 24336
rect 9364 24296 9674 24324
rect 9364 24284 9370 24296
rect 9646 24256 9674 24296
rect 14471 24296 14924 24324
rect 10870 24256 10876 24268
rect 8588 24228 9076 24256
rect 9232 24228 9449 24256
rect 9646 24228 10876 24256
rect 9048 24197 9076 24228
rect 8021 24191 8079 24197
rect 8021 24188 8033 24191
rect 7892 24160 8033 24188
rect 7892 24148 7898 24160
rect 8021 24157 8033 24160
rect 8067 24157 8079 24191
rect 8021 24151 8079 24157
rect 8114 24191 8172 24197
rect 8114 24157 8126 24191
rect 8160 24157 8172 24191
rect 8114 24151 8172 24157
rect 8297 24191 8355 24197
rect 8297 24157 8309 24191
rect 8343 24157 8355 24191
rect 8501 24191 8563 24197
rect 8501 24160 8517 24191
rect 8297 24151 8355 24157
rect 8505 24157 8517 24160
rect 8551 24157 8563 24191
rect 8929 24191 8987 24197
rect 8929 24188 8941 24191
rect 8505 24151 8563 24157
rect 8772 24160 8941 24188
rect 6052 24092 6500 24120
rect 6052 24080 6058 24092
rect 5626 24012 5632 24064
rect 5684 24012 5690 24064
rect 6564 24052 6592 24148
rect 7374 24080 7380 24132
rect 7432 24120 7438 24132
rect 8128 24120 8156 24151
rect 8312 24120 8340 24151
rect 7432 24092 8156 24120
rect 8184 24092 8340 24120
rect 7432 24080 7438 24092
rect 8184 24052 8212 24092
rect 8386 24080 8392 24132
rect 8444 24080 8450 24132
rect 8772 24120 8800 24160
rect 8929 24157 8941 24160
rect 8975 24157 8987 24191
rect 8929 24151 8987 24157
rect 9034 24191 9092 24197
rect 9034 24157 9046 24191
rect 9080 24157 9092 24191
rect 9034 24151 9092 24157
rect 8588 24092 8800 24120
rect 8588 24064 8616 24092
rect 6564 24024 8212 24052
rect 8570 24012 8576 24064
rect 8628 24012 8634 24064
rect 8662 24012 8668 24064
rect 8720 24012 8726 24064
rect 9048 24052 9076 24151
rect 9214 24148 9220 24200
rect 9272 24148 9278 24200
rect 9421 24197 9449 24228
rect 10870 24216 10876 24228
rect 10928 24216 10934 24268
rect 11330 24216 11336 24268
rect 11388 24256 11394 24268
rect 14471 24256 14499 24296
rect 14918 24284 14924 24296
rect 14976 24284 14982 24336
rect 15304 24333 15332 24364
rect 15654 24352 15660 24364
rect 15712 24352 15718 24404
rect 17310 24352 17316 24404
rect 17368 24392 17374 24404
rect 17773 24395 17831 24401
rect 17773 24392 17785 24395
rect 17368 24364 17785 24392
rect 17368 24352 17374 24364
rect 17773 24361 17785 24364
rect 17819 24361 17831 24395
rect 17773 24355 17831 24361
rect 19981 24395 20039 24401
rect 19981 24361 19993 24395
rect 20027 24392 20039 24395
rect 20349 24395 20407 24401
rect 20349 24392 20361 24395
rect 20027 24364 20361 24392
rect 20027 24361 20039 24364
rect 19981 24355 20039 24361
rect 20349 24361 20361 24364
rect 20395 24361 20407 24395
rect 20349 24355 20407 24361
rect 23400 24364 23796 24392
rect 15105 24327 15163 24333
rect 15105 24293 15117 24327
rect 15151 24293 15163 24327
rect 15105 24287 15163 24293
rect 15289 24327 15347 24333
rect 15289 24293 15301 24327
rect 15335 24293 15347 24327
rect 15289 24287 15347 24293
rect 11388 24228 14499 24256
rect 11388 24216 11394 24228
rect 9406 24191 9464 24197
rect 9406 24157 9418 24191
rect 9452 24157 9464 24191
rect 9406 24151 9464 24157
rect 10410 24148 10416 24200
rect 10468 24188 10474 24200
rect 10594 24188 10600 24200
rect 10468 24160 10600 24188
rect 10468 24148 10474 24160
rect 10594 24148 10600 24160
rect 10652 24188 10658 24200
rect 10965 24191 11023 24197
rect 10965 24188 10977 24191
rect 10652 24160 10977 24188
rect 10652 24148 10658 24160
rect 10965 24157 10977 24160
rect 11011 24157 11023 24191
rect 10965 24151 11023 24157
rect 11149 24191 11207 24197
rect 11149 24157 11161 24191
rect 11195 24188 11207 24191
rect 11238 24188 11244 24200
rect 11195 24160 11244 24188
rect 11195 24157 11207 24160
rect 11149 24151 11207 24157
rect 11238 24148 11244 24160
rect 11296 24188 11302 24200
rect 12618 24188 12624 24200
rect 11296 24160 12624 24188
rect 11296 24148 11302 24160
rect 12618 24148 12624 24160
rect 12676 24148 12682 24200
rect 13906 24148 13912 24200
rect 13964 24188 13970 24200
rect 14471 24197 14499 24228
rect 14734 24216 14740 24268
rect 14792 24256 14798 24268
rect 15120 24256 15148 24287
rect 15470 24284 15476 24336
rect 15528 24284 15534 24336
rect 15746 24284 15752 24336
rect 15804 24284 15810 24336
rect 18966 24284 18972 24336
rect 19024 24324 19030 24336
rect 19886 24324 19892 24336
rect 19024 24296 19892 24324
rect 19024 24284 19030 24296
rect 19886 24284 19892 24296
rect 19944 24284 19950 24336
rect 20441 24327 20499 24333
rect 20441 24293 20453 24327
rect 20487 24324 20499 24327
rect 20898 24324 20904 24336
rect 20487 24296 20904 24324
rect 20487 24293 20499 24296
rect 20441 24287 20499 24293
rect 20898 24284 20904 24296
rect 20956 24284 20962 24336
rect 14792 24228 15148 24256
rect 15488 24256 15516 24284
rect 15565 24259 15623 24265
rect 15565 24256 15577 24259
rect 15488 24228 15577 24256
rect 14792 24216 14798 24228
rect 15565 24225 15577 24228
rect 15611 24225 15623 24259
rect 15565 24219 15623 24225
rect 16298 24216 16304 24268
rect 16356 24256 16362 24268
rect 16577 24259 16635 24265
rect 16577 24256 16589 24259
rect 16356 24228 16589 24256
rect 16356 24216 16362 24228
rect 16577 24225 16589 24228
rect 16623 24225 16635 24259
rect 16577 24219 16635 24225
rect 18509 24259 18567 24265
rect 18509 24225 18521 24259
rect 18555 24256 18567 24259
rect 18598 24256 18604 24268
rect 18555 24228 18604 24256
rect 18555 24225 18567 24228
rect 18509 24219 18567 24225
rect 18598 24216 18604 24228
rect 18656 24256 18662 24268
rect 19518 24256 19524 24268
rect 18656 24228 19524 24256
rect 18656 24216 18662 24228
rect 19518 24216 19524 24228
rect 19576 24216 19582 24268
rect 20070 24216 20076 24268
rect 20128 24256 20134 24268
rect 20257 24259 20315 24265
rect 20257 24256 20269 24259
rect 20128 24228 20269 24256
rect 20128 24216 20134 24228
rect 20257 24225 20269 24228
rect 20303 24256 20315 24259
rect 20303 24228 23208 24256
rect 20303 24225 20315 24228
rect 20257 24219 20315 24225
rect 14093 24191 14151 24197
rect 14093 24188 14105 24191
rect 13964 24160 14105 24188
rect 13964 24148 13970 24160
rect 14093 24157 14105 24160
rect 14139 24157 14151 24191
rect 14093 24151 14151 24157
rect 14369 24191 14427 24197
rect 14369 24157 14381 24191
rect 14415 24157 14427 24191
rect 14369 24151 14427 24157
rect 14460 24191 14518 24197
rect 14460 24157 14472 24191
rect 14506 24157 14518 24191
rect 14460 24151 14518 24157
rect 9306 24080 9312 24132
rect 9364 24080 9370 24132
rect 12250 24120 12256 24132
rect 9416 24092 12256 24120
rect 9416 24052 9444 24092
rect 12250 24080 12256 24092
rect 12308 24080 12314 24132
rect 14251 24123 14309 24129
rect 14251 24120 14263 24123
rect 12406 24092 14263 24120
rect 9048 24024 9444 24052
rect 10870 24012 10876 24064
rect 10928 24052 10934 24064
rect 12406 24052 12434 24092
rect 14251 24089 14263 24092
rect 14297 24120 14309 24123
rect 14384 24120 14412 24151
rect 14550 24148 14556 24200
rect 14608 24148 14614 24200
rect 15286 24188 15292 24200
rect 14844 24160 15292 24188
rect 14844 24120 14872 24160
rect 15286 24148 15292 24160
rect 15344 24148 15350 24200
rect 15470 24148 15476 24200
rect 15528 24188 15534 24200
rect 15749 24191 15807 24197
rect 15749 24188 15761 24191
rect 15528 24160 15761 24188
rect 15528 24148 15534 24160
rect 15749 24157 15761 24160
rect 15795 24157 15807 24191
rect 15749 24151 15807 24157
rect 16025 24191 16083 24197
rect 16025 24157 16037 24191
rect 16071 24188 16083 24191
rect 16071 24160 16344 24188
rect 16071 24157 16083 24160
rect 16025 24151 16083 24157
rect 14297 24089 14320 24120
rect 14384 24092 14872 24120
rect 14251 24083 14320 24089
rect 10928 24024 12434 24052
rect 14292 24052 14320 24083
rect 14918 24080 14924 24132
rect 14976 24120 14982 24132
rect 16209 24123 16267 24129
rect 16209 24120 16221 24123
rect 14976 24092 16221 24120
rect 14976 24080 14982 24092
rect 16209 24089 16221 24092
rect 16255 24089 16267 24123
rect 16316 24120 16344 24160
rect 16390 24148 16396 24200
rect 16448 24148 16454 24200
rect 17954 24148 17960 24200
rect 18012 24148 18018 24200
rect 18141 24191 18199 24197
rect 18141 24157 18153 24191
rect 18187 24157 18199 24191
rect 18141 24151 18199 24157
rect 18233 24191 18291 24197
rect 18233 24157 18245 24191
rect 18279 24188 18291 24191
rect 19150 24188 19156 24200
rect 18279 24160 19156 24188
rect 18279 24157 18291 24160
rect 18233 24151 18291 24157
rect 17034 24120 17040 24132
rect 16316 24092 17040 24120
rect 16209 24083 16267 24089
rect 17034 24080 17040 24092
rect 17092 24080 17098 24132
rect 18156 24120 18184 24151
rect 19150 24148 19156 24160
rect 19208 24188 19214 24200
rect 19613 24191 19671 24197
rect 19613 24188 19625 24191
rect 19208 24160 19625 24188
rect 19208 24148 19214 24160
rect 19613 24157 19625 24160
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 18414 24120 18420 24132
rect 18156 24092 18420 24120
rect 18414 24080 18420 24092
rect 18472 24080 18478 24132
rect 18506 24080 18512 24132
rect 18564 24120 18570 24132
rect 18693 24123 18751 24129
rect 18693 24120 18705 24123
rect 18564 24092 18705 24120
rect 18564 24080 18570 24092
rect 18693 24089 18705 24092
rect 18739 24089 18751 24123
rect 18693 24083 18751 24089
rect 18877 24123 18935 24129
rect 18877 24089 18889 24123
rect 18923 24120 18935 24123
rect 20088 24120 20116 24216
rect 20533 24191 20591 24197
rect 20533 24157 20545 24191
rect 20579 24188 20591 24191
rect 20622 24188 20628 24200
rect 20579 24160 20628 24188
rect 20579 24157 20591 24160
rect 20533 24151 20591 24157
rect 20622 24148 20628 24160
rect 20680 24148 20686 24200
rect 23014 24148 23020 24200
rect 23072 24148 23078 24200
rect 23180 24197 23208 24228
rect 23165 24191 23223 24197
rect 23165 24157 23177 24191
rect 23211 24188 23223 24191
rect 23400 24188 23428 24364
rect 23661 24327 23719 24333
rect 23661 24293 23673 24327
rect 23707 24293 23719 24327
rect 23768 24324 23796 24364
rect 23842 24352 23848 24404
rect 23900 24352 23906 24404
rect 24118 24352 24124 24404
rect 24176 24352 24182 24404
rect 25590 24392 25596 24404
rect 24412 24364 25596 24392
rect 24412 24324 24440 24364
rect 25590 24352 25596 24364
rect 25648 24352 25654 24404
rect 25866 24352 25872 24404
rect 25924 24392 25930 24404
rect 26145 24395 26203 24401
rect 26145 24392 26157 24395
rect 25924 24364 26157 24392
rect 25924 24352 25930 24364
rect 26145 24361 26157 24364
rect 26191 24361 26203 24395
rect 26145 24355 26203 24361
rect 26605 24395 26663 24401
rect 26605 24361 26617 24395
rect 26651 24392 26663 24395
rect 26694 24392 26700 24404
rect 26651 24364 26700 24392
rect 26651 24361 26663 24364
rect 26605 24355 26663 24361
rect 26694 24352 26700 24364
rect 26752 24352 26758 24404
rect 26970 24352 26976 24404
rect 27028 24392 27034 24404
rect 27249 24395 27307 24401
rect 27249 24392 27261 24395
rect 27028 24364 27261 24392
rect 27028 24352 27034 24364
rect 27249 24361 27261 24364
rect 27295 24361 27307 24395
rect 27249 24355 27307 24361
rect 27338 24352 27344 24404
rect 27396 24392 27402 24404
rect 27396 24364 28120 24392
rect 27396 24352 27402 24364
rect 23768 24296 24440 24324
rect 23661 24287 23719 24293
rect 23676 24256 23704 24287
rect 24412 24268 24440 24296
rect 24949 24327 25007 24333
rect 24949 24293 24961 24327
rect 24995 24324 25007 24327
rect 25130 24324 25136 24336
rect 24995 24296 25136 24324
rect 24995 24293 25007 24296
rect 24949 24287 25007 24293
rect 25130 24284 25136 24296
rect 25188 24284 25194 24336
rect 27522 24284 27528 24336
rect 27580 24284 27586 24336
rect 28092 24324 28120 24364
rect 28350 24352 28356 24404
rect 28408 24392 28414 24404
rect 28813 24395 28871 24401
rect 28813 24392 28825 24395
rect 28408 24364 28825 24392
rect 28408 24352 28414 24364
rect 28813 24361 28825 24364
rect 28859 24361 28871 24395
rect 28813 24355 28871 24361
rect 30926 24352 30932 24404
rect 30984 24392 30990 24404
rect 32490 24392 32496 24404
rect 30984 24364 32496 24392
rect 30984 24352 30990 24364
rect 32490 24352 32496 24364
rect 32548 24352 32554 24404
rect 33502 24352 33508 24404
rect 33560 24392 33566 24404
rect 36078 24392 36084 24404
rect 33560 24364 36084 24392
rect 33560 24352 33566 24364
rect 36078 24352 36084 24364
rect 36136 24352 36142 24404
rect 37918 24352 37924 24404
rect 37976 24352 37982 24404
rect 39482 24392 39488 24404
rect 38396 24364 39488 24392
rect 29273 24327 29331 24333
rect 29273 24324 29285 24327
rect 28092 24296 29285 24324
rect 29273 24293 29285 24296
rect 29319 24293 29331 24327
rect 29273 24287 29331 24293
rect 29638 24284 29644 24336
rect 29696 24324 29702 24336
rect 38396 24324 38424 24364
rect 39482 24352 39488 24364
rect 39540 24352 39546 24404
rect 39666 24352 39672 24404
rect 39724 24392 39730 24404
rect 40037 24395 40095 24401
rect 40037 24392 40049 24395
rect 39724 24364 40049 24392
rect 39724 24352 39730 24364
rect 40037 24361 40049 24364
rect 40083 24361 40095 24395
rect 40037 24355 40095 24361
rect 38562 24324 38568 24336
rect 29696 24296 38424 24324
rect 38488 24296 38568 24324
rect 29696 24284 29702 24296
rect 23676 24228 23796 24256
rect 23211 24160 23428 24188
rect 23211 24157 23223 24160
rect 23165 24151 23223 24157
rect 23474 24148 23480 24200
rect 23532 24197 23538 24200
rect 23532 24188 23540 24197
rect 23532 24160 23577 24188
rect 23532 24151 23540 24160
rect 23532 24148 23538 24151
rect 23658 24148 23664 24200
rect 23716 24148 23722 24200
rect 23768 24197 23796 24228
rect 24394 24216 24400 24268
rect 24452 24256 24458 24268
rect 24489 24259 24547 24265
rect 24489 24256 24501 24259
rect 24452 24228 24501 24256
rect 24452 24216 24458 24228
rect 24489 24225 24501 24228
rect 24535 24225 24547 24259
rect 24489 24219 24547 24225
rect 24762 24216 24768 24268
rect 24820 24256 24826 24268
rect 27246 24256 27252 24268
rect 24820 24228 27252 24256
rect 24820 24216 24826 24228
rect 27246 24216 27252 24228
rect 27304 24216 27310 24268
rect 27540 24256 27568 24284
rect 27448 24228 27568 24256
rect 23753 24191 23811 24197
rect 23753 24157 23765 24191
rect 23799 24157 23811 24191
rect 23753 24151 23811 24157
rect 23842 24148 23848 24200
rect 23900 24188 23906 24200
rect 23937 24191 23995 24197
rect 23937 24188 23949 24191
rect 23900 24160 23949 24188
rect 23900 24148 23906 24160
rect 23937 24157 23949 24160
rect 23983 24188 23995 24191
rect 24670 24188 24676 24200
rect 23983 24160 24676 24188
rect 23983 24157 23995 24160
rect 23937 24151 23995 24157
rect 24670 24148 24676 24160
rect 24728 24148 24734 24200
rect 25130 24148 25136 24200
rect 25188 24188 25194 24200
rect 25225 24191 25283 24197
rect 25225 24188 25237 24191
rect 25188 24160 25237 24188
rect 25188 24148 25194 24160
rect 25225 24157 25237 24160
rect 25271 24157 25283 24191
rect 25225 24151 25283 24157
rect 25685 24191 25743 24197
rect 25685 24157 25697 24191
rect 25731 24188 25743 24191
rect 25866 24188 25872 24200
rect 25731 24160 25872 24188
rect 25731 24157 25743 24160
rect 25685 24151 25743 24157
rect 18923 24092 20116 24120
rect 18923 24089 18935 24092
rect 18877 24083 18935 24089
rect 15930 24052 15936 24064
rect 14292 24024 15936 24052
rect 10928 24012 10934 24024
rect 15930 24012 15936 24024
rect 15988 24012 15994 24064
rect 19978 24012 19984 24064
rect 20036 24012 20042 24064
rect 20070 24012 20076 24064
rect 20128 24052 20134 24064
rect 20165 24055 20223 24061
rect 20165 24052 20177 24055
rect 20128 24024 20177 24052
rect 20128 24012 20134 24024
rect 20165 24021 20177 24024
rect 20211 24021 20223 24055
rect 20640 24052 20668 24148
rect 20898 24080 20904 24132
rect 20956 24120 20962 24132
rect 23293 24123 23351 24129
rect 23293 24120 23305 24123
rect 20956 24092 23305 24120
rect 20956 24080 20962 24092
rect 23293 24089 23305 24092
rect 23339 24089 23351 24123
rect 23293 24083 23351 24089
rect 23385 24123 23443 24129
rect 23385 24089 23397 24123
rect 23431 24120 23443 24123
rect 23676 24120 23704 24148
rect 24210 24120 24216 24132
rect 23431 24092 24216 24120
rect 23431 24089 23443 24092
rect 23385 24083 23443 24089
rect 24210 24080 24216 24092
rect 24268 24080 24274 24132
rect 25240 24120 25268 24151
rect 25866 24148 25872 24160
rect 25924 24148 25930 24200
rect 26145 24191 26203 24197
rect 26145 24157 26157 24191
rect 26191 24188 26203 24191
rect 26694 24188 26700 24200
rect 26191 24160 26700 24188
rect 26191 24157 26203 24160
rect 26145 24151 26203 24157
rect 26694 24148 26700 24160
rect 26752 24148 26758 24200
rect 27448 24197 27476 24228
rect 27982 24216 27988 24268
rect 28040 24256 28046 24268
rect 28040 24228 28212 24256
rect 28040 24216 28046 24228
rect 27433 24191 27491 24197
rect 27433 24157 27445 24191
rect 27479 24157 27491 24191
rect 27433 24151 27491 24157
rect 27522 24148 27528 24200
rect 27580 24148 27586 24200
rect 27706 24148 27712 24200
rect 27764 24148 27770 24200
rect 27801 24191 27859 24197
rect 27801 24157 27813 24191
rect 27847 24157 27859 24191
rect 27801 24151 27859 24157
rect 25774 24120 25780 24132
rect 25240 24092 25780 24120
rect 25774 24080 25780 24092
rect 25832 24120 25838 24132
rect 25961 24123 26019 24129
rect 25961 24120 25973 24123
rect 25832 24092 25973 24120
rect 25832 24080 25838 24092
rect 25961 24089 25973 24092
rect 26007 24089 26019 24123
rect 25961 24083 26019 24089
rect 26237 24123 26295 24129
rect 26237 24089 26249 24123
rect 26283 24089 26295 24123
rect 26237 24083 26295 24089
rect 23474 24052 23480 24064
rect 20640 24024 23480 24052
rect 20165 24015 20223 24021
rect 23474 24012 23480 24024
rect 23532 24052 23538 24064
rect 23658 24052 23664 24064
rect 23532 24024 23664 24052
rect 23532 24012 23538 24024
rect 23658 24012 23664 24024
rect 23716 24012 23722 24064
rect 25866 24012 25872 24064
rect 25924 24052 25930 24064
rect 26252 24052 26280 24083
rect 26418 24080 26424 24132
rect 26476 24080 26482 24132
rect 27430 24052 27436 24064
rect 25924 24024 27436 24052
rect 25924 24012 25930 24024
rect 27430 24012 27436 24024
rect 27488 24012 27494 24064
rect 27522 24012 27528 24064
rect 27580 24052 27586 24064
rect 27816 24052 27844 24151
rect 28074 24148 28080 24200
rect 28132 24148 28138 24200
rect 28184 24197 28212 24228
rect 28718 24216 28724 24268
rect 28776 24256 28782 24268
rect 28776 24228 29132 24256
rect 28776 24216 28782 24228
rect 28170 24191 28228 24197
rect 28170 24157 28182 24191
rect 28216 24157 28228 24191
rect 28170 24151 28228 24157
rect 28442 24148 28448 24200
rect 28500 24148 28506 24200
rect 28534 24148 28540 24200
rect 28592 24197 28598 24200
rect 28592 24188 28600 24197
rect 28592 24160 28637 24188
rect 28592 24151 28600 24160
rect 28592 24148 28598 24151
rect 28994 24148 29000 24200
rect 29052 24148 29058 24200
rect 29104 24197 29132 24228
rect 37826 24216 37832 24268
rect 37884 24256 37890 24268
rect 37884 24228 38332 24256
rect 37884 24216 37890 24228
rect 29089 24191 29147 24197
rect 29089 24157 29101 24191
rect 29135 24157 29147 24191
rect 29089 24151 29147 24157
rect 36538 24148 36544 24200
rect 36596 24188 36602 24200
rect 38304 24197 38332 24228
rect 38488 24197 38516 24296
rect 38562 24284 38568 24296
rect 38620 24284 38626 24336
rect 38105 24191 38163 24197
rect 38105 24188 38117 24191
rect 36596 24160 38117 24188
rect 36596 24148 36602 24160
rect 38105 24157 38117 24160
rect 38151 24157 38163 24191
rect 38105 24151 38163 24157
rect 38289 24191 38347 24197
rect 38289 24157 38301 24191
rect 38335 24157 38347 24191
rect 38289 24151 38347 24157
rect 38473 24191 38531 24197
rect 38473 24157 38485 24191
rect 38519 24157 38531 24191
rect 38473 24151 38531 24157
rect 38565 24191 38623 24197
rect 38565 24157 38577 24191
rect 38611 24188 38623 24191
rect 39390 24188 39396 24200
rect 38611 24160 39396 24188
rect 38611 24157 38623 24160
rect 38565 24151 38623 24157
rect 39390 24148 39396 24160
rect 39448 24148 39454 24200
rect 39666 24148 39672 24200
rect 39724 24148 39730 24200
rect 40126 24148 40132 24200
rect 40184 24188 40190 24200
rect 40221 24191 40279 24197
rect 40221 24188 40233 24191
rect 40184 24160 40233 24188
rect 40184 24148 40190 24160
rect 40221 24157 40233 24160
rect 40267 24157 40279 24191
rect 40221 24151 40279 24157
rect 28353 24123 28411 24129
rect 28353 24089 28365 24123
rect 28399 24120 28411 24123
rect 28626 24120 28632 24132
rect 28399 24092 28632 24120
rect 28399 24089 28411 24092
rect 28353 24083 28411 24089
rect 28626 24080 28632 24092
rect 28684 24080 28690 24132
rect 28813 24123 28871 24129
rect 28813 24089 28825 24123
rect 28859 24089 28871 24123
rect 28813 24083 28871 24089
rect 27580 24024 27844 24052
rect 28721 24055 28779 24061
rect 27580 24012 27586 24024
rect 28721 24021 28733 24055
rect 28767 24052 28779 24055
rect 28828 24052 28856 24083
rect 38194 24080 38200 24132
rect 38252 24080 38258 24132
rect 28767 24024 28856 24052
rect 28767 24021 28779 24024
rect 28721 24015 28779 24021
rect 31110 24012 31116 24064
rect 31168 24052 31174 24064
rect 35342 24052 35348 24064
rect 31168 24024 35348 24052
rect 31168 24012 31174 24024
rect 35342 24012 35348 24024
rect 35400 24012 35406 24064
rect 37090 24012 37096 24064
rect 37148 24052 37154 24064
rect 39485 24055 39543 24061
rect 39485 24052 39497 24055
rect 37148 24024 39497 24052
rect 37148 24012 37154 24024
rect 39485 24021 39497 24024
rect 39531 24021 39543 24055
rect 39485 24015 39543 24021
rect 1104 23962 40572 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 40572 23962
rect 1104 23888 40572 23910
rect 1670 23808 1676 23860
rect 1728 23848 1734 23860
rect 2501 23851 2559 23857
rect 2501 23848 2513 23851
rect 1728 23820 2513 23848
rect 1728 23808 1734 23820
rect 2501 23817 2513 23820
rect 2547 23817 2559 23851
rect 2501 23811 2559 23817
rect 2869 23851 2927 23857
rect 2869 23817 2881 23851
rect 2915 23848 2927 23851
rect 2958 23848 2964 23860
rect 2915 23820 2964 23848
rect 2915 23817 2927 23820
rect 2869 23811 2927 23817
rect 2958 23808 2964 23820
rect 3016 23808 3022 23860
rect 4985 23851 5043 23857
rect 4985 23817 4997 23851
rect 5031 23848 5043 23851
rect 5626 23848 5632 23860
rect 5031 23820 5632 23848
rect 5031 23817 5043 23820
rect 4985 23811 5043 23817
rect 5626 23808 5632 23820
rect 5684 23808 5690 23860
rect 5994 23848 6000 23860
rect 5920 23820 6000 23848
rect 3694 23740 3700 23792
rect 3752 23740 3758 23792
rect 4525 23783 4583 23789
rect 4525 23749 4537 23783
rect 4571 23780 4583 23783
rect 4614 23780 4620 23792
rect 4571 23752 4620 23780
rect 4571 23749 4583 23752
rect 4525 23743 4583 23749
rect 4614 23740 4620 23752
rect 4672 23780 4678 23792
rect 5442 23780 5448 23792
rect 4672 23752 5448 23780
rect 4672 23740 4678 23752
rect 5442 23740 5448 23752
rect 5500 23740 5506 23792
rect 5920 23789 5948 23820
rect 5994 23808 6000 23820
rect 6052 23808 6058 23860
rect 6730 23808 6736 23860
rect 6788 23808 6794 23860
rect 7834 23808 7840 23860
rect 7892 23808 7898 23860
rect 10410 23848 10416 23860
rect 8312 23820 10416 23848
rect 5905 23783 5963 23789
rect 5905 23780 5917 23783
rect 5552 23752 5917 23780
rect 2961 23715 3019 23721
rect 2961 23681 2973 23715
rect 3007 23712 3019 23715
rect 3050 23712 3056 23724
rect 3007 23684 3056 23712
rect 3007 23681 3019 23684
rect 2961 23675 3019 23681
rect 3050 23672 3056 23684
rect 3108 23672 3114 23724
rect 3878 23672 3884 23724
rect 3936 23712 3942 23724
rect 5552 23712 5580 23752
rect 5905 23749 5917 23752
rect 5951 23749 5963 23783
rect 5905 23743 5963 23749
rect 6641 23783 6699 23789
rect 6641 23749 6653 23783
rect 6687 23780 6699 23783
rect 6748 23780 6776 23808
rect 6687 23752 6776 23780
rect 6687 23749 6699 23752
rect 6641 23743 6699 23749
rect 6822 23740 6828 23792
rect 6880 23780 6886 23792
rect 8113 23783 8171 23789
rect 8113 23780 8125 23783
rect 6880 23752 8125 23780
rect 6880 23740 6886 23752
rect 8113 23749 8125 23752
rect 8159 23749 8171 23783
rect 8113 23743 8171 23749
rect 3936 23684 5580 23712
rect 5813 23715 5871 23721
rect 3936 23672 3942 23684
rect 5813 23681 5825 23715
rect 5859 23712 5871 23715
rect 5997 23715 6055 23721
rect 5859 23684 5948 23712
rect 5859 23681 5871 23684
rect 5813 23675 5871 23681
rect 3145 23647 3203 23653
rect 3145 23613 3157 23647
rect 3191 23644 3203 23647
rect 3191 23616 5028 23644
rect 3191 23613 3203 23616
rect 3145 23607 3203 23613
rect 4062 23536 4068 23588
rect 4120 23576 4126 23588
rect 4617 23579 4675 23585
rect 4617 23576 4629 23579
rect 4120 23548 4629 23576
rect 4120 23536 4126 23548
rect 4617 23545 4629 23548
rect 4663 23545 4675 23579
rect 5000 23576 5028 23616
rect 5074 23604 5080 23656
rect 5132 23604 5138 23656
rect 5258 23604 5264 23656
rect 5316 23604 5322 23656
rect 5534 23604 5540 23656
rect 5592 23644 5598 23656
rect 5920 23644 5948 23684
rect 5997 23681 6009 23715
rect 6043 23681 6055 23715
rect 5997 23675 6055 23681
rect 5592 23616 5948 23644
rect 6012 23644 6040 23675
rect 6178 23672 6184 23724
rect 6236 23672 6242 23724
rect 6270 23672 6276 23724
rect 6328 23712 6334 23724
rect 6546 23712 6552 23724
rect 6328 23684 6552 23712
rect 6328 23672 6334 23684
rect 6546 23672 6552 23684
rect 6604 23672 6610 23724
rect 6733 23715 6791 23721
rect 6733 23712 6745 23715
rect 6656 23684 6745 23712
rect 6656 23644 6684 23684
rect 6733 23681 6745 23684
rect 6779 23681 6791 23715
rect 6733 23675 6791 23681
rect 6917 23715 6975 23721
rect 6917 23681 6929 23715
rect 6963 23712 6975 23715
rect 7374 23712 7380 23724
rect 6963 23684 7380 23712
rect 6963 23681 6975 23684
rect 6917 23675 6975 23681
rect 7374 23672 7380 23684
rect 7432 23672 7438 23724
rect 7926 23672 7932 23724
rect 7984 23721 7990 23724
rect 7984 23715 8033 23721
rect 7984 23681 7987 23715
rect 8021 23681 8033 23715
rect 7984 23675 8033 23681
rect 7984 23672 7990 23675
rect 8202 23672 8208 23724
rect 8260 23712 8266 23724
rect 8312 23712 8340 23820
rect 10410 23808 10416 23820
rect 10468 23808 10474 23860
rect 10502 23808 10508 23860
rect 10560 23848 10566 23860
rect 10560 23820 11376 23848
rect 10560 23808 10566 23820
rect 11054 23780 11060 23792
rect 8588 23752 11060 23780
rect 8260 23684 8340 23712
rect 8388 23715 8446 23721
rect 8260 23672 8266 23684
rect 8388 23681 8400 23715
rect 8434 23681 8446 23715
rect 8388 23675 8446 23681
rect 8474 23715 8532 23721
rect 8474 23681 8486 23715
rect 8520 23713 8532 23715
rect 8588 23713 8616 23752
rect 11054 23740 11060 23752
rect 11112 23740 11118 23792
rect 11348 23789 11376 23820
rect 18414 23808 18420 23860
rect 18472 23848 18478 23860
rect 18601 23851 18659 23857
rect 18601 23848 18613 23851
rect 18472 23820 18613 23848
rect 18472 23808 18478 23820
rect 18601 23817 18613 23820
rect 18647 23817 18659 23851
rect 18601 23811 18659 23817
rect 19150 23808 19156 23860
rect 19208 23808 19214 23860
rect 19886 23848 19892 23860
rect 19352 23820 19892 23848
rect 11333 23783 11391 23789
rect 11333 23749 11345 23783
rect 11379 23749 11391 23783
rect 18046 23780 18052 23792
rect 11333 23743 11391 23749
rect 16684 23752 18052 23780
rect 8520 23685 8616 23713
rect 8520 23681 8532 23685
rect 8474 23675 8532 23681
rect 6012 23616 6684 23644
rect 5592 23604 5598 23616
rect 5276 23576 5304 23604
rect 5000 23548 5304 23576
rect 5920 23576 5948 23616
rect 6528 23576 6556 23616
rect 8110 23604 8116 23656
rect 8168 23644 8174 23656
rect 8404 23644 8432 23675
rect 8662 23672 8668 23724
rect 8720 23712 8726 23724
rect 8757 23715 8815 23721
rect 8757 23712 8769 23715
rect 8720 23684 8769 23712
rect 8720 23672 8726 23684
rect 8757 23681 8769 23684
rect 8803 23681 8815 23715
rect 8757 23675 8815 23681
rect 8846 23672 8852 23724
rect 8904 23672 8910 23724
rect 8941 23715 8999 23721
rect 8941 23681 8953 23715
rect 8987 23681 8999 23715
rect 8941 23675 8999 23681
rect 9125 23715 9183 23721
rect 9125 23681 9137 23715
rect 9171 23712 9183 23715
rect 9398 23712 9404 23724
rect 9171 23684 9404 23712
rect 9171 23681 9183 23684
rect 9125 23675 9183 23681
rect 8956 23644 8984 23675
rect 9398 23672 9404 23684
rect 9456 23672 9462 23724
rect 9766 23672 9772 23724
rect 9824 23712 9830 23724
rect 10502 23712 10508 23724
rect 9824 23684 10508 23712
rect 9824 23672 9830 23684
rect 10502 23672 10508 23684
rect 10560 23672 10566 23724
rect 10686 23672 10692 23724
rect 10744 23712 10750 23724
rect 10965 23715 11023 23721
rect 10965 23712 10977 23715
rect 10744 23684 10977 23712
rect 10744 23672 10750 23684
rect 10965 23681 10977 23684
rect 11011 23681 11023 23715
rect 11514 23712 11520 23724
rect 10965 23675 11023 23681
rect 11164 23684 11520 23712
rect 8168 23616 8432 23644
rect 8496 23616 8984 23644
rect 8168 23604 8174 23616
rect 8294 23576 8300 23588
rect 5920 23548 6500 23576
rect 6528 23548 8300 23576
rect 4617 23539 4675 23545
rect 6196 23520 6224 23548
rect 5626 23468 5632 23520
rect 5684 23468 5690 23520
rect 6178 23468 6184 23520
rect 6236 23468 6242 23520
rect 6362 23468 6368 23520
rect 6420 23468 6426 23520
rect 6472 23508 6500 23548
rect 8294 23536 8300 23548
rect 8352 23536 8358 23588
rect 8496 23508 8524 23616
rect 6472 23480 8524 23508
rect 8570 23468 8576 23520
rect 8628 23468 8634 23520
rect 8956 23508 8984 23616
rect 10853 23647 10911 23653
rect 10853 23613 10865 23647
rect 10899 23644 10911 23647
rect 11164 23644 11192 23684
rect 11514 23672 11520 23684
rect 11572 23712 11578 23724
rect 11882 23712 11888 23724
rect 11572 23684 11888 23712
rect 11572 23672 11578 23684
rect 11882 23672 11888 23684
rect 11940 23672 11946 23724
rect 13538 23672 13544 23724
rect 13596 23672 13602 23724
rect 13722 23672 13728 23724
rect 13780 23712 13786 23724
rect 14642 23712 14648 23724
rect 13780 23684 14648 23712
rect 13780 23672 13786 23684
rect 14642 23672 14648 23684
rect 14700 23712 14706 23724
rect 15013 23715 15071 23721
rect 15013 23712 15025 23715
rect 14700 23684 15025 23712
rect 14700 23672 14706 23684
rect 15013 23681 15025 23684
rect 15059 23681 15071 23715
rect 15013 23675 15071 23681
rect 15194 23672 15200 23724
rect 15252 23672 15258 23724
rect 15470 23672 15476 23724
rect 15528 23672 15534 23724
rect 15654 23672 15660 23724
rect 15712 23712 15718 23724
rect 15749 23715 15807 23721
rect 15749 23712 15761 23715
rect 15712 23684 15761 23712
rect 15712 23672 15718 23684
rect 15749 23681 15761 23684
rect 15795 23681 15807 23715
rect 15749 23675 15807 23681
rect 15933 23715 15991 23721
rect 15933 23681 15945 23715
rect 15979 23712 15991 23715
rect 16114 23712 16120 23724
rect 15979 23684 16120 23712
rect 15979 23681 15991 23684
rect 15933 23675 15991 23681
rect 16114 23672 16120 23684
rect 16172 23672 16178 23724
rect 10899 23616 11192 23644
rect 11241 23647 11299 23653
rect 10899 23613 10911 23616
rect 10853 23607 10911 23613
rect 11241 23613 11253 23647
rect 11287 23644 11299 23647
rect 11330 23644 11336 23656
rect 11287 23616 11336 23644
rect 11287 23613 11299 23616
rect 11241 23607 11299 23613
rect 11330 23604 11336 23616
rect 11388 23644 11394 23656
rect 11698 23644 11704 23656
rect 11388 23616 11704 23644
rect 11388 23604 11394 23616
rect 11698 23604 11704 23616
rect 11756 23604 11762 23656
rect 12161 23647 12219 23653
rect 12161 23613 12173 23647
rect 12207 23613 12219 23647
rect 12161 23607 12219 23613
rect 10686 23536 10692 23588
rect 10744 23536 10750 23588
rect 11146 23508 11152 23520
rect 8956 23480 11152 23508
rect 11146 23468 11152 23480
rect 11204 23468 11210 23520
rect 11238 23468 11244 23520
rect 11296 23508 11302 23520
rect 12176 23508 12204 23607
rect 12434 23604 12440 23656
rect 12492 23604 12498 23656
rect 13906 23604 13912 23656
rect 13964 23644 13970 23656
rect 14553 23647 14611 23653
rect 14553 23644 14565 23647
rect 13964 23616 14565 23644
rect 13964 23604 13970 23616
rect 14553 23613 14565 23616
rect 14599 23613 14611 23647
rect 16684 23644 16712 23752
rect 18046 23740 18052 23752
rect 18104 23740 18110 23792
rect 18966 23780 18972 23792
rect 18800 23752 18972 23780
rect 16758 23672 16764 23724
rect 16816 23712 16822 23724
rect 17313 23715 17371 23721
rect 17313 23712 17325 23715
rect 16816 23684 17325 23712
rect 16816 23672 16822 23684
rect 17313 23681 17325 23684
rect 17359 23712 17371 23715
rect 17954 23712 17960 23724
rect 17359 23684 17960 23712
rect 17359 23681 17371 23684
rect 17313 23675 17371 23681
rect 17954 23672 17960 23684
rect 18012 23672 18018 23724
rect 18800 23721 18828 23752
rect 18966 23740 18972 23752
rect 19024 23740 19030 23792
rect 19352 23789 19380 23820
rect 19886 23808 19892 23820
rect 19944 23808 19950 23860
rect 20073 23851 20131 23857
rect 20073 23817 20085 23851
rect 20119 23848 20131 23851
rect 20119 23820 20392 23848
rect 20119 23817 20131 23820
rect 20073 23811 20131 23817
rect 20364 23792 20392 23820
rect 20438 23808 20444 23860
rect 20496 23808 20502 23860
rect 23750 23808 23756 23860
rect 23808 23808 23814 23860
rect 23860 23820 27200 23848
rect 19337 23783 19395 23789
rect 19337 23749 19349 23783
rect 19383 23749 19395 23783
rect 19337 23743 19395 23749
rect 19444 23752 20300 23780
rect 18141 23715 18199 23721
rect 18141 23681 18153 23715
rect 18187 23712 18199 23715
rect 18785 23715 18843 23721
rect 18187 23684 18736 23712
rect 18187 23681 18199 23684
rect 18141 23675 18199 23681
rect 14553 23607 14611 23613
rect 15304 23616 16712 23644
rect 13538 23536 13544 23588
rect 13596 23576 13602 23588
rect 15304 23576 15332 23616
rect 17034 23604 17040 23656
rect 17092 23604 17098 23656
rect 17402 23604 17408 23656
rect 17460 23644 17466 23656
rect 17589 23647 17647 23653
rect 17589 23644 17601 23647
rect 17460 23616 17601 23644
rect 17460 23604 17466 23616
rect 17589 23613 17601 23616
rect 17635 23613 17647 23647
rect 17589 23607 17647 23613
rect 18046 23604 18052 23656
rect 18104 23644 18110 23656
rect 18325 23647 18383 23653
rect 18325 23644 18337 23647
rect 18104 23616 18337 23644
rect 18104 23604 18110 23616
rect 18325 23613 18337 23616
rect 18371 23644 18383 23647
rect 18414 23644 18420 23656
rect 18371 23616 18420 23644
rect 18371 23613 18383 23616
rect 18325 23607 18383 23613
rect 18414 23604 18420 23616
rect 18472 23604 18478 23656
rect 18708 23644 18736 23684
rect 18785 23681 18797 23715
rect 18831 23681 18843 23715
rect 19444 23712 19472 23752
rect 18785 23675 18843 23681
rect 19076 23684 19472 23712
rect 19076 23656 19104 23684
rect 19518 23672 19524 23724
rect 19576 23672 19582 23724
rect 19886 23672 19892 23724
rect 19944 23672 19950 23724
rect 20165 23715 20223 23721
rect 20165 23681 20177 23715
rect 20211 23681 20223 23715
rect 20272 23712 20300 23752
rect 20346 23740 20352 23792
rect 20404 23740 20410 23792
rect 20622 23789 20628 23792
rect 20609 23783 20628 23789
rect 20609 23749 20621 23783
rect 20609 23743 20628 23749
rect 20622 23740 20628 23743
rect 20680 23740 20686 23792
rect 20809 23783 20867 23789
rect 20809 23749 20821 23783
rect 20855 23780 20867 23783
rect 21266 23780 21272 23792
rect 20855 23752 21272 23780
rect 20855 23749 20867 23752
rect 20809 23743 20867 23749
rect 20824 23712 20852 23743
rect 21266 23740 21272 23752
rect 21324 23740 21330 23792
rect 23201 23783 23259 23789
rect 23201 23749 23213 23783
rect 23247 23749 23259 23783
rect 23201 23746 23259 23749
rect 23124 23743 23259 23746
rect 23293 23783 23351 23789
rect 23293 23749 23305 23783
rect 23339 23780 23351 23783
rect 23339 23752 23520 23780
rect 23339 23749 23351 23752
rect 23293 23743 23351 23749
rect 23124 23724 23244 23743
rect 20272 23684 20852 23712
rect 20165 23675 20223 23681
rect 18969 23647 19027 23653
rect 18969 23644 18981 23647
rect 18708 23616 18981 23644
rect 18969 23613 18981 23616
rect 19015 23613 19027 23647
rect 18969 23607 19027 23613
rect 13596 23548 15332 23576
rect 15381 23579 15439 23585
rect 13596 23536 13602 23548
rect 15381 23545 15393 23579
rect 15427 23576 15439 23579
rect 16574 23576 16580 23588
rect 15427 23548 16580 23576
rect 15427 23545 15439 23548
rect 15381 23539 15439 23545
rect 16574 23536 16580 23548
rect 16632 23536 16638 23588
rect 11296 23480 12204 23508
rect 11296 23468 11302 23480
rect 13906 23468 13912 23520
rect 13964 23468 13970 23520
rect 13998 23468 14004 23520
rect 14056 23468 14062 23520
rect 15470 23468 15476 23520
rect 15528 23508 15534 23520
rect 15565 23511 15623 23517
rect 15565 23508 15577 23511
rect 15528 23480 15577 23508
rect 15528 23468 15534 23480
rect 15565 23477 15577 23480
rect 15611 23477 15623 23511
rect 15565 23471 15623 23477
rect 15930 23468 15936 23520
rect 15988 23468 15994 23520
rect 18984 23508 19012 23607
rect 19058 23604 19064 23656
rect 19116 23604 19122 23656
rect 19150 23604 19156 23656
rect 19208 23644 19214 23656
rect 19334 23644 19340 23656
rect 19208 23616 19340 23644
rect 19208 23604 19214 23616
rect 19334 23604 19340 23616
rect 19392 23604 19398 23656
rect 20180 23644 20208 23675
rect 22554 23672 22560 23724
rect 22612 23672 22618 23724
rect 22738 23672 22744 23724
rect 22796 23672 22802 23724
rect 22925 23715 22983 23721
rect 22925 23681 22937 23715
rect 22971 23712 22983 23715
rect 23017 23715 23075 23721
rect 23017 23712 23029 23715
rect 22971 23684 23029 23712
rect 22971 23681 22983 23684
rect 22925 23675 22983 23681
rect 23017 23681 23029 23684
rect 23063 23681 23075 23715
rect 23017 23675 23075 23681
rect 23106 23672 23112 23724
rect 23164 23718 23244 23724
rect 23164 23672 23170 23718
rect 23385 23715 23443 23721
rect 23385 23681 23397 23715
rect 23431 23681 23443 23715
rect 23492 23712 23520 23752
rect 23750 23712 23756 23724
rect 23492 23684 23756 23712
rect 23385 23675 23443 23681
rect 20806 23644 20812 23656
rect 20180 23616 20812 23644
rect 20806 23604 20812 23616
rect 20864 23604 20870 23656
rect 22094 23536 22100 23588
rect 22152 23576 22158 23588
rect 23400 23576 23428 23675
rect 23750 23672 23756 23684
rect 23808 23712 23814 23724
rect 23860 23712 23888 23820
rect 25590 23740 25596 23792
rect 25648 23780 25654 23792
rect 26418 23780 26424 23792
rect 25648 23752 26424 23780
rect 25648 23740 25654 23752
rect 26418 23740 26424 23752
rect 26476 23740 26482 23792
rect 27172 23789 27200 23820
rect 27706 23808 27712 23860
rect 27764 23848 27770 23860
rect 27893 23851 27951 23857
rect 27893 23848 27905 23851
rect 27764 23820 27905 23848
rect 27764 23808 27770 23820
rect 27893 23817 27905 23820
rect 27939 23817 27951 23851
rect 28718 23848 28724 23860
rect 27893 23811 27951 23817
rect 28460 23820 28724 23848
rect 27157 23783 27215 23789
rect 27157 23749 27169 23783
rect 27203 23749 27215 23783
rect 27157 23743 27215 23749
rect 27246 23740 27252 23792
rect 27304 23780 27310 23792
rect 28460 23780 28488 23820
rect 28718 23808 28724 23820
rect 28776 23808 28782 23860
rect 28994 23808 29000 23860
rect 29052 23848 29058 23860
rect 29089 23851 29147 23857
rect 29089 23848 29101 23851
rect 29052 23820 29101 23848
rect 29052 23808 29058 23820
rect 29089 23817 29101 23820
rect 29135 23817 29147 23851
rect 29089 23811 29147 23817
rect 31110 23808 31116 23860
rect 31168 23808 31174 23860
rect 33502 23808 33508 23860
rect 33560 23808 33566 23860
rect 33594 23808 33600 23860
rect 33652 23848 33658 23860
rect 34514 23848 34520 23860
rect 33652 23820 34520 23848
rect 33652 23808 33658 23820
rect 27304 23752 28488 23780
rect 27304 23740 27310 23752
rect 23808 23684 23888 23712
rect 23937 23715 23995 23721
rect 23808 23672 23814 23684
rect 23937 23681 23949 23715
rect 23983 23712 23995 23715
rect 24026 23712 24032 23724
rect 23983 23684 24032 23712
rect 23983 23681 23995 23684
rect 23937 23675 23995 23681
rect 24026 23672 24032 23684
rect 24084 23672 24090 23724
rect 26973 23715 27031 23721
rect 26973 23681 26985 23715
rect 27019 23681 27031 23715
rect 26973 23675 27031 23681
rect 23474 23604 23480 23656
rect 23532 23644 23538 23656
rect 24121 23647 24179 23653
rect 24121 23644 24133 23647
rect 23532 23616 24133 23644
rect 23532 23604 23538 23616
rect 24121 23613 24133 23616
rect 24167 23613 24179 23647
rect 24121 23607 24179 23613
rect 24210 23604 24216 23656
rect 24268 23644 24274 23656
rect 26694 23644 26700 23656
rect 24268 23616 26700 23644
rect 24268 23604 24274 23616
rect 26694 23604 26700 23616
rect 26752 23644 26758 23656
rect 26988 23644 27016 23675
rect 27982 23672 27988 23724
rect 28040 23712 28046 23724
rect 28077 23715 28135 23721
rect 28077 23712 28089 23715
rect 28040 23684 28089 23712
rect 28040 23672 28046 23684
rect 28077 23681 28089 23684
rect 28123 23681 28135 23715
rect 28077 23675 28135 23681
rect 28242 23715 28300 23721
rect 28242 23681 28254 23715
rect 28288 23681 28300 23715
rect 28242 23675 28300 23681
rect 28257 23644 28285 23675
rect 28350 23672 28356 23724
rect 28408 23672 28414 23724
rect 28460 23721 28488 23752
rect 28828 23752 29040 23780
rect 28828 23746 28856 23752
rect 28736 23724 28856 23746
rect 28445 23715 28503 23721
rect 28445 23681 28457 23715
rect 28491 23681 28503 23715
rect 28445 23675 28503 23681
rect 28534 23672 28540 23724
rect 28592 23672 28598 23724
rect 28718 23672 28724 23724
rect 28776 23721 28856 23724
rect 28776 23718 28871 23721
rect 28776 23672 28782 23718
rect 28813 23715 28871 23718
rect 28813 23681 28825 23715
rect 28859 23681 28871 23715
rect 28813 23675 28871 23681
rect 28902 23672 28908 23724
rect 28960 23672 28966 23724
rect 29012 23712 29040 23752
rect 29178 23740 29184 23792
rect 29236 23780 29242 23792
rect 29638 23780 29644 23792
rect 29236 23752 29644 23780
rect 29236 23740 29242 23752
rect 29638 23740 29644 23752
rect 29696 23740 29702 23792
rect 34026 23780 34054 23820
rect 34514 23808 34520 23820
rect 34572 23808 34578 23860
rect 34609 23851 34667 23857
rect 34609 23817 34621 23851
rect 34655 23848 34667 23851
rect 38838 23848 38844 23860
rect 34655 23820 34744 23848
rect 34655 23817 34667 23820
rect 34609 23811 34667 23817
rect 34716 23789 34744 23820
rect 37660 23820 38844 23848
rect 34701 23783 34759 23789
rect 33980 23752 34054 23780
rect 34164 23752 34652 23780
rect 30374 23712 30380 23724
rect 29012 23684 30380 23712
rect 30374 23672 30380 23684
rect 30432 23672 30438 23724
rect 30926 23672 30932 23724
rect 30984 23712 30990 23724
rect 31021 23715 31079 23721
rect 31021 23712 31033 23715
rect 30984 23684 31033 23712
rect 30984 23672 30990 23684
rect 31021 23681 31033 23684
rect 31067 23681 31079 23715
rect 31021 23675 31079 23681
rect 31205 23715 31263 23721
rect 31205 23681 31217 23715
rect 31251 23681 31263 23715
rect 31205 23675 31263 23681
rect 26752 23616 28285 23644
rect 28552 23644 28580 23672
rect 29181 23647 29239 23653
rect 29181 23644 29193 23647
rect 28552 23616 29193 23644
rect 26752 23604 26758 23616
rect 29181 23613 29193 23616
rect 29227 23613 29239 23647
rect 31220 23644 31248 23675
rect 31478 23672 31484 23724
rect 31536 23672 31542 23724
rect 32950 23672 32956 23724
rect 33008 23712 33014 23724
rect 33045 23715 33103 23721
rect 33045 23712 33057 23715
rect 33008 23684 33057 23712
rect 33008 23672 33014 23684
rect 33045 23681 33057 23684
rect 33091 23681 33103 23715
rect 33045 23675 33103 23681
rect 33134 23672 33140 23724
rect 33192 23712 33198 23724
rect 33980 23721 34008 23752
rect 34164 23721 34192 23752
rect 33321 23715 33379 23721
rect 33321 23712 33333 23715
rect 33192 23684 33333 23712
rect 33192 23672 33198 23684
rect 33321 23681 33333 23684
rect 33367 23681 33379 23715
rect 33321 23675 33379 23681
rect 33965 23715 34023 23721
rect 33965 23681 33977 23715
rect 34011 23681 34023 23715
rect 33965 23675 34023 23681
rect 34113 23715 34192 23721
rect 34113 23681 34125 23715
rect 34159 23684 34192 23715
rect 34241 23715 34299 23721
rect 34159 23681 34171 23684
rect 34113 23675 34171 23681
rect 34241 23681 34253 23715
rect 34287 23681 34299 23715
rect 34241 23675 34299 23681
rect 31496 23644 31524 23672
rect 32306 23644 32312 23656
rect 31220 23616 32312 23644
rect 29181 23607 29239 23613
rect 32306 23604 32312 23616
rect 32364 23604 32370 23656
rect 33229 23647 33287 23653
rect 33229 23613 33241 23647
rect 33275 23644 33287 23647
rect 33686 23644 33692 23656
rect 33275 23616 33692 23644
rect 33275 23613 33287 23616
rect 33229 23607 33287 23613
rect 33686 23604 33692 23616
rect 33744 23604 33750 23656
rect 34256 23644 34284 23675
rect 34330 23672 34336 23724
rect 34388 23672 34394 23724
rect 34430 23715 34488 23721
rect 34430 23681 34442 23715
rect 34476 23681 34488 23715
rect 34624 23712 34652 23752
rect 34701 23749 34713 23783
rect 34747 23749 34759 23783
rect 36354 23780 36360 23792
rect 34701 23743 34759 23749
rect 34808 23752 36360 23780
rect 34808 23712 34836 23752
rect 36354 23740 36360 23752
rect 36412 23740 36418 23792
rect 34624 23684 34836 23712
rect 34430 23675 34488 23681
rect 34164 23616 34284 23644
rect 34164 23588 34192 23616
rect 23569 23579 23627 23585
rect 22152 23548 23520 23576
rect 22152 23536 22158 23548
rect 19334 23508 19340 23520
rect 18984 23480 19340 23508
rect 19334 23468 19340 23480
rect 19392 23468 19398 23520
rect 19889 23511 19947 23517
rect 19889 23477 19901 23511
rect 19935 23508 19947 23511
rect 20070 23508 20076 23520
rect 19935 23480 20076 23508
rect 19935 23477 19947 23480
rect 19889 23471 19947 23477
rect 20070 23468 20076 23480
rect 20128 23468 20134 23520
rect 20625 23511 20683 23517
rect 20625 23477 20637 23511
rect 20671 23508 20683 23511
rect 21266 23508 21272 23520
rect 20671 23480 21272 23508
rect 20671 23477 20683 23480
rect 20625 23471 20683 23477
rect 21266 23468 21272 23480
rect 21324 23468 21330 23520
rect 23492 23508 23520 23548
rect 23569 23545 23581 23579
rect 23615 23576 23627 23579
rect 23842 23576 23848 23588
rect 23615 23548 23848 23576
rect 23615 23545 23627 23548
rect 23569 23539 23627 23545
rect 23842 23536 23848 23548
rect 23900 23536 23906 23588
rect 27341 23579 27399 23585
rect 27341 23545 27353 23579
rect 27387 23576 27399 23579
rect 28166 23576 28172 23588
rect 27387 23548 28172 23576
rect 27387 23545 27399 23548
rect 27341 23539 27399 23545
rect 28166 23536 28172 23548
rect 28224 23576 28230 23588
rect 28902 23576 28908 23588
rect 28224 23548 28908 23576
rect 28224 23536 28230 23548
rect 28902 23536 28908 23548
rect 28960 23536 28966 23588
rect 29270 23536 29276 23588
rect 29328 23536 29334 23588
rect 31018 23536 31024 23588
rect 31076 23576 31082 23588
rect 31478 23576 31484 23588
rect 31076 23548 31484 23576
rect 31076 23536 31082 23548
rect 31478 23536 31484 23548
rect 31536 23536 31542 23588
rect 34146 23536 34152 23588
rect 34204 23536 34210 23588
rect 34445 23576 34473 23675
rect 34882 23672 34888 23724
rect 34940 23672 34946 23724
rect 36541 23715 36599 23721
rect 36541 23681 36553 23715
rect 36587 23712 36599 23715
rect 37550 23712 37556 23724
rect 36587 23684 37556 23712
rect 36587 23681 36599 23684
rect 36541 23675 36599 23681
rect 37550 23672 37556 23684
rect 37608 23672 37614 23724
rect 34790 23604 34796 23656
rect 34848 23644 34854 23656
rect 36725 23647 36783 23653
rect 36725 23644 36737 23647
rect 34848 23616 36737 23644
rect 34848 23604 34854 23616
rect 36725 23613 36737 23616
rect 36771 23644 36783 23647
rect 37660 23644 37688 23820
rect 38838 23808 38844 23820
rect 38896 23808 38902 23860
rect 38378 23740 38384 23792
rect 38436 23780 38442 23792
rect 38473 23783 38531 23789
rect 38473 23780 38485 23783
rect 38436 23752 38485 23780
rect 38436 23740 38442 23752
rect 38473 23749 38485 23752
rect 38519 23749 38531 23783
rect 38473 23743 38531 23749
rect 39574 23672 39580 23724
rect 39632 23672 39638 23724
rect 36771 23616 37688 23644
rect 36771 23613 36783 23616
rect 36725 23607 36783 23613
rect 38194 23604 38200 23656
rect 38252 23604 38258 23656
rect 39114 23604 39120 23656
rect 39172 23644 39178 23656
rect 39482 23644 39488 23656
rect 39172 23616 39488 23644
rect 39172 23604 39178 23616
rect 39482 23604 39488 23616
rect 39540 23644 39546 23656
rect 40221 23647 40279 23653
rect 40221 23644 40233 23647
rect 39540 23616 40233 23644
rect 39540 23604 39546 23616
rect 40221 23613 40233 23616
rect 40267 23613 40279 23647
rect 40221 23607 40279 23613
rect 34445 23548 34836 23576
rect 34808 23520 34836 23548
rect 28629 23511 28687 23517
rect 28629 23508 28641 23511
rect 23492 23480 28641 23508
rect 28629 23477 28641 23480
rect 28675 23508 28687 23511
rect 28810 23508 28816 23520
rect 28675 23480 28816 23508
rect 28675 23477 28687 23480
rect 28629 23471 28687 23477
rect 28810 23468 28816 23480
rect 28868 23468 28874 23520
rect 31570 23468 31576 23520
rect 31628 23508 31634 23520
rect 32306 23508 32312 23520
rect 31628 23480 32312 23508
rect 31628 23468 31634 23480
rect 32306 23468 32312 23480
rect 32364 23468 32370 23520
rect 33042 23468 33048 23520
rect 33100 23468 33106 23520
rect 34790 23468 34796 23520
rect 34848 23468 34854 23520
rect 35069 23511 35127 23517
rect 35069 23477 35081 23511
rect 35115 23508 35127 23511
rect 37918 23508 37924 23520
rect 35115 23480 37924 23508
rect 35115 23477 35127 23480
rect 35069 23471 35127 23477
rect 37918 23468 37924 23480
rect 37976 23468 37982 23520
rect 1104 23418 40572 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 40572 23418
rect 1104 23344 40572 23366
rect 4433 23307 4491 23313
rect 4433 23273 4445 23307
rect 4479 23304 4491 23307
rect 4706 23304 4712 23316
rect 4479 23276 4712 23304
rect 4479 23273 4491 23276
rect 4433 23267 4491 23273
rect 4706 23264 4712 23276
rect 4764 23264 4770 23316
rect 9033 23307 9091 23313
rect 9033 23273 9045 23307
rect 9079 23304 9091 23307
rect 9214 23304 9220 23316
rect 9079 23276 9220 23304
rect 9079 23273 9091 23276
rect 9033 23267 9091 23273
rect 9214 23264 9220 23276
rect 9272 23264 9278 23316
rect 9490 23264 9496 23316
rect 9548 23304 9554 23316
rect 9861 23307 9919 23313
rect 9861 23304 9873 23307
rect 9548 23276 9873 23304
rect 9548 23264 9554 23276
rect 9861 23273 9873 23276
rect 9907 23273 9919 23307
rect 9861 23267 9919 23273
rect 10318 23264 10324 23316
rect 10376 23264 10382 23316
rect 11514 23264 11520 23316
rect 11572 23304 11578 23316
rect 11572 23276 12112 23304
rect 11572 23264 11578 23276
rect 5261 23239 5319 23245
rect 5261 23205 5273 23239
rect 5307 23236 5319 23239
rect 5537 23239 5595 23245
rect 5537 23236 5549 23239
rect 5307 23208 5549 23236
rect 5307 23205 5319 23208
rect 5261 23199 5319 23205
rect 5537 23205 5549 23208
rect 5583 23205 5595 23239
rect 5537 23199 5595 23205
rect 5626 23196 5632 23248
rect 5684 23196 5690 23248
rect 5905 23239 5963 23245
rect 5905 23205 5917 23239
rect 5951 23236 5963 23239
rect 5951 23208 8340 23236
rect 5951 23205 5963 23208
rect 5905 23199 5963 23205
rect 3234 23128 3240 23180
rect 3292 23168 3298 23180
rect 3605 23171 3663 23177
rect 3605 23168 3617 23171
rect 3292 23140 3617 23168
rect 3292 23128 3298 23140
rect 3605 23137 3617 23140
rect 3651 23168 3663 23171
rect 6270 23168 6276 23180
rect 3651 23140 5028 23168
rect 3651 23137 3663 23140
rect 3605 23131 3663 23137
rect 2409 23103 2467 23109
rect 2409 23069 2421 23103
rect 2455 23100 2467 23103
rect 2866 23100 2872 23112
rect 2455 23072 2872 23100
rect 2455 23069 2467 23072
rect 2409 23063 2467 23069
rect 2866 23060 2872 23072
rect 2924 23060 2930 23112
rect 3970 23060 3976 23112
rect 4028 23100 4034 23112
rect 5000 23109 5028 23140
rect 5368 23140 6276 23168
rect 4709 23103 4767 23109
rect 4709 23100 4721 23103
rect 4028 23072 4721 23100
rect 4028 23060 4034 23072
rect 4709 23069 4721 23072
rect 4755 23069 4767 23103
rect 4709 23063 4767 23069
rect 4985 23103 5043 23109
rect 4985 23069 4997 23103
rect 5031 23069 5043 23103
rect 4985 23063 5043 23069
rect 5077 23103 5135 23109
rect 5077 23069 5089 23103
rect 5123 23100 5135 23103
rect 5258 23100 5264 23112
rect 5123 23072 5264 23100
rect 5123 23069 5135 23072
rect 5077 23063 5135 23069
rect 5258 23060 5264 23072
rect 5316 23060 5322 23112
rect 4525 23035 4583 23041
rect 4525 23001 4537 23035
rect 4571 23001 4583 23035
rect 4525 22995 4583 23001
rect 4893 23035 4951 23041
rect 4893 23001 4905 23035
rect 4939 23032 4951 23035
rect 5368 23032 5396 23140
rect 6270 23128 6276 23140
rect 6328 23128 6334 23180
rect 8312 23168 8340 23208
rect 8386 23196 8392 23248
rect 8444 23236 8450 23248
rect 8938 23236 8944 23248
rect 8444 23208 8944 23236
rect 8444 23196 8450 23208
rect 8938 23196 8944 23208
rect 8996 23236 9002 23248
rect 11974 23236 11980 23248
rect 8996 23208 11980 23236
rect 8996 23196 9002 23208
rect 11974 23196 11980 23208
rect 12032 23196 12038 23248
rect 12084 23236 12112 23276
rect 12158 23264 12164 23316
rect 12216 23264 12222 23316
rect 12434 23264 12440 23316
rect 12492 23304 12498 23316
rect 12621 23307 12679 23313
rect 12621 23304 12633 23307
rect 12492 23276 12633 23304
rect 12492 23264 12498 23276
rect 12621 23273 12633 23276
rect 12667 23273 12679 23307
rect 12621 23267 12679 23273
rect 16574 23264 16580 23316
rect 16632 23264 16638 23316
rect 16666 23264 16672 23316
rect 16724 23304 16730 23316
rect 16761 23307 16819 23313
rect 16761 23304 16773 23307
rect 16724 23276 16773 23304
rect 16724 23264 16730 23276
rect 16761 23273 16773 23276
rect 16807 23273 16819 23307
rect 16761 23267 16819 23273
rect 18046 23264 18052 23316
rect 18104 23264 18110 23316
rect 18141 23307 18199 23313
rect 18141 23273 18153 23307
rect 18187 23304 18199 23307
rect 18690 23304 18696 23316
rect 18187 23276 18696 23304
rect 18187 23273 18199 23276
rect 18141 23267 18199 23273
rect 18690 23264 18696 23276
rect 18748 23264 18754 23316
rect 19518 23264 19524 23316
rect 19576 23304 19582 23316
rect 23290 23304 23296 23316
rect 19576 23276 23296 23304
rect 19576 23264 19582 23276
rect 23290 23264 23296 23276
rect 23348 23264 23354 23316
rect 24486 23264 24492 23316
rect 24544 23304 24550 23316
rect 29089 23307 29147 23313
rect 29089 23304 29101 23307
rect 24544 23276 29101 23304
rect 24544 23264 24550 23276
rect 29089 23273 29101 23276
rect 29135 23304 29147 23307
rect 29270 23304 29276 23316
rect 29135 23276 29276 23304
rect 29135 23273 29147 23276
rect 29089 23267 29147 23273
rect 29270 23264 29276 23276
rect 29328 23264 29334 23316
rect 34146 23264 34152 23316
rect 34204 23304 34210 23316
rect 37274 23304 37280 23316
rect 34204 23276 37280 23304
rect 34204 23264 34210 23276
rect 37274 23264 37280 23276
rect 37332 23264 37338 23316
rect 38289 23307 38347 23313
rect 38289 23273 38301 23307
rect 38335 23304 38347 23307
rect 38378 23304 38384 23316
rect 38335 23276 38384 23304
rect 38335 23273 38347 23276
rect 38289 23267 38347 23273
rect 38378 23264 38384 23276
rect 38436 23264 38442 23316
rect 38657 23307 38715 23313
rect 38657 23273 38669 23307
rect 38703 23273 38715 23307
rect 38657 23267 38715 23273
rect 39485 23307 39543 23313
rect 39485 23273 39497 23307
rect 39531 23304 39543 23307
rect 39574 23304 39580 23316
rect 39531 23276 39580 23304
rect 39531 23273 39543 23276
rect 39485 23267 39543 23273
rect 12084 23208 12204 23236
rect 9766 23168 9772 23180
rect 8312 23140 9772 23168
rect 9766 23128 9772 23140
rect 9824 23128 9830 23180
rect 10229 23171 10287 23177
rect 10229 23137 10241 23171
rect 10275 23168 10287 23171
rect 10870 23168 10876 23180
rect 10275 23140 10876 23168
rect 10275 23137 10287 23140
rect 10229 23131 10287 23137
rect 10870 23128 10876 23140
rect 10928 23168 10934 23180
rect 11514 23168 11520 23180
rect 10928 23140 11520 23168
rect 10928 23128 10934 23140
rect 11514 23128 11520 23140
rect 11572 23128 11578 23180
rect 11609 23171 11667 23177
rect 11609 23137 11621 23171
rect 11655 23168 11667 23171
rect 12066 23168 12072 23180
rect 11655 23140 12072 23168
rect 11655 23137 11667 23140
rect 11609 23131 11667 23137
rect 12066 23128 12072 23140
rect 12124 23128 12130 23180
rect 5445 23103 5503 23109
rect 5445 23069 5457 23103
rect 5491 23100 5503 23103
rect 5721 23103 5779 23109
rect 5491 23072 5672 23100
rect 5491 23069 5503 23072
rect 5445 23063 5503 23069
rect 5644 23044 5672 23072
rect 5721 23069 5733 23103
rect 5767 23069 5779 23103
rect 5721 23063 5779 23069
rect 4939 23004 5396 23032
rect 4939 23001 4951 23004
rect 4893 22995 4951 23001
rect 2590 22924 2596 22976
rect 2648 22964 2654 22976
rect 2961 22967 3019 22973
rect 2961 22964 2973 22967
rect 2648 22936 2973 22964
rect 2648 22924 2654 22936
rect 2961 22933 2973 22936
rect 3007 22933 3019 22967
rect 4540 22964 4568 22995
rect 5626 22992 5632 23044
rect 5684 22992 5690 23044
rect 5736 23032 5764 23063
rect 6086 23060 6092 23112
rect 6144 23060 6150 23112
rect 6362 23060 6368 23112
rect 6420 23060 6426 23112
rect 6730 23060 6736 23112
rect 6788 23060 6794 23112
rect 7469 23103 7527 23109
rect 7469 23069 7481 23103
rect 7515 23100 7527 23103
rect 7834 23100 7840 23112
rect 7515 23072 7840 23100
rect 7515 23069 7527 23072
rect 7469 23063 7527 23069
rect 7834 23060 7840 23072
rect 7892 23060 7898 23112
rect 8938 23060 8944 23112
rect 8996 23060 9002 23112
rect 9125 23103 9183 23109
rect 9125 23069 9137 23103
rect 9171 23100 9183 23103
rect 9171 23072 10456 23100
rect 9171 23069 9183 23072
rect 9125 23063 9183 23069
rect 10428 23044 10456 23072
rect 10502 23060 10508 23112
rect 10560 23060 10566 23112
rect 10597 23103 10655 23109
rect 10597 23069 10609 23103
rect 10643 23069 10655 23103
rect 10597 23063 10655 23069
rect 11146 23103 11204 23109
rect 11146 23069 11158 23103
rect 11192 23100 11204 23103
rect 11330 23100 11336 23112
rect 11192 23072 11336 23100
rect 11192 23069 11204 23072
rect 11146 23063 11204 23069
rect 6270 23032 6276 23044
rect 5736 23004 6276 23032
rect 6270 22992 6276 23004
rect 6328 22992 6334 23044
rect 7193 23035 7251 23041
rect 7193 23001 7205 23035
rect 7239 23032 7251 23035
rect 7239 23004 9674 23032
rect 7239 23001 7251 23004
rect 7193 22995 7251 23001
rect 7742 22964 7748 22976
rect 4540 22936 7748 22964
rect 2961 22927 3019 22933
rect 7742 22924 7748 22936
rect 7800 22964 7806 22976
rect 9490 22964 9496 22976
rect 7800 22936 9496 22964
rect 7800 22924 7806 22936
rect 9490 22924 9496 22936
rect 9548 22924 9554 22976
rect 9646 22964 9674 23004
rect 9766 22992 9772 23044
rect 9824 22992 9830 23044
rect 10410 22992 10416 23044
rect 10468 22992 10474 23044
rect 9950 22964 9956 22976
rect 9646 22936 9956 22964
rect 9950 22924 9956 22936
rect 10008 22964 10014 22976
rect 10612 22964 10640 23063
rect 11330 23060 11336 23072
rect 11388 23060 11394 23112
rect 11885 23103 11943 23109
rect 11885 23100 11897 23103
rect 11808 23072 11897 23100
rect 11698 22992 11704 23044
rect 11756 22992 11762 23044
rect 10008 22936 10640 22964
rect 10008 22924 10014 22936
rect 10686 22924 10692 22976
rect 10744 22964 10750 22976
rect 10781 22967 10839 22973
rect 10781 22964 10793 22967
rect 10744 22936 10793 22964
rect 10744 22924 10750 22936
rect 10781 22933 10793 22936
rect 10827 22933 10839 22967
rect 10781 22927 10839 22933
rect 10962 22924 10968 22976
rect 11020 22924 11026 22976
rect 11149 22967 11207 22973
rect 11149 22933 11161 22967
rect 11195 22964 11207 22967
rect 11422 22964 11428 22976
rect 11195 22936 11428 22964
rect 11195 22933 11207 22936
rect 11149 22927 11207 22933
rect 11422 22924 11428 22936
rect 11480 22924 11486 22976
rect 11514 22924 11520 22976
rect 11572 22964 11578 22976
rect 11808 22964 11836 23072
rect 11885 23069 11897 23072
rect 11931 23069 11943 23103
rect 11885 23063 11943 23069
rect 11977 23103 12035 23109
rect 11977 23069 11989 23103
rect 12023 23069 12035 23103
rect 12176 23100 12204 23208
rect 14734 23196 14740 23248
rect 14792 23196 14798 23248
rect 19058 23236 19064 23248
rect 17972 23208 19064 23236
rect 13081 23171 13139 23177
rect 13081 23137 13093 23171
rect 13127 23168 13139 23171
rect 13170 23168 13176 23180
rect 13127 23140 13176 23168
rect 13127 23137 13139 23140
rect 13081 23131 13139 23137
rect 13170 23128 13176 23140
rect 13228 23128 13234 23180
rect 13265 23171 13323 23177
rect 13265 23137 13277 23171
rect 13311 23168 13323 23171
rect 13446 23168 13452 23180
rect 13311 23140 13452 23168
rect 13311 23137 13323 23140
rect 13265 23131 13323 23137
rect 13446 23128 13452 23140
rect 13504 23128 13510 23180
rect 17972 23177 18000 23208
rect 19058 23196 19064 23208
rect 19116 23196 19122 23248
rect 19150 23196 19156 23248
rect 19208 23236 19214 23248
rect 25866 23236 25872 23248
rect 19208 23208 25872 23236
rect 19208 23196 19214 23208
rect 25866 23196 25872 23208
rect 25924 23196 25930 23248
rect 27798 23196 27804 23248
rect 27856 23236 27862 23248
rect 28902 23236 28908 23248
rect 27856 23208 28908 23236
rect 27856 23196 27862 23208
rect 28902 23196 28908 23208
rect 28960 23196 28966 23248
rect 29288 23236 29316 23264
rect 30190 23236 30196 23248
rect 29288 23208 30196 23236
rect 30190 23196 30196 23208
rect 30248 23196 30254 23248
rect 31757 23239 31815 23245
rect 31757 23205 31769 23239
rect 31803 23236 31815 23239
rect 31803 23208 33732 23236
rect 31803 23205 31815 23208
rect 31757 23199 31815 23205
rect 17957 23171 18015 23177
rect 17957 23137 17969 23171
rect 18003 23137 18015 23171
rect 17957 23131 18015 23137
rect 18690 23128 18696 23180
rect 18748 23168 18754 23180
rect 24026 23168 24032 23180
rect 18748 23140 24032 23168
rect 18748 23128 18754 23140
rect 24026 23128 24032 23140
rect 24084 23128 24090 23180
rect 30208 23168 30236 23196
rect 33704 23180 33732 23208
rect 34514 23196 34520 23248
rect 34572 23236 34578 23248
rect 34572 23208 36216 23236
rect 34572 23196 34578 23208
rect 30469 23171 30527 23177
rect 30469 23168 30481 23171
rect 30208 23140 30481 23168
rect 30469 23137 30481 23140
rect 30515 23137 30527 23171
rect 30469 23131 30527 23137
rect 32030 23128 32036 23180
rect 32088 23168 32094 23180
rect 33042 23168 33048 23180
rect 32088 23140 33048 23168
rect 32088 23128 32094 23140
rect 33042 23128 33048 23140
rect 33100 23128 33106 23180
rect 33137 23171 33195 23177
rect 33137 23137 33149 23171
rect 33183 23168 33195 23171
rect 33226 23168 33232 23180
rect 33183 23140 33232 23168
rect 33183 23137 33195 23140
rect 33137 23131 33195 23137
rect 33226 23128 33232 23140
rect 33284 23128 33290 23180
rect 33410 23128 33416 23180
rect 33468 23168 33474 23180
rect 33505 23171 33563 23177
rect 33505 23168 33517 23171
rect 33468 23140 33517 23168
rect 33468 23128 33474 23140
rect 33505 23137 33517 23140
rect 33551 23137 33563 23171
rect 33505 23131 33563 23137
rect 33686 23128 33692 23180
rect 33744 23168 33750 23180
rect 36188 23168 36216 23208
rect 37550 23196 37556 23248
rect 37608 23236 37614 23248
rect 38470 23236 38476 23248
rect 37608 23208 38476 23236
rect 37608 23196 37614 23208
rect 38470 23196 38476 23208
rect 38528 23236 38534 23248
rect 38672 23236 38700 23267
rect 39574 23264 39580 23276
rect 39632 23264 39638 23316
rect 38528 23208 38700 23236
rect 38528 23196 38534 23208
rect 33744 23140 36124 23168
rect 36188 23140 38516 23168
rect 33744 23128 33750 23140
rect 12253 23103 12311 23109
rect 12253 23100 12265 23103
rect 12176 23072 12265 23100
rect 11977 23063 12035 23069
rect 12253 23069 12265 23072
rect 12299 23069 12311 23103
rect 12253 23063 12311 23069
rect 12989 23103 13047 23109
rect 12989 23069 13001 23103
rect 13035 23100 13047 23103
rect 13998 23100 14004 23112
rect 13035 23072 14004 23100
rect 13035 23069 13047 23072
rect 12989 23063 13047 23069
rect 11992 23032 12020 23063
rect 13998 23060 14004 23072
rect 14056 23060 14062 23112
rect 14366 23060 14372 23112
rect 14424 23100 14430 23112
rect 14461 23103 14519 23109
rect 14461 23100 14473 23103
rect 14424 23072 14473 23100
rect 14424 23060 14430 23072
rect 14461 23069 14473 23072
rect 14507 23069 14519 23103
rect 14461 23063 14519 23069
rect 16853 23103 16911 23109
rect 16853 23069 16865 23103
rect 16899 23069 16911 23103
rect 16853 23063 16911 23069
rect 12158 23032 12164 23044
rect 11992 23004 12164 23032
rect 12158 22992 12164 23004
rect 12216 22992 12222 23044
rect 13538 22992 13544 23044
rect 13596 23032 13602 23044
rect 13633 23035 13691 23041
rect 13633 23032 13645 23035
rect 13596 23004 13645 23032
rect 13596 22992 13602 23004
rect 13633 23001 13645 23004
rect 13679 23001 13691 23035
rect 13633 22995 13691 23001
rect 13814 22992 13820 23044
rect 13872 22992 13878 23044
rect 14185 23035 14243 23041
rect 14185 23001 14197 23035
rect 14231 23001 14243 23035
rect 16868 23032 16896 23063
rect 16942 23060 16948 23112
rect 17000 23100 17006 23112
rect 17129 23103 17187 23109
rect 17129 23100 17141 23103
rect 17000 23072 17141 23100
rect 17000 23060 17006 23072
rect 17129 23069 17141 23072
rect 17175 23069 17187 23103
rect 17129 23063 17187 23069
rect 18049 23103 18107 23109
rect 18049 23069 18061 23103
rect 18095 23100 18107 23103
rect 18230 23100 18236 23112
rect 18095 23072 18236 23100
rect 18095 23069 18107 23072
rect 18049 23063 18107 23069
rect 18230 23060 18236 23072
rect 18288 23060 18294 23112
rect 18325 23103 18383 23109
rect 18325 23069 18337 23103
rect 18371 23069 18383 23103
rect 18325 23063 18383 23069
rect 18340 23032 18368 23063
rect 18414 23060 18420 23112
rect 18472 23060 18478 23112
rect 18782 23060 18788 23112
rect 18840 23060 18846 23112
rect 19334 23060 19340 23112
rect 19392 23100 19398 23112
rect 19392 23072 19656 23100
rect 19392 23060 19398 23072
rect 19518 23032 19524 23044
rect 16868 23004 18000 23032
rect 18340 23004 19524 23032
rect 14185 22995 14243 23001
rect 11572 22936 11836 22964
rect 11572 22924 11578 22936
rect 13998 22924 14004 22976
rect 14056 22964 14062 22976
rect 14200 22964 14228 22995
rect 17972 22976 18000 23004
rect 19518 22992 19524 23004
rect 19576 22992 19582 23044
rect 19628 23032 19656 23072
rect 20070 23060 20076 23112
rect 20128 23100 20134 23112
rect 20898 23100 20904 23112
rect 20128 23072 20904 23100
rect 20128 23060 20134 23072
rect 20898 23060 20904 23072
rect 20956 23060 20962 23112
rect 21358 23060 21364 23112
rect 21416 23100 21422 23112
rect 22278 23100 22284 23112
rect 21416 23072 22284 23100
rect 21416 23060 21422 23072
rect 22278 23060 22284 23072
rect 22336 23060 22342 23112
rect 22465 23103 22523 23109
rect 22465 23069 22477 23103
rect 22511 23100 22523 23103
rect 22830 23100 22836 23112
rect 22511 23072 22836 23100
rect 22511 23069 22523 23072
rect 22465 23063 22523 23069
rect 22830 23060 22836 23072
rect 22888 23100 22894 23112
rect 23106 23100 23112 23112
rect 22888 23072 23112 23100
rect 22888 23060 22894 23072
rect 23106 23060 23112 23072
rect 23164 23060 23170 23112
rect 29822 23060 29828 23112
rect 29880 23100 29886 23112
rect 30101 23103 30159 23109
rect 30101 23100 30113 23103
rect 29880 23072 30113 23100
rect 29880 23060 29886 23072
rect 30101 23069 30113 23072
rect 30147 23069 30159 23103
rect 30101 23063 30159 23069
rect 30285 23103 30343 23109
rect 30285 23069 30297 23103
rect 30331 23069 30343 23103
rect 30285 23063 30343 23069
rect 21450 23032 21456 23044
rect 19628 23004 21456 23032
rect 21450 22992 21456 23004
rect 21508 22992 21514 23044
rect 29270 22992 29276 23044
rect 29328 22992 29334 23044
rect 30300 23032 30328 23063
rect 31202 23060 31208 23112
rect 31260 23060 31266 23112
rect 31294 23060 31300 23112
rect 31352 23100 31358 23112
rect 31481 23103 31539 23109
rect 31481 23100 31493 23103
rect 31352 23072 31493 23100
rect 31352 23060 31358 23072
rect 31481 23069 31493 23072
rect 31527 23069 31539 23103
rect 31481 23063 31539 23069
rect 31573 23103 31631 23109
rect 31573 23069 31585 23103
rect 31619 23100 31631 23103
rect 31754 23100 31760 23112
rect 31619 23072 31760 23100
rect 31619 23069 31631 23072
rect 31573 23063 31631 23069
rect 31754 23060 31760 23072
rect 31812 23060 31818 23112
rect 33428 23100 33456 23128
rect 33962 23100 33968 23112
rect 32728 23072 33968 23100
rect 31110 23032 31116 23044
rect 30024 23004 31116 23032
rect 14056 22936 14228 22964
rect 14056 22924 14062 22936
rect 14274 22924 14280 22976
rect 14332 22924 14338 22976
rect 17678 22924 17684 22976
rect 17736 22924 17742 22976
rect 17954 22924 17960 22976
rect 18012 22924 18018 22976
rect 18046 22924 18052 22976
rect 18104 22964 18110 22976
rect 18509 22967 18567 22973
rect 18509 22964 18521 22967
rect 18104 22936 18521 22964
rect 18104 22924 18110 22936
rect 18509 22933 18521 22936
rect 18555 22933 18567 22967
rect 18509 22927 18567 22933
rect 18690 22924 18696 22976
rect 18748 22964 18754 22976
rect 19242 22964 19248 22976
rect 18748 22936 19248 22964
rect 18748 22924 18754 22936
rect 19242 22924 19248 22936
rect 19300 22924 19306 22976
rect 19978 22924 19984 22976
rect 20036 22964 20042 22976
rect 21358 22964 21364 22976
rect 20036 22936 21364 22964
rect 20036 22924 20042 22936
rect 21358 22924 21364 22936
rect 21416 22964 21422 22976
rect 22281 22967 22339 22973
rect 22281 22964 22293 22967
rect 21416 22936 22293 22964
rect 21416 22924 21422 22936
rect 22281 22933 22293 22936
rect 22327 22933 22339 22967
rect 22281 22927 22339 22933
rect 27706 22924 27712 22976
rect 27764 22964 27770 22976
rect 28350 22964 28356 22976
rect 27764 22936 28356 22964
rect 27764 22924 27770 22936
rect 28350 22924 28356 22936
rect 28408 22964 28414 22976
rect 28905 22967 28963 22973
rect 28905 22964 28917 22967
rect 28408 22936 28917 22964
rect 28408 22924 28414 22936
rect 28905 22933 28917 22936
rect 28951 22933 28963 22967
rect 28905 22927 28963 22933
rect 29073 22967 29131 22973
rect 29073 22933 29085 22967
rect 29119 22964 29131 22967
rect 30024 22964 30052 23004
rect 31110 22992 31116 23004
rect 31168 22992 31174 23044
rect 31389 23035 31447 23041
rect 31389 23001 31401 23035
rect 31435 23032 31447 23035
rect 32728 23032 32756 23072
rect 33962 23060 33968 23072
rect 34020 23060 34026 23112
rect 36096 23109 36124 23140
rect 36081 23103 36139 23109
rect 36081 23069 36093 23103
rect 36127 23069 36139 23103
rect 36081 23063 36139 23069
rect 36174 23103 36232 23109
rect 36174 23069 36186 23103
rect 36220 23069 36232 23103
rect 36174 23063 36232 23069
rect 33226 23032 33232 23044
rect 31435 23004 32756 23032
rect 32784 23004 33232 23032
rect 31435 23001 31447 23004
rect 31389 22995 31447 23001
rect 29119 22936 30052 22964
rect 29119 22933 29131 22936
rect 29073 22927 29131 22933
rect 31662 22924 31668 22976
rect 31720 22964 31726 22976
rect 32784 22964 32812 23004
rect 33226 22992 33232 23004
rect 33284 22992 33290 23044
rect 33413 23035 33471 23041
rect 33413 23001 33425 23035
rect 33459 23032 33471 23035
rect 33502 23032 33508 23044
rect 33459 23004 33508 23032
rect 33459 23001 33471 23004
rect 33413 22995 33471 23001
rect 33502 22992 33508 23004
rect 33560 23032 33566 23044
rect 34238 23032 34244 23044
rect 33560 23004 34244 23032
rect 33560 22992 33566 23004
rect 34238 22992 34244 23004
rect 34296 23032 34302 23044
rect 35986 23032 35992 23044
rect 34296 23004 35992 23032
rect 34296 22992 34302 23004
rect 35986 22992 35992 23004
rect 36044 22992 36050 23044
rect 31720 22936 32812 22964
rect 31720 22924 31726 22936
rect 32858 22924 32864 22976
rect 32916 22924 32922 22976
rect 33321 22967 33379 22973
rect 33321 22933 33333 22967
rect 33367 22964 33379 22967
rect 33686 22964 33692 22976
rect 33367 22936 33692 22964
rect 33367 22933 33379 22936
rect 33321 22927 33379 22933
rect 33686 22924 33692 22936
rect 33744 22964 33750 22976
rect 35894 22964 35900 22976
rect 33744 22936 35900 22964
rect 33744 22924 33750 22936
rect 35894 22924 35900 22936
rect 35952 22964 35958 22976
rect 36188 22964 36216 23063
rect 36446 23060 36452 23112
rect 36504 23060 36510 23112
rect 36538 23060 36544 23112
rect 36596 23109 36602 23112
rect 38488 23109 38516 23140
rect 39298 23128 39304 23180
rect 39356 23168 39362 23180
rect 39482 23168 39488 23180
rect 39356 23140 39488 23168
rect 39356 23128 39362 23140
rect 39482 23128 39488 23140
rect 39540 23128 39546 23180
rect 36596 23100 36604 23109
rect 38473 23103 38531 23109
rect 36596 23072 36641 23100
rect 36596 23063 36604 23072
rect 38473 23069 38485 23103
rect 38519 23069 38531 23103
rect 38473 23063 38531 23069
rect 36596 23060 36602 23063
rect 38562 23060 38568 23112
rect 38620 23060 38626 23112
rect 39577 23103 39635 23109
rect 39577 23069 39589 23103
rect 39623 23100 39635 23103
rect 39758 23100 39764 23112
rect 39623 23072 39764 23100
rect 39623 23069 39635 23072
rect 39577 23063 39635 23069
rect 39758 23060 39764 23072
rect 39816 23060 39822 23112
rect 36357 23035 36415 23041
rect 36357 23001 36369 23035
rect 36403 23032 36415 23035
rect 37366 23032 37372 23044
rect 36403 23004 37372 23032
rect 36403 23001 36415 23004
rect 36357 22995 36415 23001
rect 37366 22992 37372 23004
rect 37424 22992 37430 23044
rect 38654 22992 38660 23044
rect 38712 23032 38718 23044
rect 38749 23035 38807 23041
rect 38749 23032 38761 23035
rect 38712 23004 38761 23032
rect 38712 22992 38718 23004
rect 38749 23001 38761 23004
rect 38795 23001 38807 23035
rect 38749 22995 38807 23001
rect 35952 22936 36216 22964
rect 36725 22967 36783 22973
rect 35952 22924 35958 22936
rect 36725 22933 36737 22967
rect 36771 22964 36783 22967
rect 38010 22964 38016 22976
rect 36771 22936 38016 22964
rect 36771 22933 36783 22936
rect 36725 22927 36783 22933
rect 38010 22924 38016 22936
rect 38068 22924 38074 22976
rect 1104 22874 40572 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 40572 22874
rect 1104 22800 40572 22822
rect 2590 22720 2596 22772
rect 2648 22720 2654 22772
rect 2685 22763 2743 22769
rect 2685 22729 2697 22763
rect 2731 22760 2743 22763
rect 3050 22760 3056 22772
rect 2731 22732 3056 22760
rect 2731 22729 2743 22732
rect 2685 22723 2743 22729
rect 3050 22720 3056 22732
rect 3108 22720 3114 22772
rect 6181 22763 6239 22769
rect 6181 22729 6193 22763
rect 6227 22760 6239 22763
rect 6730 22760 6736 22772
rect 6227 22732 6736 22760
rect 6227 22729 6239 22732
rect 6181 22723 6239 22729
rect 6730 22720 6736 22732
rect 6788 22720 6794 22772
rect 8110 22720 8116 22772
rect 8168 22760 8174 22772
rect 9306 22760 9312 22772
rect 8168 22732 9312 22760
rect 8168 22720 8174 22732
rect 9306 22720 9312 22732
rect 9364 22720 9370 22772
rect 11885 22763 11943 22769
rect 11885 22729 11897 22763
rect 11931 22760 11943 22763
rect 12342 22760 12348 22772
rect 11931 22732 12348 22760
rect 11931 22729 11943 22732
rect 11885 22723 11943 22729
rect 12342 22720 12348 22732
rect 12400 22720 12406 22772
rect 12618 22720 12624 22772
rect 12676 22760 12682 22772
rect 13630 22760 13636 22772
rect 12676 22732 13636 22760
rect 12676 22720 12682 22732
rect 13630 22720 13636 22732
rect 13688 22760 13694 22772
rect 14274 22760 14280 22772
rect 13688 22732 14280 22760
rect 13688 22720 13694 22732
rect 14274 22720 14280 22732
rect 14332 22720 14338 22772
rect 18046 22720 18052 22772
rect 18104 22760 18110 22772
rect 18230 22760 18236 22772
rect 18104 22732 18236 22760
rect 18104 22720 18110 22732
rect 18230 22720 18236 22732
rect 18288 22760 18294 22772
rect 18598 22760 18604 22772
rect 18288 22732 18604 22760
rect 18288 22720 18294 22732
rect 18598 22720 18604 22732
rect 18656 22720 18662 22772
rect 20346 22720 20352 22772
rect 20404 22720 20410 22772
rect 20622 22720 20628 22772
rect 20680 22760 20686 22772
rect 21269 22763 21327 22769
rect 21269 22760 21281 22763
rect 20680 22732 21281 22760
rect 20680 22720 20686 22732
rect 21269 22729 21281 22732
rect 21315 22760 21327 22763
rect 21315 22732 22094 22760
rect 21315 22729 21327 22732
rect 21269 22723 21327 22729
rect 4706 22692 4712 22704
rect 4554 22678 4712 22692
rect 4540 22664 4712 22678
rect 2866 22584 2872 22636
rect 2924 22624 2930 22636
rect 3053 22627 3111 22633
rect 3053 22624 3065 22627
rect 2924 22596 3065 22624
rect 2924 22584 2930 22596
rect 3053 22593 3065 22596
rect 3099 22593 3111 22627
rect 3053 22587 3111 22593
rect 2777 22559 2835 22565
rect 2777 22525 2789 22559
rect 2823 22556 2835 22559
rect 2823 22528 2912 22556
rect 2823 22525 2835 22528
rect 2777 22519 2835 22525
rect 2884 22500 2912 22528
rect 3326 22516 3332 22568
rect 3384 22516 3390 22568
rect 3786 22516 3792 22568
rect 3844 22556 3850 22568
rect 4540 22556 4568 22664
rect 4706 22652 4712 22664
rect 4764 22652 4770 22704
rect 5813 22695 5871 22701
rect 5813 22661 5825 22695
rect 5859 22692 5871 22695
rect 5859 22664 6224 22692
rect 5859 22661 5871 22664
rect 5813 22655 5871 22661
rect 6196 22636 6224 22664
rect 8018 22652 8024 22704
rect 8076 22692 8082 22704
rect 8076 22664 8800 22692
rect 8076 22652 8082 22664
rect 5629 22627 5687 22633
rect 5629 22593 5641 22627
rect 5675 22624 5687 22627
rect 5718 22624 5724 22636
rect 5675 22596 5724 22624
rect 5675 22593 5687 22596
rect 5629 22587 5687 22593
rect 5718 22584 5724 22596
rect 5776 22584 5782 22636
rect 5905 22627 5963 22633
rect 5905 22593 5917 22627
rect 5951 22593 5963 22627
rect 5905 22587 5963 22593
rect 5997 22627 6055 22633
rect 5997 22593 6009 22627
rect 6043 22593 6055 22627
rect 5997 22587 6055 22593
rect 3844 22528 4568 22556
rect 4801 22559 4859 22565
rect 3844 22516 3850 22528
rect 4801 22525 4813 22559
rect 4847 22556 4859 22559
rect 5445 22559 5503 22565
rect 5445 22556 5457 22559
rect 4847 22528 5457 22556
rect 4847 22525 4859 22528
rect 4801 22519 4859 22525
rect 5445 22525 5457 22528
rect 5491 22556 5503 22559
rect 5920 22556 5948 22587
rect 5491 22528 5948 22556
rect 6012 22556 6040 22587
rect 6178 22584 6184 22636
rect 6236 22584 6242 22636
rect 8481 22627 8539 22633
rect 8481 22593 8493 22627
rect 8527 22593 8539 22627
rect 8481 22587 8539 22593
rect 6730 22556 6736 22568
rect 6012 22528 6736 22556
rect 5491 22525 5503 22528
rect 5445 22519 5503 22525
rect 2866 22448 2872 22500
rect 2924 22448 2930 22500
rect 4706 22448 4712 22500
rect 4764 22488 4770 22500
rect 4893 22491 4951 22497
rect 4893 22488 4905 22491
rect 4764 22460 4905 22488
rect 4764 22448 4770 22460
rect 4893 22457 4905 22460
rect 4939 22457 4951 22491
rect 4893 22451 4951 22457
rect 5258 22448 5264 22500
rect 5316 22488 5322 22500
rect 6012 22488 6040 22528
rect 6730 22516 6736 22528
rect 6788 22516 6794 22568
rect 8496 22556 8524 22587
rect 8570 22584 8576 22636
rect 8628 22624 8634 22636
rect 8772 22633 8800 22664
rect 10502 22652 10508 22704
rect 10560 22692 10566 22704
rect 10560 22664 11192 22692
rect 10560 22652 10566 22664
rect 8665 22627 8723 22633
rect 8665 22624 8677 22627
rect 8628 22596 8677 22624
rect 8628 22584 8634 22596
rect 8665 22593 8677 22596
rect 8711 22593 8723 22627
rect 8665 22587 8723 22593
rect 8757 22627 8815 22633
rect 8757 22593 8769 22627
rect 8803 22593 8815 22627
rect 8757 22587 8815 22593
rect 10226 22584 10232 22636
rect 10284 22624 10290 22636
rect 10781 22627 10839 22633
rect 10781 22624 10793 22627
rect 10284 22596 10793 22624
rect 10284 22584 10290 22596
rect 10781 22593 10793 22596
rect 10827 22593 10839 22627
rect 10781 22587 10839 22593
rect 10870 22584 10876 22636
rect 10928 22584 10934 22636
rect 11164 22633 11192 22664
rect 11330 22652 11336 22704
rect 11388 22692 11394 22704
rect 11388 22664 12480 22692
rect 11388 22652 11394 22664
rect 11149 22627 11207 22633
rect 11149 22593 11161 22627
rect 11195 22624 11207 22627
rect 11195 22596 11744 22624
rect 11195 22593 11207 22596
rect 11149 22587 11207 22593
rect 8496 22528 8708 22556
rect 5316 22460 6040 22488
rect 5316 22448 5322 22460
rect 8570 22448 8576 22500
rect 8628 22448 8634 22500
rect 8680 22488 8708 22528
rect 9490 22516 9496 22568
rect 9548 22516 9554 22568
rect 11606 22556 11612 22568
rect 9600 22528 11612 22556
rect 9600 22488 9628 22528
rect 11606 22516 11612 22528
rect 11664 22516 11670 22568
rect 11716 22565 11744 22596
rect 11974 22584 11980 22636
rect 12032 22584 12038 22636
rect 12452 22633 12480 22664
rect 14182 22652 14188 22704
rect 14240 22652 14246 22704
rect 20364 22692 20392 22720
rect 20364 22664 20668 22692
rect 12437 22627 12495 22633
rect 12437 22593 12449 22627
rect 12483 22624 12495 22627
rect 13998 22624 14004 22636
rect 12483 22596 14004 22624
rect 12483 22593 12495 22596
rect 12437 22587 12495 22593
rect 13998 22584 14004 22596
rect 14056 22584 14062 22636
rect 19334 22584 19340 22636
rect 19392 22624 19398 22636
rect 19886 22624 19892 22636
rect 19392 22596 19892 22624
rect 19392 22584 19398 22596
rect 19886 22584 19892 22596
rect 19944 22584 19950 22636
rect 20346 22584 20352 22636
rect 20404 22584 20410 22636
rect 20640 22633 20668 22664
rect 21450 22652 21456 22704
rect 21508 22652 21514 22704
rect 22066 22692 22094 22732
rect 22186 22720 22192 22772
rect 22244 22760 22250 22772
rect 22922 22760 22928 22772
rect 22244 22732 22928 22760
rect 22244 22720 22250 22732
rect 22922 22720 22928 22732
rect 22980 22720 22986 22772
rect 25406 22720 25412 22772
rect 25464 22720 25470 22772
rect 25682 22720 25688 22772
rect 25740 22760 25746 22772
rect 26418 22760 26424 22772
rect 25740 22732 26424 22760
rect 25740 22720 25746 22732
rect 26418 22720 26424 22732
rect 26476 22720 26482 22772
rect 27522 22720 27528 22772
rect 27580 22720 27586 22772
rect 27614 22720 27620 22772
rect 27672 22760 27678 22772
rect 27672 22732 29408 22760
rect 27672 22720 27678 22732
rect 22066 22664 24348 22692
rect 20441 22627 20499 22633
rect 20441 22593 20453 22627
rect 20487 22593 20499 22627
rect 20441 22587 20499 22593
rect 20625 22627 20683 22633
rect 20625 22593 20637 22627
rect 20671 22593 20683 22627
rect 20625 22587 20683 22593
rect 20717 22627 20775 22633
rect 20717 22593 20729 22627
rect 20763 22624 20775 22627
rect 20806 22624 20812 22636
rect 20763 22596 20812 22624
rect 20763 22593 20775 22596
rect 20717 22587 20775 22593
rect 11701 22559 11759 22565
rect 11701 22525 11713 22559
rect 11747 22556 11759 22559
rect 12158 22556 12164 22568
rect 11747 22528 12164 22556
rect 11747 22525 11759 22528
rect 11701 22519 11759 22525
rect 12158 22516 12164 22528
rect 12216 22556 12222 22568
rect 12529 22559 12587 22565
rect 12529 22556 12541 22559
rect 12216 22528 12541 22556
rect 12216 22516 12222 22528
rect 12529 22525 12541 22528
rect 12575 22556 12587 22559
rect 12986 22556 12992 22568
rect 12575 22528 12992 22556
rect 12575 22525 12587 22528
rect 12529 22519 12587 22525
rect 12986 22516 12992 22528
rect 13044 22516 13050 22568
rect 14016 22556 14044 22584
rect 14016 22528 20116 22556
rect 8680 22460 9628 22488
rect 9968 22460 10180 22488
rect 2222 22380 2228 22432
rect 2280 22380 2286 22432
rect 3878 22380 3884 22432
rect 3936 22420 3942 22432
rect 5276 22420 5304 22448
rect 3936 22392 5304 22420
rect 3936 22380 3942 22392
rect 5626 22380 5632 22432
rect 5684 22420 5690 22432
rect 7834 22420 7840 22432
rect 5684 22392 7840 22420
rect 5684 22380 5690 22392
rect 7834 22380 7840 22392
rect 7892 22420 7898 22432
rect 8680 22420 8708 22460
rect 7892 22392 8708 22420
rect 7892 22380 7898 22392
rect 8938 22380 8944 22432
rect 8996 22380 9002 22432
rect 9030 22380 9036 22432
rect 9088 22420 9094 22432
rect 9582 22420 9588 22432
rect 9088 22392 9588 22420
rect 9088 22380 9094 22392
rect 9582 22380 9588 22392
rect 9640 22420 9646 22432
rect 9968 22420 9996 22460
rect 9640 22392 9996 22420
rect 9640 22380 9646 22392
rect 10042 22380 10048 22432
rect 10100 22380 10106 22432
rect 10152 22420 10180 22460
rect 10226 22448 10232 22500
rect 10284 22488 10290 22500
rect 10597 22491 10655 22497
rect 10597 22488 10609 22491
rect 10284 22460 10609 22488
rect 10284 22448 10290 22460
rect 10597 22457 10609 22460
rect 10643 22457 10655 22491
rect 10597 22451 10655 22457
rect 16942 22448 16948 22500
rect 17000 22488 17006 22500
rect 19978 22488 19984 22500
rect 17000 22460 19984 22488
rect 17000 22448 17006 22460
rect 19978 22448 19984 22460
rect 20036 22448 20042 22500
rect 20088 22488 20116 22528
rect 20162 22516 20168 22568
rect 20220 22556 20226 22568
rect 20456 22556 20484 22587
rect 20220 22528 20484 22556
rect 20220 22516 20226 22528
rect 20438 22488 20444 22500
rect 20088 22460 20444 22488
rect 20438 22448 20444 22460
rect 20496 22448 20502 22500
rect 11057 22423 11115 22429
rect 11057 22420 11069 22423
rect 10152 22392 11069 22420
rect 11057 22389 11069 22392
rect 11103 22389 11115 22423
rect 11057 22383 11115 22389
rect 12158 22380 12164 22432
rect 12216 22420 12222 22432
rect 12345 22423 12403 22429
rect 12345 22420 12357 22423
rect 12216 22392 12357 22420
rect 12216 22380 12222 22392
rect 12345 22389 12357 22392
rect 12391 22389 12403 22423
rect 12345 22383 12403 22389
rect 13817 22423 13875 22429
rect 13817 22389 13829 22423
rect 13863 22420 13875 22423
rect 14550 22420 14556 22432
rect 13863 22392 14556 22420
rect 13863 22389 13875 22392
rect 13817 22383 13875 22389
rect 14550 22380 14556 22392
rect 14608 22380 14614 22432
rect 16482 22380 16488 22432
rect 16540 22420 16546 22432
rect 20732 22420 20760 22587
rect 20806 22584 20812 22596
rect 20864 22584 20870 22636
rect 21468 22624 21496 22652
rect 24320 22636 24348 22664
rect 25314 22652 25320 22704
rect 25372 22692 25378 22704
rect 28169 22695 28227 22701
rect 28169 22692 28181 22695
rect 25372 22664 28181 22692
rect 25372 22652 25378 22664
rect 28169 22661 28181 22664
rect 28215 22692 28227 22695
rect 29273 22695 29331 22701
rect 28215 22664 29224 22692
rect 28215 22661 28227 22664
rect 28169 22655 28227 22661
rect 23750 22624 23756 22636
rect 21468 22596 23756 22624
rect 23750 22584 23756 22596
rect 23808 22584 23814 22636
rect 24026 22584 24032 22636
rect 24084 22584 24090 22636
rect 24118 22584 24124 22636
rect 24176 22584 24182 22636
rect 24302 22584 24308 22636
rect 24360 22584 24366 22636
rect 24397 22627 24455 22633
rect 24397 22593 24409 22627
rect 24443 22624 24455 22627
rect 24486 22624 24492 22636
rect 24443 22596 24492 22624
rect 24443 22593 24455 22596
rect 24397 22587 24455 22593
rect 24412 22556 24440 22587
rect 24486 22584 24492 22596
rect 24544 22624 24550 22636
rect 24946 22624 24952 22636
rect 24544 22596 24952 22624
rect 24544 22584 24550 22596
rect 24946 22584 24952 22596
rect 25004 22584 25010 22636
rect 25568 22627 25626 22633
rect 25568 22593 25580 22627
rect 25614 22624 25626 22627
rect 26145 22627 26203 22633
rect 26145 22624 26157 22627
rect 25614 22596 26157 22624
rect 25614 22593 25626 22596
rect 25568 22587 25626 22593
rect 26145 22593 26157 22596
rect 26191 22593 26203 22627
rect 26145 22587 26203 22593
rect 26326 22584 26332 22636
rect 26384 22624 26390 22636
rect 26605 22627 26663 22633
rect 26605 22624 26617 22627
rect 26384 22596 26617 22624
rect 26384 22584 26390 22596
rect 26605 22593 26617 22596
rect 26651 22593 26663 22627
rect 26605 22587 26663 22593
rect 26697 22627 26755 22633
rect 26697 22593 26709 22627
rect 26743 22593 26755 22627
rect 26697 22587 26755 22593
rect 21284 22528 24440 22556
rect 25777 22559 25835 22565
rect 21284 22432 21312 22528
rect 25777 22525 25789 22559
rect 25823 22556 25835 22559
rect 25866 22556 25872 22568
rect 25823 22528 25872 22556
rect 25823 22525 25835 22528
rect 25777 22519 25835 22525
rect 25866 22516 25872 22528
rect 25924 22516 25930 22568
rect 25958 22516 25964 22568
rect 26016 22556 26022 22568
rect 26053 22559 26111 22565
rect 26053 22556 26065 22559
rect 26016 22528 26065 22556
rect 26016 22516 26022 22528
rect 26053 22525 26065 22528
rect 26099 22525 26111 22559
rect 26053 22519 26111 22525
rect 26421 22559 26479 22565
rect 26421 22525 26433 22559
rect 26467 22556 26479 22559
rect 26510 22556 26516 22568
rect 26467 22528 26516 22556
rect 26467 22525 26479 22528
rect 26421 22519 26479 22525
rect 26510 22516 26516 22528
rect 26568 22516 26574 22568
rect 23290 22448 23296 22500
rect 23348 22488 23354 22500
rect 26329 22491 26387 22497
rect 26329 22488 26341 22491
rect 23348 22460 26341 22488
rect 23348 22448 23354 22460
rect 26329 22457 26341 22460
rect 26375 22457 26387 22491
rect 26712 22488 26740 22587
rect 26786 22584 26792 22636
rect 26844 22624 26850 22636
rect 27709 22627 27767 22633
rect 27709 22624 27721 22627
rect 26844 22596 27721 22624
rect 26844 22584 26850 22596
rect 27709 22593 27721 22596
rect 27755 22593 27767 22627
rect 27709 22587 27767 22593
rect 28442 22584 28448 22636
rect 28500 22624 28506 22636
rect 28626 22624 28632 22636
rect 28500 22596 28632 22624
rect 28500 22584 28506 22596
rect 28626 22584 28632 22596
rect 28684 22584 28690 22636
rect 28902 22633 28908 22636
rect 28900 22587 28908 22633
rect 28902 22584 28908 22587
rect 28960 22584 28966 22636
rect 28994 22584 29000 22636
rect 29052 22584 29058 22636
rect 29089 22627 29147 22633
rect 29089 22593 29101 22627
rect 29135 22593 29147 22627
rect 29089 22587 29147 22593
rect 27893 22559 27951 22565
rect 27893 22525 27905 22559
rect 27939 22556 27951 22559
rect 28261 22559 28319 22565
rect 28261 22556 28273 22559
rect 27939 22528 28273 22556
rect 27939 22525 27951 22528
rect 27893 22519 27951 22525
rect 28261 22525 28273 22528
rect 28307 22525 28319 22559
rect 28261 22519 28319 22525
rect 28718 22516 28724 22568
rect 28776 22516 28782 22568
rect 26329 22451 26387 22457
rect 26436 22460 26740 22488
rect 16540 22392 20760 22420
rect 16540 22380 16546 22392
rect 20898 22380 20904 22432
rect 20956 22380 20962 22432
rect 21082 22380 21088 22432
rect 21140 22380 21146 22432
rect 21266 22380 21272 22432
rect 21324 22380 21330 22432
rect 24489 22423 24547 22429
rect 24489 22389 24501 22423
rect 24535 22420 24547 22423
rect 24670 22420 24676 22432
rect 24535 22392 24676 22420
rect 24535 22389 24547 22392
rect 24489 22383 24547 22389
rect 24670 22380 24676 22392
rect 24728 22380 24734 22432
rect 25682 22380 25688 22432
rect 25740 22420 25746 22432
rect 26436 22420 26464 22460
rect 27062 22448 27068 22500
rect 27120 22488 27126 22500
rect 28166 22488 28172 22500
rect 27120 22460 28172 22488
rect 27120 22448 27126 22460
rect 28166 22448 28172 22460
rect 28224 22488 28230 22500
rect 28629 22491 28687 22497
rect 28629 22488 28641 22491
rect 28224 22460 28641 22488
rect 28224 22448 28230 22460
rect 28629 22457 28641 22460
rect 28675 22488 28687 22491
rect 29104 22488 29132 22587
rect 29196 22565 29224 22664
rect 29273 22661 29285 22695
rect 29319 22692 29331 22695
rect 29380 22692 29408 22732
rect 29638 22720 29644 22772
rect 29696 22720 29702 22772
rect 30190 22720 30196 22772
rect 30248 22760 30254 22772
rect 30653 22763 30711 22769
rect 30653 22760 30665 22763
rect 30248 22732 30665 22760
rect 30248 22720 30254 22732
rect 30653 22729 30665 22732
rect 30699 22729 30711 22763
rect 31846 22760 31852 22772
rect 30653 22723 30711 22729
rect 31588 22732 31852 22760
rect 31588 22701 31616 22732
rect 31846 22720 31852 22732
rect 31904 22720 31910 22772
rect 32030 22720 32036 22772
rect 32088 22760 32094 22772
rect 32677 22763 32735 22769
rect 32677 22760 32689 22763
rect 32088 22732 32689 22760
rect 32088 22720 32094 22732
rect 32677 22729 32689 22732
rect 32723 22729 32735 22763
rect 36262 22760 36268 22772
rect 32677 22723 32735 22729
rect 36096 22732 36268 22760
rect 31573 22695 31631 22701
rect 29319 22664 31524 22692
rect 29319 22661 29331 22664
rect 29273 22655 29331 22661
rect 29454 22584 29460 22636
rect 29512 22624 29518 22636
rect 29825 22627 29883 22633
rect 29825 22624 29837 22627
rect 29512 22596 29837 22624
rect 29512 22584 29518 22596
rect 29825 22593 29837 22596
rect 29871 22593 29883 22627
rect 29825 22587 29883 22593
rect 29181 22559 29239 22565
rect 29181 22525 29193 22559
rect 29227 22525 29239 22559
rect 29840 22556 29868 22587
rect 29914 22584 29920 22636
rect 29972 22584 29978 22636
rect 30285 22627 30343 22633
rect 30285 22593 30297 22627
rect 30331 22593 30343 22627
rect 30285 22587 30343 22593
rect 30300 22556 30328 22587
rect 30374 22584 30380 22636
rect 30432 22584 30438 22636
rect 30837 22627 30895 22633
rect 30837 22593 30849 22627
rect 30883 22593 30895 22627
rect 30837 22587 30895 22593
rect 30558 22556 30564 22568
rect 29840 22528 30564 22556
rect 29181 22519 29239 22525
rect 30558 22516 30564 22528
rect 30616 22516 30622 22568
rect 30852 22556 30880 22587
rect 31386 22584 31392 22636
rect 31444 22584 31450 22636
rect 31496 22624 31524 22664
rect 31573 22661 31585 22695
rect 31619 22661 31631 22695
rect 31573 22655 31631 22661
rect 32232 22664 33180 22692
rect 31662 22624 31668 22636
rect 31496 22596 31668 22624
rect 31662 22584 31668 22596
rect 31720 22584 31726 22636
rect 31754 22584 31760 22636
rect 31812 22584 31818 22636
rect 31846 22584 31852 22636
rect 31904 22624 31910 22636
rect 32125 22627 32183 22633
rect 32125 22624 32137 22627
rect 31904 22596 32137 22624
rect 31904 22584 31910 22596
rect 32125 22593 32137 22596
rect 32171 22593 32183 22627
rect 32125 22587 32183 22593
rect 31570 22556 31576 22568
rect 30852 22528 31576 22556
rect 31570 22516 31576 22528
rect 31628 22516 31634 22568
rect 31772 22556 31800 22584
rect 32232 22556 32260 22664
rect 32309 22627 32367 22633
rect 32309 22593 32321 22627
rect 32355 22593 32367 22627
rect 32309 22587 32367 22593
rect 31772 22528 32260 22556
rect 32324 22556 32352 22587
rect 32398 22584 32404 22636
rect 32456 22584 32462 22636
rect 32508 22633 32536 22664
rect 32493 22627 32551 22633
rect 32493 22593 32505 22627
rect 32539 22593 32551 22627
rect 32493 22587 32551 22593
rect 32858 22584 32864 22636
rect 32916 22584 32922 22636
rect 33042 22584 33048 22636
rect 33100 22584 33106 22636
rect 32674 22556 32680 22568
rect 32324 22528 32680 22556
rect 32674 22516 32680 22528
rect 32732 22516 32738 22568
rect 33152 22565 33180 22664
rect 34422 22652 34428 22704
rect 34480 22692 34486 22704
rect 36096 22701 36124 22732
rect 36262 22720 36268 22732
rect 36320 22720 36326 22772
rect 36081 22695 36139 22701
rect 34480 22664 35940 22692
rect 34480 22652 34486 22664
rect 33410 22584 33416 22636
rect 33468 22624 33474 22636
rect 33870 22624 33876 22636
rect 33468 22596 33876 22624
rect 33468 22584 33474 22596
rect 33870 22584 33876 22596
rect 33928 22584 33934 22636
rect 35434 22584 35440 22636
rect 35492 22624 35498 22636
rect 35912 22633 35940 22664
rect 36081 22661 36093 22695
rect 36127 22661 36139 22695
rect 36081 22655 36139 22661
rect 35805 22627 35863 22633
rect 35805 22624 35817 22627
rect 35492 22596 35817 22624
rect 35492 22584 35498 22596
rect 35805 22593 35817 22596
rect 35851 22593 35863 22627
rect 35805 22587 35863 22593
rect 35898 22627 35956 22633
rect 35898 22593 35910 22627
rect 35944 22593 35956 22627
rect 35898 22587 35956 22593
rect 36170 22584 36176 22636
rect 36228 22584 36234 22636
rect 36311 22627 36369 22633
rect 36311 22593 36323 22627
rect 36357 22624 36369 22627
rect 36538 22624 36544 22636
rect 36357 22596 36544 22624
rect 36357 22593 36369 22596
rect 36311 22587 36369 22593
rect 36538 22584 36544 22596
rect 36596 22584 36602 22636
rect 38010 22584 38016 22636
rect 38068 22584 38074 22636
rect 32953 22559 33011 22565
rect 32953 22556 32965 22559
rect 32784 22528 32965 22556
rect 30282 22488 30288 22500
rect 28675 22460 29132 22488
rect 29748 22460 30288 22488
rect 28675 22457 28687 22460
rect 28629 22451 28687 22457
rect 25740 22392 26464 22420
rect 26513 22423 26571 22429
rect 25740 22380 25746 22392
rect 26513 22389 26525 22423
rect 26559 22420 26571 22423
rect 27338 22420 27344 22432
rect 26559 22392 27344 22420
rect 26559 22389 26571 22392
rect 26513 22383 26571 22389
rect 27338 22380 27344 22392
rect 27396 22380 27402 22432
rect 27614 22380 27620 22432
rect 27672 22420 27678 22432
rect 28074 22420 28080 22432
rect 27672 22392 28080 22420
rect 27672 22380 27678 22392
rect 28074 22380 28080 22392
rect 28132 22380 28138 22432
rect 28442 22380 28448 22432
rect 28500 22420 28506 22432
rect 29748 22420 29776 22460
rect 30282 22448 30288 22460
rect 30340 22448 30346 22500
rect 30576 22488 30604 22516
rect 31941 22491 31999 22497
rect 30576 22460 31616 22488
rect 28500 22392 29776 22420
rect 28500 22380 28506 22392
rect 30006 22380 30012 22432
rect 30064 22420 30070 22432
rect 30101 22423 30159 22429
rect 30101 22420 30113 22423
rect 30064 22392 30113 22420
rect 30064 22380 30070 22392
rect 30101 22389 30113 22392
rect 30147 22420 30159 22423
rect 31294 22420 31300 22432
rect 30147 22392 31300 22420
rect 30147 22389 30159 22392
rect 30101 22383 30159 22389
rect 31294 22380 31300 22392
rect 31352 22380 31358 22432
rect 31588 22420 31616 22460
rect 31941 22457 31953 22491
rect 31987 22488 31999 22491
rect 32122 22488 32128 22500
rect 31987 22460 32128 22488
rect 31987 22457 31999 22460
rect 31941 22451 31999 22457
rect 32122 22448 32128 22460
rect 32180 22448 32186 22500
rect 32784 22488 32812 22528
rect 32953 22525 32965 22528
rect 32999 22525 33011 22559
rect 32953 22519 33011 22525
rect 33137 22559 33195 22565
rect 33137 22525 33149 22559
rect 33183 22556 33195 22559
rect 34790 22556 34796 22568
rect 33183 22528 34796 22556
rect 33183 22525 33195 22528
rect 33137 22519 33195 22525
rect 34790 22516 34796 22528
rect 34848 22516 34854 22568
rect 37918 22516 37924 22568
rect 37976 22556 37982 22568
rect 38105 22559 38163 22565
rect 38105 22556 38117 22559
rect 37976 22528 38117 22556
rect 37976 22516 37982 22528
rect 38105 22525 38117 22528
rect 38151 22556 38163 22559
rect 38378 22556 38384 22568
rect 38151 22528 38384 22556
rect 38151 22525 38163 22528
rect 38105 22519 38163 22525
rect 38378 22516 38384 22528
rect 38436 22516 38442 22568
rect 32858 22488 32864 22500
rect 32784 22460 32864 22488
rect 32858 22448 32864 22460
rect 32916 22448 32922 22500
rect 33321 22491 33379 22497
rect 33321 22457 33333 22491
rect 33367 22488 33379 22491
rect 37458 22488 37464 22500
rect 33367 22460 37464 22488
rect 33367 22457 33379 22460
rect 33321 22451 33379 22457
rect 37458 22448 37464 22460
rect 37516 22488 37522 22500
rect 37516 22460 38056 22488
rect 37516 22448 37522 22460
rect 33042 22420 33048 22432
rect 31588 22392 33048 22420
rect 33042 22380 33048 22392
rect 33100 22380 33106 22432
rect 36449 22423 36507 22429
rect 36449 22389 36461 22423
rect 36495 22420 36507 22423
rect 37918 22420 37924 22432
rect 36495 22392 37924 22420
rect 36495 22389 36507 22392
rect 36449 22383 36507 22389
rect 37918 22380 37924 22392
rect 37976 22380 37982 22432
rect 38028 22429 38056 22460
rect 38013 22423 38071 22429
rect 38013 22389 38025 22423
rect 38059 22389 38071 22423
rect 38013 22383 38071 22389
rect 38381 22423 38439 22429
rect 38381 22389 38393 22423
rect 38427 22420 38439 22423
rect 39758 22420 39764 22432
rect 38427 22392 39764 22420
rect 38427 22389 38439 22392
rect 38381 22383 38439 22389
rect 39758 22380 39764 22392
rect 39816 22380 39822 22432
rect 1104 22330 40572 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 40572 22330
rect 1104 22256 40572 22278
rect 1752 22219 1810 22225
rect 1752 22185 1764 22219
rect 1798 22216 1810 22219
rect 2222 22216 2228 22228
rect 1798 22188 2228 22216
rect 1798 22185 1810 22188
rect 1752 22179 1810 22185
rect 2222 22176 2228 22188
rect 2280 22176 2286 22228
rect 3234 22176 3240 22228
rect 3292 22176 3298 22228
rect 6288 22188 6914 22216
rect 6288 22148 6316 22188
rect 6454 22148 6460 22160
rect 6196 22120 6316 22148
rect 6380 22120 6460 22148
rect 1486 21972 1492 22024
rect 1544 21972 1550 22024
rect 3050 22012 3056 22024
rect 2898 21984 3056 22012
rect 3050 21972 3056 21984
rect 3108 22012 3114 22024
rect 3786 22012 3792 22024
rect 3108 21984 3792 22012
rect 3108 21972 3114 21984
rect 3786 21972 3792 21984
rect 3844 21972 3850 22024
rect 4341 22015 4399 22021
rect 4341 21981 4353 22015
rect 4387 22012 4399 22015
rect 4614 22012 4620 22024
rect 4387 21984 4620 22012
rect 4387 21981 4399 21984
rect 4341 21975 4399 21981
rect 4614 21972 4620 21984
rect 4672 21972 4678 22024
rect 5626 21972 5632 22024
rect 5684 22012 5690 22024
rect 6196 22021 6224 22120
rect 5905 22015 5963 22021
rect 5905 22012 5917 22015
rect 5684 21984 5917 22012
rect 5684 21972 5690 21984
rect 5905 21981 5917 21984
rect 5951 21981 5963 22015
rect 5905 21975 5963 21981
rect 6181 22015 6239 22021
rect 6181 21981 6193 22015
rect 6227 21981 6239 22015
rect 6181 21975 6239 21981
rect 5169 21947 5227 21953
rect 5169 21913 5181 21947
rect 5215 21944 5227 21947
rect 5442 21944 5448 21956
rect 5215 21916 5448 21944
rect 5215 21913 5227 21916
rect 5169 21907 5227 21913
rect 5442 21904 5448 21916
rect 5500 21904 5506 21956
rect 5718 21904 5724 21956
rect 5776 21944 5782 21956
rect 6196 21944 6224 21975
rect 6270 21972 6276 22024
rect 6328 21972 6334 22024
rect 6380 22021 6408 22120
rect 6454 22108 6460 22120
rect 6512 22108 6518 22160
rect 6886 22080 6914 22188
rect 8570 22176 8576 22228
rect 8628 22216 8634 22228
rect 8665 22219 8723 22225
rect 8665 22216 8677 22219
rect 8628 22188 8677 22216
rect 8628 22176 8634 22188
rect 8665 22185 8677 22188
rect 8711 22185 8723 22219
rect 8665 22179 8723 22185
rect 8938 22176 8944 22228
rect 8996 22216 9002 22228
rect 8996 22188 11652 22216
rect 8996 22176 9002 22188
rect 7285 22151 7343 22157
rect 7285 22117 7297 22151
rect 7331 22148 7343 22151
rect 8202 22148 8208 22160
rect 7331 22120 8208 22148
rect 7331 22117 7343 22120
rect 7285 22111 7343 22117
rect 8202 22108 8208 22120
rect 8260 22108 8266 22160
rect 11238 22148 11244 22160
rect 10704 22120 11244 22148
rect 10410 22080 10416 22092
rect 6886 22052 7420 22080
rect 6365 22015 6423 22021
rect 6365 21981 6377 22015
rect 6411 21981 6423 22015
rect 6365 21975 6423 21981
rect 6454 21972 6460 22024
rect 6512 21972 6518 22024
rect 7006 21972 7012 22024
rect 7064 21972 7070 22024
rect 7392 22021 7420 22052
rect 7944 22052 10416 22080
rect 7193 22015 7251 22021
rect 7193 21981 7205 22015
rect 7239 21981 7251 22015
rect 7193 21975 7251 21981
rect 7377 22015 7435 22021
rect 7377 21981 7389 22015
rect 7423 22012 7435 22015
rect 7834 22012 7840 22024
rect 7423 21984 7840 22012
rect 7423 21981 7435 21984
rect 7377 21975 7435 21981
rect 5776 21916 6224 21944
rect 5776 21904 5782 21916
rect 7098 21904 7104 21956
rect 7156 21944 7162 21956
rect 7208 21944 7236 21975
rect 7834 21972 7840 21984
rect 7892 21972 7898 22024
rect 7944 21944 7972 22052
rect 10410 22040 10416 22052
rect 10468 22040 10474 22092
rect 10704 22089 10732 22120
rect 11238 22108 11244 22120
rect 11296 22108 11302 22160
rect 11514 22108 11520 22160
rect 11572 22108 11578 22160
rect 11624 22148 11652 22188
rect 12066 22176 12072 22228
rect 12124 22216 12130 22228
rect 18230 22216 18236 22228
rect 12124 22188 14412 22216
rect 12124 22176 12130 22188
rect 12618 22148 12624 22160
rect 11624 22120 12624 22148
rect 12618 22108 12624 22120
rect 12676 22108 12682 22160
rect 14384 22157 14412 22188
rect 17788 22188 18236 22216
rect 14369 22151 14427 22157
rect 12820 22120 13032 22148
rect 10689 22083 10747 22089
rect 10689 22049 10701 22083
rect 10735 22049 10747 22083
rect 10689 22043 10747 22049
rect 12437 22083 12495 22089
rect 12437 22049 12449 22083
rect 12483 22080 12495 22083
rect 12820 22080 12848 22120
rect 12483 22052 12848 22080
rect 12483 22049 12495 22052
rect 12437 22043 12495 22049
rect 12894 22040 12900 22092
rect 12952 22040 12958 22092
rect 13004 22080 13032 22120
rect 14369 22117 14381 22151
rect 14415 22117 14427 22151
rect 14369 22111 14427 22117
rect 13817 22083 13875 22089
rect 13817 22080 13829 22083
rect 13004 22052 13124 22080
rect 13096 22024 13124 22052
rect 13280 22052 13829 22080
rect 8110 21972 8116 22024
rect 8168 21972 8174 22024
rect 8478 21972 8484 22024
rect 8536 21972 8542 22024
rect 10781 22015 10839 22021
rect 10781 21981 10793 22015
rect 10827 21981 10839 22015
rect 10781 21975 10839 21981
rect 7156 21916 7972 21944
rect 7156 21904 7162 21916
rect 8294 21904 8300 21956
rect 8352 21904 8358 21956
rect 8389 21947 8447 21953
rect 8389 21913 8401 21947
rect 8435 21944 8447 21947
rect 8570 21944 8576 21956
rect 8435 21916 8576 21944
rect 8435 21913 8447 21916
rect 8389 21907 8447 21913
rect 8570 21904 8576 21916
rect 8628 21904 8634 21956
rect 8680 21916 9246 21944
rect 5350 21836 5356 21888
rect 5408 21836 5414 21888
rect 6638 21836 6644 21888
rect 6696 21836 6702 21888
rect 7742 21836 7748 21888
rect 7800 21876 7806 21888
rect 8202 21876 8208 21888
rect 7800 21848 8208 21876
rect 7800 21836 7806 21848
rect 8202 21836 8208 21848
rect 8260 21876 8266 21888
rect 8680 21876 8708 21916
rect 10410 21904 10416 21956
rect 10468 21904 10474 21956
rect 10502 21904 10508 21956
rect 10560 21944 10566 21956
rect 10796 21944 10824 21975
rect 10870 21972 10876 22024
rect 10928 21972 10934 22024
rect 11054 21972 11060 22024
rect 11112 21972 11118 22024
rect 11146 21972 11152 22024
rect 11204 21972 11210 22024
rect 11333 22015 11391 22021
rect 11333 21981 11345 22015
rect 11379 22012 11391 22015
rect 11425 22015 11483 22021
rect 11425 22012 11437 22015
rect 11379 21984 11437 22012
rect 11379 21981 11391 21984
rect 11333 21975 11391 21981
rect 11425 21981 11437 21984
rect 11471 21981 11483 22015
rect 11425 21975 11483 21981
rect 11606 21972 11612 22024
rect 11664 22012 11670 22024
rect 12066 22012 12072 22024
rect 11664 21984 12072 22012
rect 11664 21972 11670 21984
rect 12066 21972 12072 21984
rect 12124 21972 12130 22024
rect 12529 22015 12587 22021
rect 12529 21981 12541 22015
rect 12575 21981 12587 22015
rect 12529 21975 12587 21981
rect 10560 21916 10824 21944
rect 10560 21904 10566 21916
rect 8260 21848 8708 21876
rect 8941 21879 8999 21885
rect 8260 21836 8266 21848
rect 8941 21845 8953 21879
rect 8987 21876 8999 21879
rect 9490 21876 9496 21888
rect 8987 21848 9496 21876
rect 8987 21845 8999 21848
rect 8941 21839 8999 21845
rect 9490 21836 9496 21848
rect 9548 21876 9554 21888
rect 11072 21876 11100 21972
rect 12544 21944 12572 21975
rect 12618 21972 12624 22024
rect 12676 21972 12682 22024
rect 12710 21972 12716 22024
rect 12768 21972 12774 22024
rect 12986 21972 12992 22024
rect 13044 21972 13050 22024
rect 13078 21972 13084 22024
rect 13136 21972 13142 22024
rect 13280 21953 13308 22052
rect 13817 22049 13829 22052
rect 13863 22049 13875 22083
rect 17678 22080 17684 22092
rect 13817 22043 13875 22049
rect 17328 22052 17684 22080
rect 13449 22015 13507 22021
rect 13449 21981 13461 22015
rect 13495 21981 13507 22015
rect 13449 21975 13507 21981
rect 13265 21947 13323 21953
rect 13265 21944 13277 21947
rect 12544 21916 13277 21944
rect 13265 21913 13277 21916
rect 13311 21913 13323 21947
rect 13265 21907 13323 21913
rect 13354 21904 13360 21956
rect 13412 21904 13418 21956
rect 9548 21848 11100 21876
rect 9548 21836 9554 21848
rect 12710 21836 12716 21888
rect 12768 21876 12774 21888
rect 13464 21876 13492 21975
rect 13538 21972 13544 22024
rect 13596 22012 13602 22024
rect 13725 22015 13783 22021
rect 13725 22012 13737 22015
rect 13596 21984 13737 22012
rect 13596 21972 13602 21984
rect 13725 21981 13737 21984
rect 13771 21981 13783 22015
rect 13725 21975 13783 21981
rect 13909 22015 13967 22021
rect 13909 21981 13921 22015
rect 13955 22012 13967 22015
rect 13998 22012 14004 22024
rect 13955 21984 14004 22012
rect 13955 21981 13967 21984
rect 13909 21975 13967 21981
rect 13998 21972 14004 21984
rect 14056 21972 14062 22024
rect 14366 21972 14372 22024
rect 14424 21972 14430 22024
rect 14734 21972 14740 22024
rect 14792 21972 14798 22024
rect 15105 22015 15163 22021
rect 15105 21981 15117 22015
rect 15151 22012 15163 22015
rect 16574 22012 16580 22024
rect 15151 21984 16580 22012
rect 15151 21981 15163 21984
rect 15105 21975 15163 21981
rect 16574 21972 16580 21984
rect 16632 21972 16638 22024
rect 16942 21972 16948 22024
rect 17000 22012 17006 22024
rect 17037 22015 17095 22021
rect 17037 22012 17049 22015
rect 17000 21984 17049 22012
rect 17000 21972 17006 21984
rect 17037 21981 17049 21984
rect 17083 21981 17095 22015
rect 17037 21975 17095 21981
rect 17052 21944 17080 21975
rect 17126 21972 17132 22024
rect 17184 22012 17190 22024
rect 17328 22021 17356 22052
rect 17678 22040 17684 22052
rect 17736 22040 17742 22092
rect 17313 22015 17371 22021
rect 17184 21984 17229 22012
rect 17184 21972 17190 21984
rect 17313 21981 17325 22015
rect 17359 21981 17371 22015
rect 17313 21975 17371 21981
rect 17543 22015 17601 22021
rect 17543 21981 17555 22015
rect 17589 22012 17601 22015
rect 17788 22012 17816 22188
rect 18230 22176 18236 22188
rect 18288 22176 18294 22228
rect 19334 22176 19340 22228
rect 19392 22216 19398 22228
rect 19705 22219 19763 22225
rect 19705 22216 19717 22219
rect 19392 22188 19717 22216
rect 19392 22176 19398 22188
rect 19705 22185 19717 22188
rect 19751 22185 19763 22219
rect 20073 22219 20131 22225
rect 20073 22216 20085 22219
rect 19705 22179 19763 22185
rect 19904 22188 20085 22216
rect 18782 22108 18788 22160
rect 18840 22148 18846 22160
rect 19904 22148 19932 22188
rect 20073 22185 20085 22188
rect 20119 22185 20131 22219
rect 20073 22179 20131 22185
rect 20162 22176 20168 22228
rect 20220 22176 20226 22228
rect 21082 22216 21088 22228
rect 20272 22188 21088 22216
rect 18840 22120 19932 22148
rect 18840 22108 18846 22120
rect 19978 22108 19984 22160
rect 20036 22148 20042 22160
rect 20272 22148 20300 22188
rect 21082 22176 21088 22188
rect 21140 22176 21146 22228
rect 25314 22176 25320 22228
rect 25372 22176 25378 22228
rect 26053 22219 26111 22225
rect 26053 22185 26065 22219
rect 26099 22216 26111 22219
rect 26510 22216 26516 22228
rect 26099 22188 26516 22216
rect 26099 22185 26111 22188
rect 26053 22179 26111 22185
rect 26510 22176 26516 22188
rect 26568 22176 26574 22228
rect 27154 22176 27160 22228
rect 27212 22216 27218 22228
rect 27338 22216 27344 22228
rect 27212 22188 27344 22216
rect 27212 22176 27218 22188
rect 27338 22176 27344 22188
rect 27396 22176 27402 22228
rect 30006 22176 30012 22228
rect 30064 22176 30070 22228
rect 31662 22176 31668 22228
rect 31720 22216 31726 22228
rect 31941 22219 31999 22225
rect 31941 22216 31953 22219
rect 31720 22188 31953 22216
rect 31720 22176 31726 22188
rect 31941 22185 31953 22188
rect 31987 22185 31999 22219
rect 31941 22179 31999 22185
rect 33134 22176 33140 22228
rect 33192 22216 33198 22228
rect 34054 22216 34060 22228
rect 33192 22188 34060 22216
rect 33192 22176 33198 22188
rect 34054 22176 34060 22188
rect 34112 22176 34118 22228
rect 37734 22176 37740 22228
rect 37792 22216 37798 22228
rect 37918 22216 37924 22228
rect 37792 22188 37924 22216
rect 37792 22176 37798 22188
rect 37918 22176 37924 22188
rect 37976 22216 37982 22228
rect 38197 22219 38255 22225
rect 38197 22216 38209 22219
rect 37976 22188 38209 22216
rect 37976 22176 37982 22188
rect 38197 22185 38209 22188
rect 38243 22185 38255 22219
rect 38197 22179 38255 22185
rect 38289 22219 38347 22225
rect 38289 22185 38301 22219
rect 38335 22216 38347 22219
rect 38335 22188 38608 22216
rect 38335 22185 38347 22188
rect 38289 22179 38347 22185
rect 20036 22120 20300 22148
rect 20640 22120 21680 22148
rect 20036 22108 20042 22120
rect 18322 22080 18328 22092
rect 18156 22052 18328 22080
rect 17589 21984 17816 22012
rect 17957 22015 18015 22021
rect 17589 21981 17601 21984
rect 17543 21975 17601 21981
rect 17957 21981 17969 22015
rect 18003 22006 18015 22015
rect 18156 22006 18184 22052
rect 18322 22040 18328 22052
rect 18380 22080 18386 22092
rect 18598 22080 18604 22092
rect 18380 22052 18604 22080
rect 18380 22040 18386 22052
rect 18598 22040 18604 22052
rect 18656 22040 18662 22092
rect 19610 22040 19616 22092
rect 19668 22080 19674 22092
rect 20640 22080 20668 22120
rect 20993 22083 21051 22089
rect 20993 22080 21005 22083
rect 19668 22052 20668 22080
rect 20732 22052 21005 22080
rect 19668 22040 19674 22052
rect 18003 21981 18184 22006
rect 17957 21978 18184 21981
rect 17957 21975 18015 21978
rect 17052 21916 17264 21944
rect 17236 21888 17264 21916
rect 12768 21848 13492 21876
rect 13633 21879 13691 21885
rect 12768 21836 12774 21848
rect 13633 21845 13645 21879
rect 13679 21876 13691 21879
rect 13722 21876 13728 21888
rect 13679 21848 13728 21876
rect 13679 21845 13691 21848
rect 13633 21839 13691 21845
rect 13722 21836 13728 21848
rect 13780 21836 13786 21888
rect 17218 21836 17224 21888
rect 17276 21836 17282 21888
rect 17328 21876 17356 21975
rect 18230 21972 18236 22024
rect 18288 21972 18294 22024
rect 19886 21972 19892 22024
rect 19944 21972 19950 22024
rect 20254 21972 20260 22024
rect 20312 21972 20318 22024
rect 20441 22015 20499 22021
rect 20441 21981 20453 22015
rect 20487 21981 20499 22015
rect 20441 21975 20499 21981
rect 17402 21904 17408 21956
rect 17460 21904 17466 21956
rect 19904 21944 19932 21972
rect 20456 21944 20484 21975
rect 17604 21916 20484 21944
rect 20533 21947 20591 21953
rect 17604 21876 17632 21916
rect 20533 21913 20545 21947
rect 20579 21944 20591 21947
rect 20732 21944 20760 22052
rect 20993 22049 21005 22052
rect 21039 22049 21051 22083
rect 20993 22043 21051 22049
rect 21453 22083 21511 22089
rect 21453 22049 21465 22083
rect 21499 22080 21511 22083
rect 21542 22080 21548 22092
rect 21499 22052 21548 22080
rect 21499 22049 21511 22052
rect 21453 22043 21511 22049
rect 21542 22040 21548 22052
rect 21600 22040 21606 22092
rect 21652 22080 21680 22120
rect 21818 22108 21824 22160
rect 21876 22148 21882 22160
rect 22097 22151 22155 22157
rect 22097 22148 22109 22151
rect 21876 22120 22109 22148
rect 21876 22108 21882 22120
rect 22097 22117 22109 22120
rect 22143 22117 22155 22151
rect 22097 22111 22155 22117
rect 23474 22108 23480 22160
rect 23532 22148 23538 22160
rect 30024 22148 30052 22176
rect 23532 22120 30052 22148
rect 23532 22108 23538 22120
rect 32858 22108 32864 22160
rect 32916 22148 32922 22160
rect 33226 22148 33232 22160
rect 32916 22120 33232 22148
rect 32916 22108 32922 22120
rect 33226 22108 33232 22120
rect 33284 22108 33290 22160
rect 37458 22108 37464 22160
rect 37516 22148 37522 22160
rect 38381 22151 38439 22157
rect 38381 22148 38393 22151
rect 37516 22120 38393 22148
rect 37516 22108 37522 22120
rect 38381 22117 38393 22120
rect 38427 22117 38439 22151
rect 38580 22148 38608 22188
rect 38654 22176 38660 22228
rect 38712 22176 38718 22228
rect 38749 22151 38807 22157
rect 38749 22148 38761 22151
rect 38580 22120 38761 22148
rect 38381 22111 38439 22117
rect 38749 22117 38761 22120
rect 38795 22117 38807 22151
rect 38749 22111 38807 22117
rect 23753 22083 23811 22089
rect 23753 22080 23765 22083
rect 21652 22052 22094 22080
rect 22770 22066 23765 22080
rect 20809 22015 20867 22021
rect 20809 21981 20821 22015
rect 20855 22012 20867 22015
rect 20898 22012 20904 22024
rect 20855 21984 20904 22012
rect 20855 21981 20867 21984
rect 20809 21975 20867 21981
rect 20898 21972 20904 21984
rect 20956 21972 20962 22024
rect 21177 22015 21235 22021
rect 21177 21981 21189 22015
rect 21223 21981 21235 22015
rect 21177 21975 21235 21981
rect 21269 22015 21327 22021
rect 21269 21981 21281 22015
rect 21315 21981 21327 22015
rect 21269 21975 21327 21981
rect 20579 21916 20760 21944
rect 20579 21913 20591 21916
rect 20533 21907 20591 21913
rect 20990 21904 20996 21956
rect 21048 21944 21054 21956
rect 21192 21944 21220 21975
rect 21048 21916 21220 21944
rect 21284 21944 21312 21975
rect 21358 21972 21364 22024
rect 21416 21972 21422 22024
rect 21542 21944 21548 21956
rect 21284 21916 21548 21944
rect 21048 21904 21054 21916
rect 21542 21904 21548 21916
rect 21600 21904 21606 21956
rect 22066 21944 22094 22052
rect 22756 22052 23765 22066
rect 22462 21972 22468 22024
rect 22520 21972 22526 22024
rect 22756 21944 22784 22052
rect 23753 22049 23765 22052
rect 23799 22049 23811 22083
rect 23753 22043 23811 22049
rect 23842 22040 23848 22092
rect 23900 22080 23906 22092
rect 24765 22083 24823 22089
rect 24765 22080 24777 22083
rect 23900 22052 24777 22080
rect 23900 22040 23906 22052
rect 24765 22049 24777 22052
rect 24811 22049 24823 22083
rect 24765 22043 24823 22049
rect 25038 22040 25044 22092
rect 25096 22040 25102 22092
rect 25961 22083 26019 22089
rect 25332 22052 25912 22080
rect 22922 21972 22928 22024
rect 22980 21972 22986 22024
rect 23385 22015 23443 22021
rect 23385 21981 23397 22015
rect 23431 21981 23443 22015
rect 23385 21975 23443 21981
rect 22066 21916 22784 21944
rect 23400 21944 23428 21975
rect 24026 21972 24032 22024
rect 24084 21972 24090 22024
rect 24857 22015 24915 22021
rect 24857 21981 24869 22015
rect 24903 22012 24915 22015
rect 25332 22012 25360 22052
rect 25774 22012 25780 22024
rect 24903 21984 25360 22012
rect 25424 21984 25780 22012
rect 24903 21981 24915 21984
rect 24857 21975 24915 21981
rect 25038 21944 25044 21956
rect 23400 21916 25044 21944
rect 25038 21904 25044 21916
rect 25096 21904 25102 21956
rect 25133 21947 25191 21953
rect 25133 21913 25145 21947
rect 25179 21913 25191 21947
rect 25133 21907 25191 21913
rect 25338 21947 25396 21953
rect 25338 21913 25350 21947
rect 25384 21944 25396 21947
rect 25424 21944 25452 21984
rect 25774 21972 25780 21984
rect 25832 21972 25838 22024
rect 25593 21947 25651 21953
rect 25593 21944 25605 21947
rect 25384 21916 25452 21944
rect 25516 21916 25605 21944
rect 25384 21913 25396 21916
rect 25338 21907 25396 21913
rect 17328 21848 17632 21876
rect 17678 21836 17684 21888
rect 17736 21836 17742 21888
rect 17773 21879 17831 21885
rect 17773 21845 17785 21879
rect 17819 21876 17831 21879
rect 17862 21876 17868 21888
rect 17819 21848 17868 21876
rect 17819 21845 17831 21848
rect 17773 21839 17831 21845
rect 17862 21836 17868 21848
rect 17920 21836 17926 21888
rect 18141 21879 18199 21885
rect 18141 21845 18153 21879
rect 18187 21876 18199 21879
rect 19334 21876 19340 21888
rect 18187 21848 19340 21876
rect 18187 21845 18199 21848
rect 18141 21839 18199 21845
rect 19334 21836 19340 21848
rect 19392 21876 19398 21888
rect 19794 21876 19800 21888
rect 19392 21848 19800 21876
rect 19392 21836 19398 21848
rect 19794 21836 19800 21848
rect 19852 21836 19858 21888
rect 19886 21836 19892 21888
rect 19944 21876 19950 21888
rect 20631 21879 20689 21885
rect 20631 21876 20643 21879
rect 19944 21848 20643 21876
rect 19944 21836 19950 21848
rect 20631 21845 20643 21848
rect 20677 21845 20689 21879
rect 20631 21839 20689 21845
rect 20717 21879 20775 21885
rect 20717 21845 20729 21879
rect 20763 21876 20775 21879
rect 21726 21876 21732 21888
rect 20763 21848 21732 21876
rect 20763 21845 20775 21848
rect 20717 21839 20775 21845
rect 21726 21836 21732 21848
rect 21784 21836 21790 21888
rect 24394 21836 24400 21888
rect 24452 21876 24458 21888
rect 25148 21876 25176 21907
rect 25516 21885 25544 21916
rect 25593 21913 25605 21916
rect 25639 21913 25651 21947
rect 25884 21944 25912 22052
rect 25961 22049 25973 22083
rect 26007 22080 26019 22083
rect 26605 22083 26663 22089
rect 26605 22080 26617 22083
rect 26007 22052 26617 22080
rect 26007 22049 26019 22052
rect 25961 22043 26019 22049
rect 26605 22049 26617 22052
rect 26651 22049 26663 22083
rect 26605 22043 26663 22049
rect 29638 22040 29644 22092
rect 29696 22080 29702 22092
rect 30285 22083 30343 22089
rect 30285 22080 30297 22083
rect 29696 22052 30297 22080
rect 29696 22040 29702 22052
rect 30285 22049 30297 22052
rect 30331 22080 30343 22083
rect 30466 22080 30472 22092
rect 30331 22052 30472 22080
rect 30331 22049 30343 22052
rect 30285 22043 30343 22049
rect 30466 22040 30472 22052
rect 30524 22040 30530 22092
rect 32122 22040 32128 22092
rect 32180 22080 32186 22092
rect 32950 22080 32956 22092
rect 32180 22052 32956 22080
rect 32180 22040 32186 22052
rect 32950 22040 32956 22052
rect 33008 22040 33014 22092
rect 26053 22015 26111 22021
rect 26053 21981 26065 22015
rect 26099 22012 26111 22015
rect 26142 22012 26148 22024
rect 26099 21984 26148 22012
rect 26099 21981 26111 21984
rect 26053 21975 26111 21981
rect 26142 21972 26148 21984
rect 26200 21972 26206 22024
rect 26789 22015 26847 22021
rect 26789 21981 26801 22015
rect 26835 21981 26847 22015
rect 26789 21975 26847 21981
rect 26804 21944 26832 21975
rect 27062 21972 27068 22024
rect 27120 21972 27126 22024
rect 27433 22015 27491 22021
rect 27433 21981 27445 22015
rect 27479 21981 27491 22015
rect 27433 21975 27491 21981
rect 27448 21944 27476 21975
rect 27522 21972 27528 22024
rect 27580 21972 27586 22024
rect 30101 22015 30159 22021
rect 30101 21981 30113 22015
rect 30147 22012 30159 22015
rect 30190 22012 30196 22024
rect 30147 21984 30196 22012
rect 30147 21981 30159 21984
rect 30101 21975 30159 21981
rect 30190 21972 30196 21984
rect 30248 21972 30254 22024
rect 30558 21972 30564 22024
rect 30616 21972 30622 22024
rect 30745 22015 30803 22021
rect 30745 21981 30757 22015
rect 30791 22012 30803 22015
rect 32214 22012 32220 22024
rect 30791 21984 32220 22012
rect 30791 21981 30803 21984
rect 30745 21975 30803 21981
rect 32214 21972 32220 21984
rect 32272 21972 32278 22024
rect 37918 21972 37924 22024
rect 37976 21972 37982 22024
rect 38933 22015 38991 22021
rect 38933 21981 38945 22015
rect 38979 21981 38991 22015
rect 38933 21975 38991 21981
rect 27614 21944 27620 21956
rect 25884 21916 26372 21944
rect 26804 21916 27200 21944
rect 27448 21916 27620 21944
rect 25593 21907 25651 21913
rect 24452 21848 25176 21876
rect 25501 21879 25559 21885
rect 24452 21836 24458 21848
rect 25501 21845 25513 21879
rect 25547 21845 25559 21879
rect 25501 21839 25559 21845
rect 25958 21836 25964 21888
rect 26016 21876 26022 21888
rect 26142 21876 26148 21888
rect 26016 21848 26148 21876
rect 26016 21836 26022 21848
rect 26142 21836 26148 21848
rect 26200 21836 26206 21888
rect 26234 21836 26240 21888
rect 26292 21836 26298 21888
rect 26344 21876 26372 21916
rect 26970 21876 26976 21888
rect 26344 21848 26976 21876
rect 26970 21836 26976 21848
rect 27028 21836 27034 21888
rect 27172 21885 27200 21916
rect 27614 21904 27620 21916
rect 27672 21904 27678 21956
rect 31849 21947 31907 21953
rect 31849 21944 31861 21947
rect 29932 21916 31861 21944
rect 27157 21879 27215 21885
rect 27157 21845 27169 21879
rect 27203 21845 27215 21879
rect 27157 21839 27215 21845
rect 28534 21836 28540 21888
rect 28592 21876 28598 21888
rect 29932 21885 29960 21916
rect 31849 21913 31861 21916
rect 31895 21913 31907 21947
rect 31849 21907 31907 21913
rect 36538 21904 36544 21956
rect 36596 21944 36602 21956
rect 38948 21944 38976 21975
rect 39114 21972 39120 22024
rect 39172 21972 39178 22024
rect 39298 21972 39304 22024
rect 39356 21972 39362 22024
rect 39390 21972 39396 22024
rect 39448 21972 39454 22024
rect 36596 21916 38976 21944
rect 39025 21947 39083 21953
rect 36596 21904 36602 21916
rect 39025 21913 39037 21947
rect 39071 21913 39083 21947
rect 39025 21907 39083 21913
rect 29917 21879 29975 21885
rect 29917 21876 29929 21879
rect 28592 21848 29929 21876
rect 28592 21836 28598 21848
rect 29917 21845 29929 21848
rect 29963 21845 29975 21879
rect 29917 21839 29975 21845
rect 30006 21836 30012 21888
rect 30064 21876 30070 21888
rect 30377 21879 30435 21885
rect 30377 21876 30389 21879
rect 30064 21848 30389 21876
rect 30064 21836 30070 21848
rect 30377 21845 30389 21848
rect 30423 21876 30435 21879
rect 32398 21876 32404 21888
rect 30423 21848 32404 21876
rect 30423 21845 30435 21848
rect 30377 21839 30435 21845
rect 32398 21836 32404 21848
rect 32456 21836 32462 21888
rect 33962 21836 33968 21888
rect 34020 21876 34026 21888
rect 34422 21876 34428 21888
rect 34020 21848 34428 21876
rect 34020 21836 34026 21848
rect 34422 21836 34428 21848
rect 34480 21836 34486 21888
rect 37274 21836 37280 21888
rect 37332 21876 37338 21888
rect 38013 21879 38071 21885
rect 38013 21876 38025 21879
rect 37332 21848 38025 21876
rect 37332 21836 37338 21848
rect 38013 21845 38025 21848
rect 38059 21845 38071 21879
rect 38013 21839 38071 21845
rect 38102 21836 38108 21888
rect 38160 21876 38166 21888
rect 39040 21876 39068 21907
rect 38160 21848 39068 21876
rect 38160 21836 38166 21848
rect 1104 21786 40572 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 40572 21786
rect 1104 21712 40572 21734
rect 3326 21632 3332 21684
rect 3384 21672 3390 21684
rect 3973 21675 4031 21681
rect 3973 21672 3985 21675
rect 3384 21644 3985 21672
rect 3384 21632 3390 21644
rect 3973 21641 3985 21644
rect 4019 21641 4031 21675
rect 3973 21635 4031 21641
rect 4341 21675 4399 21681
rect 4341 21641 4353 21675
rect 4387 21672 4399 21675
rect 4706 21672 4712 21684
rect 4387 21644 4712 21672
rect 4387 21641 4399 21644
rect 4341 21635 4399 21641
rect 4706 21632 4712 21644
rect 4764 21632 4770 21684
rect 5169 21675 5227 21681
rect 5169 21641 5181 21675
rect 5215 21672 5227 21675
rect 5350 21672 5356 21684
rect 5215 21644 5356 21672
rect 5215 21641 5227 21644
rect 5169 21635 5227 21641
rect 5350 21632 5356 21644
rect 5408 21632 5414 21684
rect 5810 21632 5816 21684
rect 5868 21672 5874 21684
rect 6086 21672 6092 21684
rect 5868 21644 6092 21672
rect 5868 21632 5874 21644
rect 6086 21632 6092 21644
rect 6144 21632 6150 21684
rect 6181 21675 6239 21681
rect 6181 21641 6193 21675
rect 6227 21672 6239 21675
rect 6227 21644 8524 21672
rect 6227 21641 6239 21644
rect 6181 21635 6239 21641
rect 3050 21604 3056 21616
rect 2990 21576 3056 21604
rect 3050 21564 3056 21576
rect 3108 21564 3114 21616
rect 3421 21607 3479 21613
rect 3421 21573 3433 21607
rect 3467 21604 3479 21607
rect 8496 21604 8524 21644
rect 8570 21632 8576 21684
rect 8628 21632 8634 21684
rect 9769 21675 9827 21681
rect 9769 21641 9781 21675
rect 9815 21672 9827 21675
rect 10042 21672 10048 21684
rect 9815 21644 10048 21672
rect 9815 21641 9827 21644
rect 9769 21635 9827 21641
rect 10042 21632 10048 21644
rect 10100 21632 10106 21684
rect 10137 21675 10195 21681
rect 10137 21641 10149 21675
rect 10183 21672 10195 21675
rect 10410 21672 10416 21684
rect 10183 21644 10416 21672
rect 10183 21641 10195 21644
rect 10137 21635 10195 21641
rect 10410 21632 10416 21644
rect 10468 21632 10474 21684
rect 11974 21672 11980 21684
rect 11072 21644 11980 21672
rect 11072 21604 11100 21644
rect 11974 21632 11980 21644
rect 12032 21632 12038 21684
rect 13078 21632 13084 21684
rect 13136 21672 13142 21684
rect 14093 21675 14151 21681
rect 14093 21672 14105 21675
rect 13136 21644 14105 21672
rect 13136 21632 13142 21644
rect 14093 21641 14105 21644
rect 14139 21641 14151 21675
rect 14093 21635 14151 21641
rect 17126 21632 17132 21684
rect 17184 21672 17190 21684
rect 17770 21672 17776 21684
rect 17184 21644 17776 21672
rect 17184 21632 17190 21644
rect 17770 21632 17776 21644
rect 17828 21672 17834 21684
rect 20254 21672 20260 21684
rect 17828 21644 20260 21672
rect 17828 21632 17834 21644
rect 20254 21632 20260 21644
rect 20312 21632 20318 21684
rect 20346 21632 20352 21684
rect 20404 21672 20410 21684
rect 20809 21675 20867 21681
rect 20809 21672 20821 21675
rect 20404 21644 20821 21672
rect 20404 21632 20410 21644
rect 20809 21641 20821 21644
rect 20855 21641 20867 21675
rect 21358 21672 21364 21684
rect 20809 21635 20867 21641
rect 21100 21644 21364 21672
rect 3467 21576 6040 21604
rect 8496 21576 11100 21604
rect 3467 21573 3479 21576
rect 3421 21567 3479 21573
rect 3602 21496 3608 21548
rect 3660 21496 3666 21548
rect 3694 21496 3700 21548
rect 3752 21536 3758 21548
rect 3789 21539 3847 21545
rect 3789 21536 3801 21539
rect 3752 21508 3801 21536
rect 3752 21496 3758 21508
rect 3789 21505 3801 21508
rect 3835 21505 3847 21539
rect 3789 21499 3847 21505
rect 3878 21496 3884 21548
rect 3936 21496 3942 21548
rect 4430 21496 4436 21548
rect 4488 21496 4494 21548
rect 5718 21496 5724 21548
rect 5776 21496 5782 21548
rect 5902 21496 5908 21548
rect 5960 21496 5966 21548
rect 6012 21545 6040 21576
rect 11146 21564 11152 21616
rect 11204 21604 11210 21616
rect 11204 21576 12572 21604
rect 11204 21564 11210 21576
rect 5997 21539 6055 21545
rect 5997 21505 6009 21539
rect 6043 21505 6055 21539
rect 5997 21499 6055 21505
rect 8202 21496 8208 21548
rect 8260 21496 8266 21548
rect 8570 21496 8576 21548
rect 8628 21536 8634 21548
rect 9217 21539 9275 21545
rect 9217 21536 9229 21539
rect 8628 21508 9229 21536
rect 8628 21496 8634 21508
rect 9217 21505 9229 21508
rect 9263 21505 9275 21539
rect 10502 21536 10508 21548
rect 9217 21499 9275 21505
rect 9600 21508 10508 21536
rect 1486 21428 1492 21480
rect 1544 21428 1550 21480
rect 1765 21471 1823 21477
rect 1765 21437 1777 21471
rect 1811 21468 1823 21471
rect 4617 21471 4675 21477
rect 1811 21440 3832 21468
rect 1811 21437 1823 21440
rect 1765 21431 1823 21437
rect 3804 21400 3832 21440
rect 4617 21437 4629 21471
rect 4663 21468 4675 21471
rect 4663 21440 5120 21468
rect 4663 21437 4675 21440
rect 4617 21431 4675 21437
rect 5092 21412 5120 21440
rect 5166 21428 5172 21480
rect 5224 21468 5230 21480
rect 5261 21471 5319 21477
rect 5261 21468 5273 21471
rect 5224 21440 5273 21468
rect 5224 21428 5230 21440
rect 5261 21437 5273 21440
rect 5307 21437 5319 21471
rect 5261 21431 5319 21437
rect 5353 21471 5411 21477
rect 5353 21437 5365 21471
rect 5399 21437 5411 21471
rect 5353 21431 5411 21437
rect 4801 21403 4859 21409
rect 4801 21400 4813 21403
rect 3804 21372 4813 21400
rect 4801 21369 4813 21372
rect 4847 21369 4859 21403
rect 4801 21363 4859 21369
rect 5074 21360 5080 21412
rect 5132 21400 5138 21412
rect 5368 21400 5396 21431
rect 5442 21428 5448 21480
rect 5500 21468 5506 21480
rect 6822 21468 6828 21480
rect 5500 21440 6828 21468
rect 5500 21428 5506 21440
rect 6822 21428 6828 21440
rect 6880 21428 6886 21480
rect 7101 21471 7159 21477
rect 7101 21437 7113 21471
rect 7147 21468 7159 21471
rect 7650 21468 7656 21480
rect 7147 21440 7656 21468
rect 7147 21437 7159 21440
rect 7101 21431 7159 21437
rect 7650 21428 7656 21440
rect 7708 21428 7714 21480
rect 8386 21428 8392 21480
rect 8444 21468 8450 21480
rect 9600 21477 9628 21508
rect 10502 21496 10508 21508
rect 10560 21496 10566 21548
rect 9585 21471 9643 21477
rect 9585 21468 9597 21471
rect 8444 21440 9597 21468
rect 8444 21428 8450 21440
rect 9585 21437 9597 21440
rect 9631 21437 9643 21471
rect 9585 21431 9643 21437
rect 9677 21471 9735 21477
rect 9677 21437 9689 21471
rect 9723 21468 9735 21471
rect 9858 21468 9864 21480
rect 9723 21440 9864 21468
rect 9723 21437 9735 21440
rect 9677 21431 9735 21437
rect 9858 21428 9864 21440
rect 9916 21428 9922 21480
rect 5132 21372 5396 21400
rect 5132 21360 5138 21372
rect 5810 21360 5816 21412
rect 5868 21360 5874 21412
rect 11422 21400 11428 21412
rect 8128 21372 11428 21400
rect 3237 21335 3295 21341
rect 3237 21301 3249 21335
rect 3283 21332 3295 21335
rect 5626 21332 5632 21344
rect 3283 21304 5632 21332
rect 3283 21301 3295 21304
rect 3237 21295 3295 21301
rect 5626 21292 5632 21304
rect 5684 21292 5690 21344
rect 6638 21292 6644 21344
rect 6696 21332 6702 21344
rect 8128 21332 8156 21372
rect 11422 21360 11428 21372
rect 11480 21360 11486 21412
rect 6696 21304 8156 21332
rect 6696 21292 6702 21304
rect 8662 21292 8668 21344
rect 8720 21292 8726 21344
rect 12544 21332 12572 21576
rect 12618 21564 12624 21616
rect 12676 21604 12682 21616
rect 13173 21607 13231 21613
rect 12676 21576 13124 21604
rect 12676 21564 12682 21576
rect 12800 21539 12858 21545
rect 12800 21505 12812 21539
rect 12846 21505 12858 21539
rect 12800 21499 12858 21505
rect 12820 21468 12848 21499
rect 12894 21496 12900 21548
rect 12952 21496 12958 21548
rect 12986 21496 12992 21548
rect 13044 21496 13050 21548
rect 13096 21536 13124 21576
rect 13173 21573 13185 21607
rect 13219 21604 13231 21607
rect 13906 21604 13912 21616
rect 13219 21576 13912 21604
rect 13219 21573 13231 21576
rect 13173 21567 13231 21573
rect 13906 21564 13912 21576
rect 13964 21564 13970 21616
rect 16761 21607 16819 21613
rect 16761 21604 16773 21607
rect 14752 21576 16773 21604
rect 14752 21548 14780 21576
rect 16761 21573 16773 21576
rect 16807 21604 16819 21607
rect 20622 21604 20628 21616
rect 16807 21576 16988 21604
rect 16807 21573 16819 21576
rect 16761 21567 16819 21573
rect 13354 21536 13360 21548
rect 13096 21508 13360 21536
rect 13354 21496 13360 21508
rect 13412 21496 13418 21548
rect 14277 21539 14335 21545
rect 14277 21505 14289 21539
rect 14323 21536 14335 21539
rect 14366 21536 14372 21548
rect 14323 21508 14372 21536
rect 14323 21505 14335 21508
rect 14277 21499 14335 21505
rect 14366 21496 14372 21508
rect 14424 21496 14430 21548
rect 14461 21539 14519 21545
rect 14461 21505 14473 21539
rect 14507 21536 14519 21539
rect 14734 21536 14740 21548
rect 14507 21508 14740 21536
rect 14507 21505 14519 21508
rect 14461 21499 14519 21505
rect 14734 21496 14740 21508
rect 14792 21496 14798 21548
rect 16960 21545 16988 21576
rect 17144 21576 20628 21604
rect 17144 21545 17172 21576
rect 20622 21564 20628 21576
rect 20680 21564 20686 21616
rect 21100 21613 21128 21644
rect 21358 21632 21364 21644
rect 21416 21672 21422 21684
rect 22186 21672 22192 21684
rect 21416 21644 22192 21672
rect 21416 21632 21422 21644
rect 22186 21632 22192 21644
rect 22244 21632 22250 21684
rect 23851 21675 23909 21681
rect 23851 21641 23863 21675
rect 23897 21672 23909 21675
rect 24394 21672 24400 21684
rect 23897 21644 24400 21672
rect 23897 21641 23909 21644
rect 23851 21635 23909 21641
rect 24394 21632 24400 21644
rect 24452 21632 24458 21684
rect 25038 21632 25044 21684
rect 25096 21672 25102 21684
rect 25774 21672 25780 21684
rect 25096 21644 25780 21672
rect 25096 21632 25102 21644
rect 25774 21632 25780 21644
rect 25832 21632 25838 21684
rect 26694 21632 26700 21684
rect 26752 21672 26758 21684
rect 26752 21644 27660 21672
rect 26752 21632 26758 21644
rect 21085 21607 21143 21613
rect 21085 21573 21097 21607
rect 21131 21573 21143 21607
rect 21085 21567 21143 21573
rect 23382 21564 23388 21616
rect 23440 21604 23446 21616
rect 23937 21607 23995 21613
rect 23937 21604 23949 21607
rect 23440 21576 23949 21604
rect 23440 21564 23446 21576
rect 23937 21573 23949 21576
rect 23983 21604 23995 21607
rect 25590 21604 25596 21616
rect 23983 21576 25596 21604
rect 23983 21573 23995 21576
rect 23937 21567 23995 21573
rect 25590 21564 25596 21576
rect 25648 21564 25654 21616
rect 27062 21564 27068 21616
rect 27120 21604 27126 21616
rect 27632 21613 27660 21644
rect 33226 21632 33232 21684
rect 33284 21672 33290 21684
rect 33689 21675 33747 21681
rect 33689 21672 33701 21675
rect 33284 21644 33701 21672
rect 33284 21632 33290 21644
rect 33689 21641 33701 21644
rect 33735 21672 33747 21675
rect 33778 21672 33784 21684
rect 33735 21644 33784 21672
rect 33735 21641 33747 21644
rect 33689 21635 33747 21641
rect 33778 21632 33784 21644
rect 33836 21632 33842 21684
rect 34057 21675 34115 21681
rect 34057 21641 34069 21675
rect 34103 21641 34115 21675
rect 34057 21635 34115 21641
rect 27525 21607 27583 21613
rect 27525 21604 27537 21607
rect 27120 21576 27537 21604
rect 27120 21564 27126 21576
rect 27525 21573 27537 21576
rect 27571 21573 27583 21607
rect 27525 21567 27583 21573
rect 27617 21607 27675 21613
rect 27617 21573 27629 21607
rect 27663 21604 27675 21607
rect 27890 21604 27896 21616
rect 27663 21576 27896 21604
rect 27663 21573 27675 21576
rect 27617 21567 27675 21573
rect 27890 21564 27896 21576
rect 27948 21564 27954 21616
rect 28077 21607 28135 21613
rect 28077 21573 28089 21607
rect 28123 21604 28135 21607
rect 28994 21604 29000 21616
rect 28123 21576 29000 21604
rect 28123 21573 28135 21576
rect 28077 21567 28135 21573
rect 28994 21564 29000 21576
rect 29052 21564 29058 21616
rect 31478 21564 31484 21616
rect 31536 21604 31542 21616
rect 34072 21604 34100 21635
rect 34146 21632 34152 21684
rect 34204 21672 34210 21684
rect 34606 21672 34612 21684
rect 34204 21644 34612 21672
rect 34204 21632 34210 21644
rect 34606 21632 34612 21644
rect 34664 21672 34670 21684
rect 34664 21644 34744 21672
rect 34664 21632 34670 21644
rect 34716 21613 34744 21644
rect 34790 21632 34796 21684
rect 34848 21672 34854 21684
rect 34848 21644 35848 21672
rect 34848 21632 34854 21644
rect 31536 21576 34100 21604
rect 34701 21607 34759 21613
rect 31536 21564 31542 21576
rect 16669 21539 16727 21545
rect 16669 21505 16681 21539
rect 16715 21536 16727 21539
rect 16853 21539 16911 21545
rect 16715 21508 16804 21536
rect 16715 21505 16727 21508
rect 16669 21499 16727 21505
rect 13262 21468 13268 21480
rect 12820 21440 13268 21468
rect 13262 21428 13268 21440
rect 13320 21428 13326 21480
rect 12710 21360 12716 21412
rect 12768 21400 12774 21412
rect 13173 21403 13231 21409
rect 13173 21400 13185 21403
rect 12768 21372 13185 21400
rect 12768 21360 12774 21372
rect 13173 21369 13185 21372
rect 13219 21369 13231 21403
rect 14384 21400 14412 21496
rect 14553 21471 14611 21477
rect 14553 21437 14565 21471
rect 14599 21468 14611 21471
rect 16574 21468 16580 21480
rect 14599 21440 16580 21468
rect 14599 21437 14611 21440
rect 14553 21431 14611 21437
rect 16574 21428 16580 21440
rect 16632 21428 16638 21480
rect 15102 21400 15108 21412
rect 14384 21372 15108 21400
rect 13173 21363 13231 21369
rect 15102 21360 15108 21372
rect 15160 21360 15166 21412
rect 16776 21400 16804 21508
rect 16853 21505 16865 21539
rect 16899 21505 16911 21539
rect 16853 21499 16911 21505
rect 16945 21539 17003 21545
rect 16945 21505 16957 21539
rect 16991 21505 17003 21539
rect 16945 21499 17003 21505
rect 17129 21539 17187 21545
rect 17129 21505 17141 21539
rect 17175 21505 17187 21539
rect 17129 21499 17187 21505
rect 16868 21468 16896 21499
rect 17862 21496 17868 21548
rect 17920 21536 17926 21548
rect 18782 21536 18788 21548
rect 17920 21508 18788 21536
rect 17920 21496 17926 21508
rect 18782 21496 18788 21508
rect 18840 21496 18846 21548
rect 20806 21496 20812 21548
rect 20864 21536 20870 21548
rect 20947 21539 21005 21545
rect 20947 21536 20959 21539
rect 20864 21508 20959 21536
rect 20864 21496 20870 21508
rect 20947 21505 20959 21508
rect 20993 21505 21005 21539
rect 21177 21539 21235 21545
rect 21177 21536 21189 21539
rect 20947 21499 21005 21505
rect 21100 21508 21189 21536
rect 17034 21468 17040 21480
rect 16868 21440 17040 21468
rect 17034 21428 17040 21440
rect 17092 21468 17098 21480
rect 18230 21468 18236 21480
rect 17092 21440 18236 21468
rect 17092 21428 17098 21440
rect 18230 21428 18236 21440
rect 18288 21468 18294 21480
rect 19426 21468 19432 21480
rect 18288 21440 19432 21468
rect 18288 21428 18294 21440
rect 19426 21428 19432 21440
rect 19484 21468 19490 21480
rect 21100 21468 21128 21508
rect 21177 21505 21189 21508
rect 21223 21505 21235 21539
rect 21177 21499 21235 21505
rect 21360 21539 21418 21545
rect 21360 21505 21372 21539
rect 21406 21505 21418 21539
rect 21360 21499 21418 21505
rect 21453 21539 21511 21545
rect 21453 21505 21465 21539
rect 21499 21536 21511 21539
rect 21818 21536 21824 21548
rect 21499 21508 21824 21536
rect 21499 21505 21511 21508
rect 21453 21499 21511 21505
rect 19484 21440 21128 21468
rect 19484 21428 19490 21440
rect 17402 21400 17408 21412
rect 16776 21372 17408 21400
rect 17402 21360 17408 21372
rect 17460 21360 17466 21412
rect 20254 21360 20260 21412
rect 20312 21400 20318 21412
rect 21376 21400 21404 21499
rect 21818 21496 21824 21508
rect 21876 21496 21882 21548
rect 23750 21496 23756 21548
rect 23808 21496 23814 21548
rect 24029 21539 24087 21545
rect 24029 21505 24041 21539
rect 24075 21536 24087 21539
rect 24118 21536 24124 21548
rect 24075 21508 24124 21536
rect 24075 21505 24087 21508
rect 24029 21499 24087 21505
rect 24118 21496 24124 21508
rect 24176 21496 24182 21548
rect 24394 21496 24400 21548
rect 24452 21536 24458 21548
rect 24578 21536 24584 21548
rect 24452 21508 24584 21536
rect 24452 21496 24458 21508
rect 24578 21496 24584 21508
rect 24636 21496 24642 21548
rect 24854 21496 24860 21548
rect 24912 21536 24918 21548
rect 25682 21536 25688 21548
rect 24912 21508 25688 21536
rect 24912 21496 24918 21508
rect 25682 21496 25688 21508
rect 25740 21496 25746 21548
rect 27246 21496 27252 21548
rect 27304 21496 27310 21548
rect 27338 21496 27344 21548
rect 27396 21536 27402 21548
rect 27396 21508 27441 21536
rect 27396 21496 27402 21508
rect 27706 21496 27712 21548
rect 27764 21545 27770 21548
rect 27764 21536 27772 21545
rect 27764 21508 27809 21536
rect 27764 21499 27772 21508
rect 27764 21496 27770 21499
rect 27982 21496 27988 21548
rect 28040 21496 28046 21548
rect 28261 21539 28319 21545
rect 28261 21505 28273 21539
rect 28307 21536 28319 21539
rect 29086 21536 29092 21548
rect 28307 21508 29092 21536
rect 28307 21505 28319 21508
rect 28261 21499 28319 21505
rect 29086 21496 29092 21508
rect 29144 21496 29150 21548
rect 31846 21496 31852 21548
rect 31904 21536 31910 21548
rect 33042 21536 33048 21548
rect 31904 21508 33048 21536
rect 31904 21496 31910 21508
rect 33042 21496 33048 21508
rect 33100 21496 33106 21548
rect 33520 21545 33548 21576
rect 34701 21573 34713 21607
rect 34747 21573 34759 21607
rect 34701 21567 34759 21573
rect 35250 21564 35256 21616
rect 35308 21604 35314 21616
rect 35820 21613 35848 21644
rect 35575 21607 35633 21613
rect 35575 21604 35587 21607
rect 35308 21576 35587 21604
rect 35308 21564 35314 21576
rect 35575 21573 35587 21576
rect 35621 21573 35633 21607
rect 35575 21567 35633 21573
rect 35805 21607 35863 21613
rect 35805 21573 35817 21607
rect 35851 21573 35863 21607
rect 35805 21567 35863 21573
rect 36262 21564 36268 21616
rect 36320 21604 36326 21616
rect 36357 21607 36415 21613
rect 36357 21604 36369 21607
rect 36320 21576 36369 21604
rect 36320 21564 36326 21576
rect 36357 21573 36369 21576
rect 36403 21573 36415 21607
rect 36357 21567 36415 21573
rect 33505 21539 33563 21545
rect 33505 21505 33517 21539
rect 33551 21505 33563 21539
rect 33505 21499 33563 21505
rect 33873 21539 33931 21545
rect 33873 21505 33885 21539
rect 33919 21505 33931 21539
rect 33873 21499 33931 21505
rect 34517 21539 34575 21545
rect 34517 21505 34529 21539
rect 34563 21536 34575 21539
rect 34606 21536 34612 21548
rect 34563 21508 34612 21536
rect 34563 21505 34575 21508
rect 34517 21499 34575 21505
rect 22094 21400 22100 21412
rect 20312 21372 22100 21400
rect 20312 21360 20318 21372
rect 22094 21360 22100 21372
rect 22152 21360 22158 21412
rect 22186 21360 22192 21412
rect 22244 21400 22250 21412
rect 24118 21400 24124 21412
rect 22244 21372 24124 21400
rect 22244 21360 22250 21372
rect 24118 21360 24124 21372
rect 24176 21400 24182 21412
rect 27356 21400 27384 21496
rect 28353 21471 28411 21477
rect 28353 21468 28365 21471
rect 24176 21372 27384 21400
rect 27448 21440 28365 21468
rect 24176 21360 24182 21372
rect 12986 21332 12992 21344
rect 12544 21304 12992 21332
rect 12986 21292 12992 21304
rect 13044 21292 13050 21344
rect 14734 21292 14740 21344
rect 14792 21332 14798 21344
rect 15010 21332 15016 21344
rect 14792 21304 15016 21332
rect 14792 21292 14798 21304
rect 15010 21292 15016 21304
rect 15068 21292 15074 21344
rect 17037 21335 17095 21341
rect 17037 21301 17049 21335
rect 17083 21332 17095 21335
rect 17310 21332 17316 21344
rect 17083 21304 17316 21332
rect 17083 21301 17095 21304
rect 17037 21295 17095 21301
rect 17310 21292 17316 21304
rect 17368 21292 17374 21344
rect 20622 21292 20628 21344
rect 20680 21332 20686 21344
rect 21542 21332 21548 21344
rect 20680 21304 21548 21332
rect 20680 21292 20686 21304
rect 21542 21292 21548 21304
rect 21600 21332 21606 21344
rect 26602 21332 26608 21344
rect 21600 21304 26608 21332
rect 21600 21292 21606 21304
rect 26602 21292 26608 21304
rect 26660 21332 26666 21344
rect 27448 21332 27476 21440
rect 28353 21437 28365 21440
rect 28399 21437 28411 21471
rect 28353 21431 28411 21437
rect 32766 21360 32772 21412
rect 32824 21400 32830 21412
rect 33888 21400 33916 21499
rect 34606 21496 34612 21508
rect 34664 21496 34670 21548
rect 34793 21539 34851 21545
rect 34793 21505 34805 21539
rect 34839 21505 34851 21539
rect 34793 21499 34851 21505
rect 33962 21428 33968 21480
rect 34020 21468 34026 21480
rect 34808 21468 34836 21499
rect 34882 21496 34888 21548
rect 34940 21496 34946 21548
rect 35437 21539 35495 21545
rect 35437 21536 35449 21539
rect 34992 21508 35449 21536
rect 34992 21468 35020 21508
rect 35437 21505 35449 21508
rect 35483 21505 35495 21539
rect 35437 21499 35495 21505
rect 35710 21496 35716 21548
rect 35768 21496 35774 21548
rect 35894 21496 35900 21548
rect 35952 21496 35958 21548
rect 35986 21496 35992 21548
rect 36044 21536 36050 21548
rect 36173 21539 36231 21545
rect 36173 21536 36185 21539
rect 36044 21508 36185 21536
rect 36044 21496 36050 21508
rect 36173 21505 36185 21508
rect 36219 21505 36231 21539
rect 36173 21499 36231 21505
rect 34020 21440 34836 21468
rect 34900 21440 35020 21468
rect 36188 21468 36216 21499
rect 36446 21496 36452 21548
rect 36504 21496 36510 21548
rect 36538 21496 36544 21548
rect 36596 21496 36602 21548
rect 38930 21468 38936 21480
rect 36188 21440 38936 21468
rect 34020 21428 34026 21440
rect 32824 21372 33916 21400
rect 32824 21360 32830 21372
rect 34422 21360 34428 21412
rect 34480 21400 34486 21412
rect 34900 21400 34928 21440
rect 38930 21428 38936 21440
rect 38988 21428 38994 21480
rect 34480 21372 34928 21400
rect 34480 21360 34486 21372
rect 26660 21304 27476 21332
rect 27893 21335 27951 21341
rect 26660 21292 26666 21304
rect 27893 21301 27905 21335
rect 27939 21332 27951 21335
rect 27982 21332 27988 21344
rect 27939 21304 27988 21332
rect 27939 21301 27951 21304
rect 27893 21295 27951 21301
rect 27982 21292 27988 21304
rect 28040 21292 28046 21344
rect 28350 21292 28356 21344
rect 28408 21292 28414 21344
rect 29730 21292 29736 21344
rect 29788 21332 29794 21344
rect 30190 21332 30196 21344
rect 29788 21304 30196 21332
rect 29788 21292 29794 21304
rect 30190 21292 30196 21304
rect 30248 21292 30254 21344
rect 30926 21292 30932 21344
rect 30984 21332 30990 21344
rect 31294 21332 31300 21344
rect 30984 21304 31300 21332
rect 30984 21292 30990 21304
rect 31294 21292 31300 21304
rect 31352 21292 31358 21344
rect 31662 21292 31668 21344
rect 31720 21292 31726 21344
rect 32214 21292 32220 21344
rect 32272 21332 32278 21344
rect 33226 21332 33232 21344
rect 32272 21304 33232 21332
rect 32272 21292 32278 21304
rect 33226 21292 33232 21304
rect 33284 21292 33290 21344
rect 35069 21335 35127 21341
rect 35069 21301 35081 21335
rect 35115 21332 35127 21335
rect 35986 21332 35992 21344
rect 35115 21304 35992 21332
rect 35115 21301 35127 21304
rect 35069 21295 35127 21301
rect 35986 21292 35992 21304
rect 36044 21292 36050 21344
rect 36081 21335 36139 21341
rect 36081 21301 36093 21335
rect 36127 21332 36139 21335
rect 36170 21332 36176 21344
rect 36127 21304 36176 21332
rect 36127 21301 36139 21304
rect 36081 21295 36139 21301
rect 36170 21292 36176 21304
rect 36228 21292 36234 21344
rect 36725 21335 36783 21341
rect 36725 21301 36737 21335
rect 36771 21332 36783 21335
rect 37274 21332 37280 21344
rect 36771 21304 37280 21332
rect 36771 21301 36783 21304
rect 36725 21295 36783 21301
rect 37274 21292 37280 21304
rect 37332 21292 37338 21344
rect 1104 21242 40572 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 40572 21242
rect 1104 21168 40572 21190
rect 6270 21088 6276 21140
rect 6328 21128 6334 21140
rect 6641 21131 6699 21137
rect 6641 21128 6653 21131
rect 6328 21100 6653 21128
rect 6328 21088 6334 21100
rect 6641 21097 6653 21100
rect 6687 21097 6699 21131
rect 6641 21091 6699 21097
rect 6730 21088 6736 21140
rect 6788 21128 6794 21140
rect 6788 21100 7144 21128
rect 6788 21088 6794 21100
rect 6178 21020 6184 21072
rect 6236 21060 6242 21072
rect 6549 21063 6607 21069
rect 6236 21032 6316 21060
rect 6236 21020 6242 21032
rect 2866 20952 2872 21004
rect 2924 20992 2930 21004
rect 3326 20992 3332 21004
rect 2924 20964 3332 20992
rect 2924 20952 2930 20964
rect 3326 20952 3332 20964
rect 3384 20992 3390 21004
rect 5074 20992 5080 21004
rect 3384 20964 5080 20992
rect 3384 20952 3390 20964
rect 5074 20952 5080 20964
rect 5132 20952 5138 21004
rect 1578 20884 1584 20936
rect 1636 20924 1642 20936
rect 1857 20927 1915 20933
rect 1857 20924 1869 20927
rect 1636 20896 1869 20924
rect 1636 20884 1642 20896
rect 1857 20893 1869 20896
rect 1903 20893 1915 20927
rect 1857 20887 1915 20893
rect 4890 20884 4896 20936
rect 4948 20924 4954 20936
rect 5442 20924 5448 20936
rect 4948 20896 5448 20924
rect 4948 20884 4954 20896
rect 5442 20884 5448 20896
rect 5500 20884 5506 20936
rect 5905 20927 5963 20933
rect 5905 20893 5917 20927
rect 5951 20893 5963 20927
rect 5905 20887 5963 20893
rect 2130 20816 2136 20868
rect 2188 20816 2194 20868
rect 3786 20856 3792 20868
rect 3358 20828 3792 20856
rect 3786 20816 3792 20828
rect 3844 20816 3850 20868
rect 4801 20859 4859 20865
rect 4801 20825 4813 20859
rect 4847 20856 4859 20859
rect 5261 20859 5319 20865
rect 5261 20856 5273 20859
rect 4847 20828 5273 20856
rect 4847 20825 4859 20828
rect 4801 20819 4859 20825
rect 5261 20825 5273 20828
rect 5307 20825 5319 20859
rect 5261 20819 5319 20825
rect 5350 20816 5356 20868
rect 5408 20856 5414 20868
rect 5920 20856 5948 20887
rect 5994 20884 6000 20936
rect 6052 20884 6058 20936
rect 6089 20927 6147 20933
rect 6089 20893 6101 20927
rect 6135 20893 6147 20927
rect 6089 20887 6147 20893
rect 6104 20856 6132 20887
rect 6178 20884 6184 20936
rect 6236 20933 6242 20936
rect 6288 20934 6316 21032
rect 6549 21029 6561 21063
rect 6595 21060 6607 21063
rect 7006 21060 7012 21072
rect 6595 21032 7012 21060
rect 6595 21029 6607 21032
rect 6549 21023 6607 21029
rect 7006 21020 7012 21032
rect 7064 21020 7070 21072
rect 7116 21060 7144 21100
rect 7650 21088 7656 21140
rect 7708 21088 7714 21140
rect 10226 21088 10232 21140
rect 10284 21128 10290 21140
rect 10502 21128 10508 21140
rect 10284 21100 10508 21128
rect 10284 21088 10290 21100
rect 10502 21088 10508 21100
rect 10560 21088 10566 21140
rect 10870 21088 10876 21140
rect 10928 21088 10934 21140
rect 13262 21128 13268 21140
rect 10980 21100 13268 21128
rect 8478 21060 8484 21072
rect 7116 21032 8484 21060
rect 6288 20933 6408 20934
rect 6236 20927 6258 20933
rect 6246 20893 6258 20927
rect 6288 20927 6423 20933
rect 6288 20906 6377 20927
rect 6236 20887 6258 20893
rect 6365 20893 6377 20906
rect 6411 20893 6423 20927
rect 6730 20924 6736 20936
rect 6365 20887 6423 20893
rect 6564 20896 6736 20924
rect 6236 20884 6242 20887
rect 6564 20856 6592 20896
rect 6730 20884 6736 20896
rect 6788 20884 6794 20936
rect 6825 20927 6883 20933
rect 6825 20893 6837 20927
rect 6871 20924 6883 20927
rect 7116 20924 7144 21032
rect 8478 21020 8484 21032
rect 8536 21060 8542 21072
rect 10980 21060 11008 21100
rect 13262 21088 13268 21100
rect 13320 21088 13326 21140
rect 15470 21088 15476 21140
rect 15528 21128 15534 21140
rect 23385 21131 23443 21137
rect 23385 21128 23397 21131
rect 15528 21100 23397 21128
rect 15528 21088 15534 21100
rect 23385 21097 23397 21100
rect 23431 21097 23443 21131
rect 23385 21091 23443 21097
rect 23569 21131 23627 21137
rect 23569 21097 23581 21131
rect 23615 21097 23627 21131
rect 23569 21091 23627 21097
rect 8536 21032 11008 21060
rect 8536 21020 8542 21032
rect 7466 20952 7472 21004
rect 7524 20992 7530 21004
rect 8297 20995 8355 21001
rect 8297 20992 8309 20995
rect 7524 20964 8309 20992
rect 7524 20952 7530 20964
rect 8297 20961 8309 20964
rect 8343 20992 8355 20995
rect 9858 20992 9864 21004
rect 8343 20964 9864 20992
rect 8343 20961 8355 20964
rect 8297 20955 8355 20961
rect 9858 20952 9864 20964
rect 9916 20952 9922 21004
rect 10134 20952 10140 21004
rect 10192 20992 10198 21004
rect 10192 20964 10365 20992
rect 10192 20952 10198 20964
rect 6871 20896 7144 20924
rect 6871 20893 6883 20896
rect 6825 20887 6883 20893
rect 7190 20884 7196 20936
rect 7248 20884 7254 20936
rect 8021 20927 8079 20933
rect 8021 20893 8033 20927
rect 8067 20924 8079 20927
rect 8662 20924 8668 20936
rect 8067 20896 8668 20924
rect 8067 20893 8079 20896
rect 8021 20887 8079 20893
rect 8662 20884 8668 20896
rect 8720 20884 8726 20936
rect 10226 20884 10232 20936
rect 10284 20884 10290 20936
rect 10337 20933 10365 20964
rect 10322 20927 10380 20933
rect 10322 20893 10334 20927
rect 10368 20893 10380 20927
rect 10322 20887 10380 20893
rect 10694 20927 10752 20933
rect 10694 20893 10706 20927
rect 10740 20924 10752 20927
rect 10796 20924 10824 21032
rect 17126 21020 17132 21072
rect 17184 21060 17190 21072
rect 17313 21063 17371 21069
rect 17313 21060 17325 21063
rect 17184 21032 17325 21060
rect 17184 21020 17190 21032
rect 17313 21029 17325 21032
rect 17359 21029 17371 21063
rect 17313 21023 17371 21029
rect 18414 21020 18420 21072
rect 18472 21060 18478 21072
rect 18693 21063 18751 21069
rect 18693 21060 18705 21063
rect 18472 21032 18705 21060
rect 18472 21020 18478 21032
rect 18693 21029 18705 21032
rect 18739 21029 18751 21063
rect 18693 21023 18751 21029
rect 20806 21020 20812 21072
rect 20864 21060 20870 21072
rect 21910 21060 21916 21072
rect 20864 21032 21916 21060
rect 20864 21020 20870 21032
rect 21910 21020 21916 21032
rect 21968 21020 21974 21072
rect 23198 21020 23204 21072
rect 23256 21060 23262 21072
rect 23584 21060 23612 21091
rect 28994 21088 29000 21140
rect 29052 21128 29058 21140
rect 36446 21128 36452 21140
rect 29052 21100 36452 21128
rect 29052 21088 29058 21100
rect 36446 21088 36452 21100
rect 36504 21088 36510 21140
rect 36541 21131 36599 21137
rect 36541 21097 36553 21131
rect 36587 21097 36599 21131
rect 36541 21091 36599 21097
rect 25038 21060 25044 21072
rect 23256 21032 23612 21060
rect 23676 21032 25044 21060
rect 23256 21020 23262 21032
rect 10965 20995 11023 21001
rect 10965 20961 10977 20995
rect 11011 20992 11023 20995
rect 11238 20992 11244 21004
rect 11011 20964 11244 20992
rect 11011 20961 11023 20964
rect 10965 20955 11023 20961
rect 11238 20952 11244 20964
rect 11296 20952 11302 21004
rect 12713 20995 12771 21001
rect 12713 20961 12725 20995
rect 12759 20992 12771 20995
rect 12894 20992 12900 21004
rect 12759 20964 12900 20992
rect 12759 20961 12771 20964
rect 12713 20955 12771 20961
rect 12894 20952 12900 20964
rect 12952 20992 12958 21004
rect 13357 20995 13415 21001
rect 13357 20992 13369 20995
rect 12952 20964 13369 20992
rect 12952 20952 12958 20964
rect 13357 20961 13369 20964
rect 13403 20961 13415 20995
rect 15470 20992 15476 21004
rect 13357 20955 13415 20961
rect 14752 20964 15476 20992
rect 10740 20896 10824 20924
rect 13725 20927 13783 20933
rect 10740 20893 10752 20896
rect 10694 20887 10752 20893
rect 13725 20893 13737 20927
rect 13771 20893 13783 20927
rect 13725 20887 13783 20893
rect 5408 20828 6040 20856
rect 6104 20828 6592 20856
rect 6917 20859 6975 20865
rect 5408 20816 5414 20828
rect 3602 20748 3608 20800
rect 3660 20748 3666 20800
rect 4430 20748 4436 20800
rect 4488 20748 4494 20800
rect 6012 20788 6040 20828
rect 6917 20825 6929 20859
rect 6963 20825 6975 20859
rect 6917 20819 6975 20825
rect 6932 20788 6960 20819
rect 7006 20816 7012 20868
rect 7064 20856 7070 20868
rect 7064 20828 8340 20856
rect 7064 20816 7070 20828
rect 8312 20800 8340 20828
rect 8570 20816 8576 20868
rect 8628 20856 8634 20868
rect 10505 20859 10563 20865
rect 10505 20856 10517 20859
rect 8628 20828 10517 20856
rect 8628 20816 8634 20828
rect 10505 20825 10517 20828
rect 10551 20825 10563 20859
rect 10505 20819 10563 20825
rect 6012 20760 6960 20788
rect 8113 20791 8171 20797
rect 8113 20757 8125 20791
rect 8159 20788 8171 20791
rect 8202 20788 8208 20800
rect 8159 20760 8208 20788
rect 8159 20757 8171 20760
rect 8113 20751 8171 20757
rect 8202 20748 8208 20760
rect 8260 20748 8266 20800
rect 8294 20748 8300 20800
rect 8352 20788 8358 20800
rect 10042 20788 10048 20800
rect 8352 20760 10048 20788
rect 8352 20748 8358 20760
rect 10042 20748 10048 20760
rect 10100 20748 10106 20800
rect 10520 20788 10548 20819
rect 10594 20816 10600 20868
rect 10652 20816 10658 20868
rect 11241 20859 11299 20865
rect 11241 20825 11253 20859
rect 11287 20856 11299 20859
rect 11514 20856 11520 20868
rect 11287 20828 11520 20856
rect 11287 20825 11299 20828
rect 11241 20819 11299 20825
rect 11514 20816 11520 20828
rect 11572 20816 11578 20868
rect 12250 20816 12256 20868
rect 12308 20816 12314 20868
rect 12894 20856 12900 20868
rect 12728 20828 12900 20856
rect 12728 20788 12756 20828
rect 12894 20816 12900 20828
rect 12952 20856 12958 20868
rect 13541 20859 13599 20865
rect 13541 20856 13553 20859
rect 12952 20828 13553 20856
rect 12952 20816 12958 20828
rect 13541 20825 13553 20828
rect 13587 20825 13599 20859
rect 13740 20856 13768 20887
rect 13814 20884 13820 20936
rect 13872 20884 13878 20936
rect 14752 20933 14780 20964
rect 15470 20952 15476 20964
rect 15528 20952 15534 21004
rect 18966 20992 18972 21004
rect 18432 20964 18972 20992
rect 14461 20927 14519 20933
rect 14461 20893 14473 20927
rect 14507 20893 14519 20927
rect 14461 20887 14519 20893
rect 14645 20927 14703 20933
rect 14645 20893 14657 20927
rect 14691 20924 14703 20927
rect 14737 20927 14795 20933
rect 14737 20924 14749 20927
rect 14691 20896 14749 20924
rect 14691 20893 14703 20896
rect 14645 20887 14703 20893
rect 14737 20893 14749 20896
rect 14783 20893 14795 20927
rect 14737 20887 14795 20893
rect 14921 20927 14979 20933
rect 14921 20893 14933 20927
rect 14967 20924 14979 20927
rect 15654 20924 15660 20936
rect 14967 20896 15660 20924
rect 14967 20893 14979 20896
rect 14921 20887 14979 20893
rect 14476 20856 14504 20887
rect 14936 20856 14964 20887
rect 15654 20884 15660 20896
rect 15712 20884 15718 20936
rect 17034 20884 17040 20936
rect 17092 20884 17098 20936
rect 18230 20884 18236 20936
rect 18288 20924 18294 20936
rect 18432 20933 18460 20964
rect 18966 20952 18972 20964
rect 19024 20952 19030 21004
rect 19794 20952 19800 21004
rect 19852 20952 19858 21004
rect 23676 20992 23704 21032
rect 25038 21020 25044 21032
rect 25096 21020 25102 21072
rect 26234 21020 26240 21072
rect 26292 21060 26298 21072
rect 29638 21060 29644 21072
rect 26292 21032 29644 21060
rect 26292 21020 26298 21032
rect 29638 21020 29644 21032
rect 29696 21060 29702 21072
rect 34790 21060 34796 21072
rect 29696 21032 34796 21060
rect 29696 21020 29702 21032
rect 34790 21020 34796 21032
rect 34848 21060 34854 21072
rect 35710 21060 35716 21072
rect 34848 21032 35716 21060
rect 34848 21020 34854 21032
rect 35710 21020 35716 21032
rect 35768 21020 35774 21072
rect 36078 21020 36084 21072
rect 36136 21060 36142 21072
rect 36556 21060 36584 21091
rect 36998 21088 37004 21140
rect 37056 21088 37062 21140
rect 36136 21032 36584 21060
rect 36136 21020 36142 21032
rect 20272 20964 23704 20992
rect 23753 20995 23811 21001
rect 18417 20927 18475 20933
rect 18417 20924 18429 20927
rect 18288 20896 18429 20924
rect 18288 20884 18294 20896
rect 18417 20893 18429 20896
rect 18463 20893 18475 20927
rect 18417 20887 18475 20893
rect 18506 20884 18512 20936
rect 18564 20884 18570 20936
rect 18693 20927 18751 20933
rect 18693 20893 18705 20927
rect 18739 20924 18751 20927
rect 18739 20896 19564 20924
rect 18739 20893 18751 20896
rect 18693 20887 18751 20893
rect 13740 20828 14412 20856
rect 14476 20828 14964 20856
rect 17313 20859 17371 20865
rect 13541 20819 13599 20825
rect 14384 20800 14412 20828
rect 17313 20825 17325 20859
rect 17359 20856 17371 20859
rect 18598 20856 18604 20868
rect 17359 20828 18604 20856
rect 17359 20825 17371 20828
rect 17313 20819 17371 20825
rect 18598 20816 18604 20828
rect 18656 20816 18662 20868
rect 18782 20816 18788 20868
rect 18840 20856 18846 20868
rect 19245 20859 19303 20865
rect 19245 20856 19257 20859
rect 18840 20828 19257 20856
rect 18840 20816 18846 20828
rect 19245 20825 19257 20828
rect 19291 20825 19303 20859
rect 19536 20856 19564 20896
rect 19610 20884 19616 20936
rect 19668 20924 19674 20936
rect 20272 20933 20300 20964
rect 23753 20961 23765 20995
rect 23799 20992 23811 20995
rect 28350 20992 28356 21004
rect 23799 20964 28356 20992
rect 23799 20961 23811 20964
rect 23753 20955 23811 20961
rect 28350 20952 28356 20964
rect 28408 20952 28414 21004
rect 30116 20964 31800 20992
rect 19889 20927 19947 20933
rect 19889 20924 19901 20927
rect 19668 20896 19901 20924
rect 19668 20884 19674 20896
rect 19889 20893 19901 20896
rect 19935 20893 19947 20927
rect 19889 20887 19947 20893
rect 20257 20927 20315 20933
rect 20257 20893 20269 20927
rect 20303 20893 20315 20927
rect 20257 20887 20315 20893
rect 20438 20884 20444 20936
rect 20496 20884 20502 20936
rect 20622 20884 20628 20936
rect 20680 20924 20686 20936
rect 23566 20924 23572 20936
rect 20680 20896 23572 20924
rect 20680 20884 20686 20896
rect 23566 20884 23572 20896
rect 23624 20884 23630 20936
rect 23845 20927 23903 20933
rect 23845 20893 23857 20927
rect 23891 20924 23903 20927
rect 28813 20927 28871 20933
rect 28813 20924 28825 20927
rect 23891 20896 28825 20924
rect 23891 20893 23903 20896
rect 23845 20887 23903 20893
rect 28813 20893 28825 20896
rect 28859 20893 28871 20927
rect 28813 20887 28871 20893
rect 28902 20884 28908 20936
rect 28960 20884 28966 20936
rect 28997 20927 29055 20933
rect 28997 20893 29009 20927
rect 29043 20924 29055 20927
rect 29086 20924 29092 20936
rect 29043 20896 29092 20924
rect 29043 20893 29055 20896
rect 28997 20887 29055 20893
rect 29086 20884 29092 20896
rect 29144 20884 29150 20936
rect 29914 20884 29920 20936
rect 29972 20884 29978 20936
rect 30006 20884 30012 20936
rect 30064 20924 30070 20936
rect 30116 20933 30144 20964
rect 30101 20927 30159 20933
rect 30101 20924 30113 20927
rect 30064 20896 30113 20924
rect 30064 20884 30070 20896
rect 30101 20893 30113 20896
rect 30147 20893 30159 20927
rect 30101 20887 30159 20893
rect 30193 20927 30251 20933
rect 30193 20893 30205 20927
rect 30239 20924 30251 20927
rect 30466 20924 30472 20936
rect 30239 20896 30472 20924
rect 30239 20893 30251 20896
rect 30193 20887 30251 20893
rect 30466 20884 30472 20896
rect 30524 20884 30530 20936
rect 19536 20828 20576 20856
rect 19245 20819 19303 20825
rect 10520 20760 12756 20788
rect 12802 20748 12808 20800
rect 12860 20748 12866 20800
rect 13906 20748 13912 20800
rect 13964 20788 13970 20800
rect 14277 20791 14335 20797
rect 14277 20788 14289 20791
rect 13964 20760 14289 20788
rect 13964 20748 13970 20760
rect 14277 20757 14289 20760
rect 14323 20757 14335 20791
rect 14277 20751 14335 20757
rect 14366 20748 14372 20800
rect 14424 20788 14430 20800
rect 14737 20791 14795 20797
rect 14737 20788 14749 20791
rect 14424 20760 14749 20788
rect 14424 20748 14430 20760
rect 14737 20757 14749 20760
rect 14783 20757 14795 20791
rect 14737 20751 14795 20757
rect 16114 20748 16120 20800
rect 16172 20788 16178 20800
rect 16850 20788 16856 20800
rect 16172 20760 16856 20788
rect 16172 20748 16178 20760
rect 16850 20748 16856 20760
rect 16908 20748 16914 20800
rect 17129 20791 17187 20797
rect 17129 20757 17141 20791
rect 17175 20788 17187 20791
rect 17402 20788 17408 20800
rect 17175 20760 17408 20788
rect 17175 20757 17187 20760
rect 17129 20751 17187 20757
rect 17402 20748 17408 20760
rect 17460 20788 17466 20800
rect 18690 20788 18696 20800
rect 17460 20760 18696 20788
rect 17460 20748 17466 20760
rect 18690 20748 18696 20760
rect 18748 20788 18754 20800
rect 18966 20788 18972 20800
rect 18748 20760 18972 20788
rect 18748 20748 18754 20760
rect 18966 20748 18972 20760
rect 19024 20748 19030 20800
rect 20548 20788 20576 20828
rect 20806 20816 20812 20868
rect 20864 20816 20870 20868
rect 21726 20816 21732 20868
rect 21784 20856 21790 20868
rect 23934 20856 23940 20868
rect 21784 20828 23940 20856
rect 21784 20816 21790 20828
rect 23934 20816 23940 20828
rect 23992 20816 23998 20868
rect 25958 20816 25964 20868
rect 26016 20856 26022 20868
rect 26237 20859 26295 20865
rect 26237 20856 26249 20859
rect 26016 20828 26249 20856
rect 26016 20816 26022 20828
rect 26237 20825 26249 20828
rect 26283 20825 26295 20859
rect 26237 20819 26295 20825
rect 26421 20859 26479 20865
rect 26421 20825 26433 20859
rect 26467 20856 26479 20859
rect 27614 20856 27620 20868
rect 26467 20828 27620 20856
rect 26467 20825 26479 20828
rect 26421 20819 26479 20825
rect 27614 20816 27620 20828
rect 27672 20816 27678 20868
rect 27706 20816 27712 20868
rect 27764 20856 27770 20868
rect 28350 20856 28356 20868
rect 27764 20828 28356 20856
rect 27764 20816 27770 20828
rect 28350 20816 28356 20828
rect 28408 20816 28414 20868
rect 28718 20816 28724 20868
rect 28776 20856 28782 20868
rect 29181 20859 29239 20865
rect 29181 20856 29193 20859
rect 28776 20828 29193 20856
rect 28776 20816 28782 20828
rect 20898 20788 20904 20800
rect 20548 20760 20904 20788
rect 20898 20748 20904 20760
rect 20956 20748 20962 20800
rect 21542 20748 21548 20800
rect 21600 20788 21606 20800
rect 21818 20788 21824 20800
rect 21600 20760 21824 20788
rect 21600 20748 21606 20760
rect 21818 20748 21824 20760
rect 21876 20748 21882 20800
rect 22002 20748 22008 20800
rect 22060 20788 22066 20800
rect 22097 20791 22155 20797
rect 22097 20788 22109 20791
rect 22060 20760 22109 20788
rect 22060 20748 22066 20760
rect 22097 20757 22109 20760
rect 22143 20757 22155 20791
rect 22097 20751 22155 20757
rect 26602 20748 26608 20800
rect 26660 20748 26666 20800
rect 28368 20788 28396 20816
rect 29012 20800 29040 20828
rect 29181 20825 29193 20828
rect 29227 20825 29239 20859
rect 29181 20819 29239 20825
rect 29273 20859 29331 20865
rect 29273 20825 29285 20859
rect 29319 20856 29331 20859
rect 29733 20859 29791 20865
rect 29733 20856 29745 20859
rect 29319 20828 29745 20856
rect 29319 20825 29331 20828
rect 29273 20819 29331 20825
rect 29733 20825 29745 20828
rect 29779 20825 29791 20859
rect 29733 20819 29791 20825
rect 30282 20816 30288 20868
rect 30340 20856 30346 20868
rect 31205 20859 31263 20865
rect 31205 20856 31217 20859
rect 30340 20828 31217 20856
rect 30340 20816 30346 20828
rect 31205 20825 31217 20828
rect 31251 20825 31263 20859
rect 31772 20856 31800 20964
rect 32490 20952 32496 21004
rect 32548 20952 32554 21004
rect 33042 20952 33048 21004
rect 33100 20992 33106 21004
rect 33100 20964 35756 20992
rect 33100 20952 33106 20964
rect 31846 20884 31852 20936
rect 31904 20924 31910 20936
rect 32214 20924 32220 20936
rect 31904 20896 32220 20924
rect 31904 20884 31910 20896
rect 32214 20884 32220 20896
rect 32272 20884 32278 20936
rect 32858 20884 32864 20936
rect 32916 20924 32922 20936
rect 33689 20927 33747 20933
rect 33689 20924 33701 20927
rect 32916 20896 33701 20924
rect 32916 20884 32922 20896
rect 33689 20893 33701 20896
rect 33735 20893 33747 20927
rect 33689 20887 33747 20893
rect 33778 20884 33784 20936
rect 33836 20884 33842 20936
rect 34149 20927 34207 20933
rect 34149 20893 34161 20927
rect 34195 20924 34207 20927
rect 34422 20924 34428 20936
rect 34195 20896 34428 20924
rect 34195 20893 34207 20896
rect 34149 20887 34207 20893
rect 34422 20884 34428 20896
rect 34480 20884 34486 20936
rect 35728 20933 35756 20964
rect 36170 20952 36176 21004
rect 36228 20992 36234 21004
rect 36725 20995 36783 21001
rect 36725 20992 36737 20995
rect 36228 20964 36737 20992
rect 36228 20952 36234 20964
rect 36725 20961 36737 20964
rect 36771 20992 36783 20995
rect 36998 20992 37004 21004
rect 36771 20964 37004 20992
rect 36771 20961 36783 20964
rect 36725 20955 36783 20961
rect 36998 20952 37004 20964
rect 37056 20952 37062 21004
rect 35713 20927 35771 20933
rect 35713 20893 35725 20927
rect 35759 20893 35771 20927
rect 36354 20924 36360 20936
rect 35713 20887 35771 20893
rect 35820 20896 36360 20924
rect 33796 20856 33824 20884
rect 31772 20828 33824 20856
rect 31205 20819 31263 20825
rect 33870 20816 33876 20868
rect 33928 20816 33934 20868
rect 34011 20859 34069 20865
rect 34011 20825 34023 20859
rect 34057 20856 34069 20859
rect 35820 20856 35848 20896
rect 36354 20884 36360 20896
rect 36412 20884 36418 20936
rect 36817 20927 36875 20933
rect 36817 20893 36829 20927
rect 36863 20924 36875 20927
rect 37274 20924 37280 20936
rect 36863 20896 37280 20924
rect 36863 20893 36875 20896
rect 36817 20887 36875 20893
rect 37274 20884 37280 20896
rect 37332 20924 37338 20936
rect 38102 20924 38108 20936
rect 37332 20896 38108 20924
rect 37332 20884 37338 20896
rect 38102 20884 38108 20896
rect 38160 20884 38166 20936
rect 38470 20884 38476 20936
rect 38528 20924 38534 20936
rect 38749 20927 38807 20933
rect 38749 20924 38761 20927
rect 38528 20896 38761 20924
rect 38528 20884 38534 20896
rect 38749 20893 38761 20896
rect 38795 20893 38807 20927
rect 38749 20887 38807 20893
rect 34057 20828 35848 20856
rect 34057 20825 34069 20828
rect 34011 20819 34069 20825
rect 36262 20816 36268 20868
rect 36320 20856 36326 20868
rect 36541 20859 36599 20865
rect 36541 20856 36553 20859
rect 36320 20828 36553 20856
rect 36320 20816 36326 20828
rect 36541 20825 36553 20828
rect 36587 20825 36599 20859
rect 36541 20819 36599 20825
rect 38286 20816 38292 20868
rect 38344 20856 38350 20868
rect 38838 20856 38844 20868
rect 38344 20828 38844 20856
rect 38344 20816 38350 20828
rect 38838 20816 38844 20828
rect 38896 20816 38902 20868
rect 28810 20788 28816 20800
rect 28368 20760 28816 20788
rect 28810 20748 28816 20760
rect 28868 20748 28874 20800
rect 28994 20748 29000 20800
rect 29052 20748 29058 20800
rect 30466 20748 30472 20800
rect 30524 20788 30530 20800
rect 31297 20791 31355 20797
rect 31297 20788 31309 20791
rect 30524 20760 31309 20788
rect 30524 20748 30530 20760
rect 31297 20757 31309 20760
rect 31343 20757 31355 20791
rect 31297 20751 31355 20757
rect 33502 20748 33508 20800
rect 33560 20748 33566 20800
rect 35250 20748 35256 20800
rect 35308 20788 35314 20800
rect 35894 20788 35900 20800
rect 35308 20760 35900 20788
rect 35308 20748 35314 20760
rect 35894 20748 35900 20760
rect 35952 20788 35958 20800
rect 37274 20788 37280 20800
rect 35952 20760 37280 20788
rect 35952 20748 35958 20760
rect 37274 20748 37280 20760
rect 37332 20748 37338 20800
rect 38378 20748 38384 20800
rect 38436 20788 38442 20800
rect 38473 20791 38531 20797
rect 38473 20788 38485 20791
rect 38436 20760 38485 20788
rect 38436 20748 38442 20760
rect 38473 20757 38485 20760
rect 38519 20757 38531 20791
rect 38473 20751 38531 20757
rect 1104 20698 40572 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 40572 20698
rect 1104 20624 40572 20646
rect 1578 20544 1584 20596
rect 1636 20584 1642 20596
rect 5261 20587 5319 20593
rect 1636 20556 3556 20584
rect 1636 20544 1642 20556
rect 3050 20408 3056 20460
rect 3108 20408 3114 20460
rect 2774 20340 2780 20392
rect 2832 20380 2838 20392
rect 3142 20380 3148 20392
rect 2832 20352 3148 20380
rect 2832 20340 2838 20352
rect 3142 20340 3148 20352
rect 3200 20340 3206 20392
rect 3326 20340 3332 20392
rect 3384 20340 3390 20392
rect 3528 20389 3556 20556
rect 5261 20553 5273 20587
rect 5307 20584 5319 20587
rect 5350 20584 5356 20596
rect 5307 20556 5356 20584
rect 5307 20553 5319 20556
rect 5261 20547 5319 20553
rect 5350 20544 5356 20556
rect 5408 20544 5414 20596
rect 5905 20587 5963 20593
rect 5905 20553 5917 20587
rect 5951 20584 5963 20587
rect 5994 20584 6000 20596
rect 5951 20556 6000 20584
rect 5951 20553 5963 20556
rect 5905 20547 5963 20553
rect 5994 20544 6000 20556
rect 6052 20544 6058 20596
rect 6362 20544 6368 20596
rect 6420 20544 6426 20596
rect 10321 20587 10379 20593
rect 10321 20553 10333 20587
rect 10367 20584 10379 20587
rect 10594 20584 10600 20596
rect 10367 20556 10600 20584
rect 10367 20553 10379 20556
rect 10321 20547 10379 20553
rect 10594 20544 10600 20556
rect 10652 20544 10658 20596
rect 11514 20544 11520 20596
rect 11572 20584 11578 20596
rect 11793 20587 11851 20593
rect 11793 20584 11805 20587
rect 11572 20556 11805 20584
rect 11572 20544 11578 20556
rect 11793 20553 11805 20556
rect 11839 20553 11851 20587
rect 11793 20547 11851 20553
rect 12161 20587 12219 20593
rect 12161 20553 12173 20587
rect 12207 20584 12219 20587
rect 12802 20584 12808 20596
rect 12207 20556 12808 20584
rect 12207 20553 12219 20556
rect 12161 20547 12219 20553
rect 12802 20544 12808 20556
rect 12860 20544 12866 20596
rect 15841 20587 15899 20593
rect 15841 20584 15853 20587
rect 13188 20556 15853 20584
rect 3786 20476 3792 20528
rect 3844 20516 3850 20528
rect 3844 20488 4278 20516
rect 3844 20476 3850 20488
rect 5534 20476 5540 20528
rect 5592 20476 5598 20528
rect 5626 20476 5632 20528
rect 5684 20476 5690 20528
rect 7098 20516 7104 20528
rect 6564 20488 7104 20516
rect 5258 20408 5264 20460
rect 5316 20448 5322 20460
rect 5353 20451 5411 20457
rect 5353 20448 5365 20451
rect 5316 20420 5365 20448
rect 5316 20408 5322 20420
rect 5353 20417 5365 20420
rect 5399 20417 5411 20451
rect 5353 20411 5411 20417
rect 5718 20408 5724 20460
rect 5776 20408 5782 20460
rect 6564 20457 6592 20488
rect 7098 20476 7104 20488
rect 7156 20476 7162 20528
rect 9490 20476 9496 20528
rect 9548 20476 9554 20528
rect 6549 20451 6607 20457
rect 6549 20417 6561 20451
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 6733 20451 6791 20457
rect 6733 20417 6745 20451
rect 6779 20417 6791 20451
rect 6733 20411 6791 20417
rect 6825 20451 6883 20457
rect 6825 20417 6837 20451
rect 6871 20417 6883 20451
rect 10612 20448 10640 20544
rect 12253 20519 12311 20525
rect 12253 20485 12265 20519
rect 12299 20516 12311 20519
rect 13078 20516 13084 20528
rect 12299 20488 13084 20516
rect 12299 20485 12311 20488
rect 12253 20479 12311 20485
rect 12820 20460 12848 20488
rect 13078 20476 13084 20488
rect 13136 20476 13142 20528
rect 10965 20451 11023 20457
rect 10965 20448 10977 20451
rect 10612 20420 10977 20448
rect 6825 20411 6883 20417
rect 10965 20417 10977 20420
rect 11011 20417 11023 20451
rect 10965 20411 11023 20417
rect 3513 20383 3571 20389
rect 3513 20349 3525 20383
rect 3559 20380 3571 20383
rect 3789 20383 3847 20389
rect 3559 20352 3648 20380
rect 3559 20349 3571 20352
rect 3513 20343 3571 20349
rect 2130 20272 2136 20324
rect 2188 20312 2194 20324
rect 2685 20315 2743 20321
rect 2685 20312 2697 20315
rect 2188 20284 2697 20312
rect 2188 20272 2194 20284
rect 2685 20281 2697 20284
rect 2731 20281 2743 20315
rect 2685 20275 2743 20281
rect 3620 20244 3648 20352
rect 3789 20349 3801 20383
rect 3835 20380 3847 20383
rect 4430 20380 4436 20392
rect 3835 20352 4436 20380
rect 3835 20349 3847 20352
rect 3789 20343 3847 20349
rect 4430 20340 4436 20352
rect 4488 20340 4494 20392
rect 5442 20340 5448 20392
rect 5500 20380 5506 20392
rect 6748 20380 6776 20411
rect 5500 20352 6776 20380
rect 5500 20340 5506 20352
rect 6638 20272 6644 20324
rect 6696 20312 6702 20324
rect 6840 20312 6868 20411
rect 12802 20408 12808 20460
rect 12860 20408 12866 20460
rect 8570 20340 8576 20392
rect 8628 20340 8634 20392
rect 8849 20383 8907 20389
rect 8849 20349 8861 20383
rect 8895 20380 8907 20383
rect 9306 20380 9312 20392
rect 8895 20352 9312 20380
rect 8895 20349 8907 20352
rect 8849 20343 8907 20349
rect 9306 20340 9312 20352
rect 9364 20340 9370 20392
rect 12345 20383 12403 20389
rect 12345 20349 12357 20383
rect 12391 20349 12403 20383
rect 12345 20343 12403 20349
rect 6696 20284 6868 20312
rect 6696 20272 6702 20284
rect 9858 20272 9864 20324
rect 9916 20312 9922 20324
rect 12360 20312 12388 20343
rect 13188 20312 13216 20556
rect 15841 20553 15853 20556
rect 15887 20553 15899 20587
rect 15841 20547 15899 20553
rect 18601 20587 18659 20593
rect 18601 20553 18613 20587
rect 18647 20584 18659 20587
rect 19794 20584 19800 20596
rect 18647 20556 19800 20584
rect 18647 20553 18659 20556
rect 18601 20547 18659 20553
rect 19794 20544 19800 20556
rect 19852 20544 19858 20596
rect 23032 20556 24992 20584
rect 13906 20516 13912 20528
rect 13372 20488 13912 20516
rect 13372 20457 13400 20488
rect 13906 20476 13912 20488
rect 13964 20476 13970 20528
rect 14093 20519 14151 20525
rect 14093 20485 14105 20519
rect 14139 20516 14151 20519
rect 14274 20516 14280 20528
rect 14139 20488 14280 20516
rect 14139 20485 14151 20488
rect 14093 20479 14151 20485
rect 14274 20476 14280 20488
rect 14332 20476 14338 20528
rect 17126 20476 17132 20528
rect 17184 20516 17190 20528
rect 18233 20519 18291 20525
rect 18233 20516 18245 20519
rect 17184 20488 18245 20516
rect 17184 20476 17190 20488
rect 18233 20485 18245 20488
rect 18279 20485 18291 20519
rect 18233 20479 18291 20485
rect 18322 20476 18328 20528
rect 18380 20516 18386 20528
rect 18433 20519 18491 20525
rect 18433 20516 18445 20519
rect 18380 20488 18445 20516
rect 18380 20476 18386 20488
rect 18433 20485 18445 20488
rect 18479 20485 18491 20519
rect 18433 20479 18491 20485
rect 22002 20476 22008 20528
rect 22060 20516 22066 20528
rect 23032 20516 23060 20556
rect 22060 20488 23060 20516
rect 22060 20476 22066 20488
rect 23106 20476 23112 20528
rect 23164 20476 23170 20528
rect 24964 20525 24992 20556
rect 26418 20544 26424 20596
rect 26476 20584 26482 20596
rect 26697 20587 26755 20593
rect 26697 20584 26709 20587
rect 26476 20556 26709 20584
rect 26476 20544 26482 20556
rect 26697 20553 26709 20556
rect 26743 20553 26755 20587
rect 30466 20584 30472 20596
rect 26697 20547 26755 20553
rect 27632 20556 30472 20584
rect 24949 20519 25007 20525
rect 24949 20485 24961 20519
rect 24995 20516 25007 20519
rect 25314 20516 25320 20528
rect 24995 20488 25320 20516
rect 24995 20485 25007 20488
rect 24949 20479 25007 20485
rect 25314 20476 25320 20488
rect 25372 20476 25378 20528
rect 25409 20519 25467 20525
rect 25409 20485 25421 20519
rect 25455 20516 25467 20519
rect 25866 20516 25872 20528
rect 25455 20488 25872 20516
rect 25455 20485 25467 20488
rect 25409 20479 25467 20485
rect 25866 20476 25872 20488
rect 25924 20476 25930 20528
rect 26524 20519 26582 20525
rect 26524 20485 26536 20519
rect 26570 20516 26582 20519
rect 26570 20488 27384 20516
rect 26570 20485 26582 20488
rect 26524 20479 26582 20485
rect 13357 20451 13415 20457
rect 13357 20417 13369 20451
rect 13403 20417 13415 20451
rect 13357 20411 13415 20417
rect 13541 20451 13599 20457
rect 13541 20417 13553 20451
rect 13587 20448 13599 20451
rect 13814 20448 13820 20460
rect 13587 20420 13820 20448
rect 13587 20417 13599 20420
rect 13541 20411 13599 20417
rect 13814 20408 13820 20420
rect 13872 20448 13878 20460
rect 13872 20420 14320 20448
rect 13872 20408 13878 20420
rect 14182 20340 14188 20392
rect 14240 20340 14246 20392
rect 14292 20380 14320 20420
rect 14366 20408 14372 20460
rect 14424 20408 14430 20460
rect 14458 20408 14464 20460
rect 14516 20448 14522 20460
rect 14737 20451 14795 20457
rect 14737 20448 14749 20451
rect 14516 20420 14749 20448
rect 14516 20408 14522 20420
rect 14737 20417 14749 20420
rect 14783 20417 14795 20451
rect 14737 20411 14795 20417
rect 15470 20408 15476 20460
rect 15528 20408 15534 20460
rect 15562 20408 15568 20460
rect 15620 20448 15626 20460
rect 15657 20451 15715 20457
rect 15657 20448 15669 20451
rect 15620 20420 15669 20448
rect 15620 20408 15626 20420
rect 15657 20417 15669 20420
rect 15703 20417 15715 20451
rect 15657 20411 15715 20417
rect 15746 20408 15752 20460
rect 15804 20408 15810 20460
rect 16298 20408 16304 20460
rect 16356 20408 16362 20460
rect 16390 20408 16396 20460
rect 16448 20448 16454 20460
rect 20901 20451 20959 20457
rect 16448 20420 20760 20448
rect 16448 20408 16454 20420
rect 14476 20380 14504 20408
rect 14292 20352 14504 20380
rect 14829 20383 14887 20389
rect 14829 20349 14841 20383
rect 14875 20380 14887 20383
rect 15010 20380 15016 20392
rect 14875 20352 15016 20380
rect 14875 20349 14887 20352
rect 14829 20343 14887 20349
rect 15010 20340 15016 20352
rect 15068 20340 15074 20392
rect 15102 20340 15108 20392
rect 15160 20340 15166 20392
rect 15764 20380 15792 20408
rect 16574 20380 16580 20392
rect 15764 20352 16580 20380
rect 16574 20340 16580 20352
rect 16632 20380 16638 20392
rect 17586 20380 17592 20392
rect 16632 20352 17592 20380
rect 16632 20340 16638 20352
rect 17586 20340 17592 20352
rect 17644 20340 17650 20392
rect 20622 20340 20628 20392
rect 20680 20340 20686 20392
rect 20732 20380 20760 20420
rect 20901 20417 20913 20451
rect 20947 20448 20959 20451
rect 21358 20448 21364 20460
rect 20947 20420 21364 20448
rect 20947 20417 20959 20420
rect 20901 20411 20959 20417
rect 21358 20408 21364 20420
rect 21416 20408 21422 20460
rect 22278 20408 22284 20460
rect 22336 20448 22342 20460
rect 22741 20451 22799 20457
rect 22741 20448 22753 20451
rect 22336 20420 22753 20448
rect 22336 20408 22342 20420
rect 22741 20417 22753 20420
rect 22787 20417 22799 20451
rect 22741 20411 22799 20417
rect 22830 20408 22836 20460
rect 22888 20408 22894 20460
rect 23017 20451 23075 20457
rect 23017 20417 23029 20451
rect 23063 20446 23075 20451
rect 23124 20446 23152 20476
rect 27356 20460 27384 20488
rect 23063 20418 23152 20446
rect 23063 20417 23075 20418
rect 23017 20411 23075 20417
rect 25038 20408 25044 20460
rect 25096 20408 25102 20460
rect 25501 20451 25559 20457
rect 25501 20448 25513 20451
rect 25332 20420 25513 20448
rect 23201 20383 23259 20389
rect 23201 20380 23213 20383
rect 20732 20352 23213 20380
rect 23201 20349 23213 20352
rect 23247 20349 23259 20383
rect 23201 20343 23259 20349
rect 23382 20340 23388 20392
rect 23440 20380 23446 20392
rect 24946 20380 24952 20392
rect 23440 20352 24952 20380
rect 23440 20340 23446 20352
rect 24946 20340 24952 20352
rect 25004 20340 25010 20392
rect 25130 20340 25136 20392
rect 25188 20380 25194 20392
rect 25332 20389 25360 20420
rect 25501 20417 25513 20420
rect 25547 20417 25559 20451
rect 25501 20411 25559 20417
rect 25682 20408 25688 20460
rect 25740 20448 25746 20460
rect 25777 20451 25835 20457
rect 25777 20448 25789 20451
rect 25740 20420 25789 20448
rect 25740 20408 25746 20420
rect 25777 20417 25789 20420
rect 25823 20448 25835 20451
rect 26237 20451 26295 20457
rect 26237 20448 26249 20451
rect 25823 20420 26249 20448
rect 25823 20417 25835 20420
rect 25777 20411 25835 20417
rect 26237 20417 26249 20420
rect 26283 20417 26295 20451
rect 26605 20451 26663 20457
rect 26605 20448 26617 20451
rect 26237 20411 26295 20417
rect 26344 20420 26617 20448
rect 25317 20383 25375 20389
rect 25317 20380 25329 20383
rect 25188 20352 25329 20380
rect 25188 20340 25194 20352
rect 25317 20349 25329 20352
rect 25363 20349 25375 20383
rect 25317 20343 25375 20349
rect 25593 20383 25651 20389
rect 25593 20349 25605 20383
rect 25639 20349 25651 20383
rect 26344 20380 26372 20420
rect 26605 20417 26617 20420
rect 26651 20417 26663 20451
rect 26605 20411 26663 20417
rect 26694 20408 26700 20460
rect 26752 20448 26758 20460
rect 26789 20451 26847 20457
rect 26789 20448 26801 20451
rect 26752 20420 26801 20448
rect 26752 20408 26758 20420
rect 26789 20417 26801 20420
rect 26835 20417 26847 20451
rect 26789 20411 26847 20417
rect 27338 20408 27344 20460
rect 27396 20408 27402 20460
rect 27430 20408 27436 20460
rect 27488 20408 27494 20460
rect 27632 20457 27660 20556
rect 30466 20544 30472 20556
rect 30524 20544 30530 20596
rect 33781 20587 33839 20593
rect 33781 20584 33793 20587
rect 30760 20556 33793 20584
rect 28718 20476 28724 20528
rect 28776 20476 28782 20528
rect 29730 20476 29736 20528
rect 29788 20516 29794 20528
rect 29788 20488 30144 20516
rect 29788 20476 29794 20488
rect 27617 20451 27675 20457
rect 27617 20417 27629 20451
rect 27663 20417 27675 20451
rect 27617 20411 27675 20417
rect 25593 20343 25651 20349
rect 26068 20352 26372 20380
rect 26421 20383 26479 20389
rect 9916 20284 13216 20312
rect 9916 20272 9922 20284
rect 13262 20272 13268 20324
rect 13320 20272 13326 20324
rect 15654 20272 15660 20324
rect 15712 20312 15718 20324
rect 20349 20315 20407 20321
rect 20349 20312 20361 20315
rect 15712 20284 20361 20312
rect 15712 20272 15718 20284
rect 20349 20281 20361 20284
rect 20395 20281 20407 20315
rect 20349 20275 20407 20281
rect 22925 20315 22983 20321
rect 22925 20281 22937 20315
rect 22971 20312 22983 20315
rect 23474 20312 23480 20324
rect 22971 20284 23480 20312
rect 22971 20281 22983 20284
rect 22925 20275 22983 20281
rect 23474 20272 23480 20284
rect 23532 20312 23538 20324
rect 23658 20312 23664 20324
rect 23532 20284 23664 20312
rect 23532 20272 23538 20284
rect 23658 20272 23664 20284
rect 23716 20272 23722 20324
rect 25225 20315 25283 20321
rect 25225 20281 25237 20315
rect 25271 20312 25283 20315
rect 25406 20312 25412 20324
rect 25271 20284 25412 20312
rect 25271 20281 25283 20284
rect 25225 20275 25283 20281
rect 25406 20272 25412 20284
rect 25464 20312 25470 20324
rect 25608 20312 25636 20343
rect 25464 20284 25636 20312
rect 25464 20272 25470 20284
rect 25958 20272 25964 20324
rect 26016 20272 26022 20324
rect 26068 20321 26096 20352
rect 26421 20349 26433 20383
rect 26467 20380 26479 20383
rect 26467 20352 27017 20380
rect 26467 20349 26479 20352
rect 26421 20343 26479 20349
rect 26053 20315 26111 20321
rect 26053 20281 26065 20315
rect 26099 20281 26111 20315
rect 26053 20275 26111 20281
rect 4798 20244 4804 20256
rect 3620 20216 4804 20244
rect 4798 20204 4804 20216
rect 4856 20204 4862 20256
rect 5626 20204 5632 20256
rect 5684 20244 5690 20256
rect 6546 20244 6552 20256
rect 5684 20216 6552 20244
rect 5684 20204 5690 20216
rect 6546 20204 6552 20216
rect 6604 20204 6610 20256
rect 9950 20204 9956 20256
rect 10008 20244 10014 20256
rect 10413 20247 10471 20253
rect 10413 20244 10425 20247
rect 10008 20216 10425 20244
rect 10008 20204 10014 20216
rect 10413 20213 10425 20216
rect 10459 20213 10471 20247
rect 10413 20207 10471 20213
rect 12986 20204 12992 20256
rect 13044 20244 13050 20256
rect 13725 20247 13783 20253
rect 13725 20244 13737 20247
rect 13044 20216 13737 20244
rect 13044 20204 13050 20216
rect 13725 20213 13737 20216
rect 13771 20213 13783 20247
rect 13725 20207 13783 20213
rect 13909 20247 13967 20253
rect 13909 20213 13921 20247
rect 13955 20244 13967 20247
rect 14090 20244 14096 20256
rect 13955 20216 14096 20244
rect 13955 20213 13967 20216
rect 13909 20207 13967 20213
rect 14090 20204 14096 20216
rect 14148 20244 14154 20256
rect 15565 20247 15623 20253
rect 15565 20244 15577 20247
rect 14148 20216 15577 20244
rect 14148 20204 14154 20216
rect 15565 20213 15577 20216
rect 15611 20213 15623 20247
rect 15565 20207 15623 20213
rect 18414 20204 18420 20256
rect 18472 20204 18478 20256
rect 20438 20204 20444 20256
rect 20496 20244 20502 20256
rect 20533 20247 20591 20253
rect 20533 20244 20545 20247
rect 20496 20216 20545 20244
rect 20496 20204 20502 20216
rect 20533 20213 20545 20216
rect 20579 20244 20591 20247
rect 23198 20244 23204 20256
rect 20579 20216 23204 20244
rect 20579 20213 20591 20216
rect 20533 20207 20591 20213
rect 23198 20204 23204 20216
rect 23256 20204 23262 20256
rect 24302 20204 24308 20256
rect 24360 20244 24366 20256
rect 25314 20244 25320 20256
rect 24360 20216 25320 20244
rect 24360 20204 24366 20216
rect 25314 20204 25320 20216
rect 25372 20204 25378 20256
rect 25498 20204 25504 20256
rect 25556 20244 25562 20256
rect 26237 20247 26295 20253
rect 26237 20244 26249 20247
rect 25556 20216 26249 20244
rect 25556 20204 25562 20216
rect 26237 20213 26249 20216
rect 26283 20213 26295 20247
rect 26989 20244 27017 20352
rect 27062 20340 27068 20392
rect 27120 20380 27126 20392
rect 27632 20380 27660 20411
rect 27706 20408 27712 20460
rect 27764 20408 27770 20460
rect 27893 20451 27951 20457
rect 27893 20417 27905 20451
rect 27939 20448 27951 20451
rect 27985 20451 28043 20457
rect 27985 20448 27997 20451
rect 27939 20420 27997 20448
rect 27939 20417 27951 20420
rect 27893 20411 27951 20417
rect 27985 20417 27997 20420
rect 28031 20417 28043 20451
rect 27985 20411 28043 20417
rect 28258 20408 28264 20460
rect 28316 20408 28322 20460
rect 28994 20408 29000 20460
rect 29052 20408 29058 20460
rect 29822 20408 29828 20460
rect 29880 20408 29886 20460
rect 29917 20451 29975 20457
rect 29917 20417 29929 20451
rect 29963 20448 29975 20451
rect 30006 20448 30012 20460
rect 29963 20420 30012 20448
rect 29963 20417 29975 20420
rect 29917 20411 29975 20417
rect 30006 20408 30012 20420
rect 30064 20408 30070 20460
rect 30116 20457 30144 20488
rect 30101 20451 30159 20457
rect 30101 20417 30113 20451
rect 30147 20417 30159 20451
rect 30101 20411 30159 20417
rect 30193 20451 30251 20457
rect 30193 20417 30205 20451
rect 30239 20446 30251 20451
rect 30760 20448 30788 20556
rect 33781 20553 33793 20556
rect 33827 20584 33839 20587
rect 33962 20584 33968 20596
rect 33827 20556 33968 20584
rect 33827 20553 33839 20556
rect 33781 20547 33839 20553
rect 33962 20544 33968 20556
rect 34020 20544 34026 20596
rect 30834 20476 30840 20528
rect 30892 20516 30898 20528
rect 31363 20519 31421 20525
rect 31363 20516 31375 20519
rect 30892 20488 31375 20516
rect 30892 20476 30898 20488
rect 31363 20485 31375 20488
rect 31409 20485 31421 20519
rect 31363 20479 31421 20485
rect 31754 20476 31760 20528
rect 31812 20516 31818 20528
rect 32769 20519 32827 20525
rect 32769 20516 32781 20519
rect 31812 20488 32781 20516
rect 31812 20476 31818 20488
rect 32769 20485 32781 20488
rect 32815 20485 32827 20519
rect 32769 20479 32827 20485
rect 36538 20476 36544 20528
rect 36596 20516 36602 20528
rect 38010 20516 38016 20528
rect 36596 20488 38016 20516
rect 36596 20476 36602 20488
rect 38010 20476 38016 20488
rect 38068 20516 38074 20528
rect 38378 20516 38384 20528
rect 38068 20488 38384 20516
rect 38068 20476 38074 20488
rect 38378 20476 38384 20488
rect 38436 20476 38442 20528
rect 30300 20446 30788 20448
rect 30239 20420 30788 20446
rect 30239 20418 30328 20420
rect 30239 20417 30251 20418
rect 30193 20411 30251 20417
rect 27120 20352 27660 20380
rect 27120 20340 27126 20352
rect 27798 20340 27804 20392
rect 27856 20380 27862 20392
rect 28074 20380 28080 20392
rect 27856 20352 28080 20380
rect 27856 20340 27862 20352
rect 28074 20340 28080 20352
rect 28132 20340 28138 20392
rect 28626 20340 28632 20392
rect 28684 20340 28690 20392
rect 29181 20383 29239 20389
rect 29181 20349 29193 20383
rect 29227 20380 29239 20383
rect 29641 20383 29699 20389
rect 29641 20380 29653 20383
rect 29227 20352 29653 20380
rect 29227 20349 29239 20352
rect 29181 20343 29239 20349
rect 29641 20349 29653 20352
rect 29687 20349 29699 20383
rect 29641 20343 29699 20349
rect 27522 20272 27528 20324
rect 27580 20312 27586 20324
rect 30300 20312 30328 20418
rect 31478 20408 31484 20460
rect 31536 20408 31542 20460
rect 31570 20408 31576 20460
rect 31628 20408 31634 20460
rect 31665 20451 31723 20457
rect 31665 20417 31677 20451
rect 31711 20448 31723 20451
rect 31846 20448 31852 20460
rect 31711 20420 31852 20448
rect 31711 20417 31723 20420
rect 31665 20411 31723 20417
rect 31846 20408 31852 20420
rect 31904 20408 31910 20460
rect 32030 20408 32036 20460
rect 32088 20448 32094 20460
rect 32490 20448 32496 20460
rect 32088 20420 32496 20448
rect 32088 20408 32094 20420
rect 32490 20408 32496 20420
rect 32548 20408 32554 20460
rect 32582 20408 32588 20460
rect 32640 20448 32646 20460
rect 32677 20451 32735 20457
rect 32677 20448 32689 20451
rect 32640 20420 32689 20448
rect 32640 20408 32646 20420
rect 32677 20417 32689 20420
rect 32723 20417 32735 20451
rect 32677 20411 32735 20417
rect 32858 20408 32864 20460
rect 32916 20408 32922 20460
rect 33594 20408 33600 20460
rect 33652 20448 33658 20460
rect 33965 20451 34023 20457
rect 33965 20448 33977 20451
rect 33652 20420 33977 20448
rect 33652 20408 33658 20420
rect 33965 20417 33977 20420
rect 34011 20448 34023 20451
rect 34698 20448 34704 20460
rect 34011 20420 34704 20448
rect 34011 20417 34023 20420
rect 33965 20411 34023 20417
rect 34698 20408 34704 20420
rect 34756 20408 34762 20460
rect 38102 20408 38108 20460
rect 38160 20408 38166 20460
rect 38198 20451 38256 20457
rect 38198 20417 38210 20451
rect 38244 20417 38256 20451
rect 38198 20411 38256 20417
rect 31202 20340 31208 20392
rect 31260 20340 31266 20392
rect 31754 20340 31760 20392
rect 31812 20380 31818 20392
rect 32876 20380 32904 20408
rect 31812 20352 32904 20380
rect 31812 20340 31818 20352
rect 33226 20340 33232 20392
rect 33284 20380 33290 20392
rect 33778 20380 33784 20392
rect 33284 20352 33784 20380
rect 33284 20340 33290 20352
rect 33778 20340 33784 20352
rect 33836 20380 33842 20392
rect 34149 20383 34207 20389
rect 34149 20380 34161 20383
rect 33836 20352 34161 20380
rect 33836 20340 33842 20352
rect 34149 20349 34161 20352
rect 34195 20349 34207 20383
rect 34149 20343 34207 20349
rect 37090 20340 37096 20392
rect 37148 20380 37154 20392
rect 37642 20380 37648 20392
rect 37148 20352 37648 20380
rect 37148 20340 37154 20352
rect 37642 20340 37648 20352
rect 37700 20380 37706 20392
rect 38212 20380 38240 20411
rect 38286 20408 38292 20460
rect 38344 20448 38350 20460
rect 38473 20451 38531 20457
rect 38473 20448 38485 20451
rect 38344 20420 38485 20448
rect 38344 20408 38350 20420
rect 38473 20417 38485 20420
rect 38519 20417 38531 20451
rect 38473 20411 38531 20417
rect 38570 20451 38628 20457
rect 38570 20417 38582 20451
rect 38616 20417 38628 20451
rect 38570 20411 38628 20417
rect 37700 20352 38240 20380
rect 37700 20340 37706 20352
rect 27580 20284 30328 20312
rect 27580 20272 27586 20284
rect 30926 20272 30932 20324
rect 30984 20312 30990 20324
rect 31478 20312 31484 20324
rect 30984 20284 31484 20312
rect 30984 20272 30990 20284
rect 31478 20272 31484 20284
rect 31536 20272 31542 20324
rect 34422 20272 34428 20324
rect 34480 20312 34486 20324
rect 35986 20312 35992 20324
rect 34480 20284 35992 20312
rect 34480 20272 34486 20284
rect 35986 20272 35992 20284
rect 36044 20272 36050 20324
rect 38010 20272 38016 20324
rect 38068 20312 38074 20324
rect 38580 20312 38608 20411
rect 38068 20284 38608 20312
rect 38068 20272 38074 20284
rect 27798 20244 27804 20256
rect 26989 20216 27804 20244
rect 26237 20207 26295 20213
rect 27798 20204 27804 20216
rect 27856 20204 27862 20256
rect 27982 20204 27988 20256
rect 28040 20204 28046 20256
rect 28442 20204 28448 20256
rect 28500 20204 28506 20256
rect 29822 20204 29828 20256
rect 29880 20244 29886 20256
rect 30650 20244 30656 20256
rect 29880 20216 30656 20244
rect 29880 20204 29886 20216
rect 30650 20204 30656 20216
rect 30708 20204 30714 20256
rect 30834 20204 30840 20256
rect 30892 20244 30898 20256
rect 31570 20244 31576 20256
rect 30892 20216 31576 20244
rect 30892 20204 30898 20216
rect 31570 20204 31576 20216
rect 31628 20204 31634 20256
rect 31754 20204 31760 20256
rect 31812 20244 31818 20256
rect 31849 20247 31907 20253
rect 31849 20244 31861 20247
rect 31812 20216 31861 20244
rect 31812 20204 31818 20216
rect 31849 20213 31861 20216
rect 31895 20213 31907 20247
rect 31849 20207 31907 20213
rect 32214 20204 32220 20256
rect 32272 20244 32278 20256
rect 32858 20244 32864 20256
rect 32272 20216 32864 20244
rect 32272 20204 32278 20216
rect 32858 20204 32864 20216
rect 32916 20204 32922 20256
rect 33042 20204 33048 20256
rect 33100 20204 33106 20256
rect 33962 20204 33968 20256
rect 34020 20244 34026 20256
rect 35250 20244 35256 20256
rect 34020 20216 35256 20244
rect 34020 20204 34026 20216
rect 35250 20204 35256 20216
rect 35308 20204 35314 20256
rect 38749 20247 38807 20253
rect 38749 20213 38761 20247
rect 38795 20244 38807 20247
rect 39298 20244 39304 20256
rect 38795 20216 39304 20244
rect 38795 20213 38807 20216
rect 38749 20207 38807 20213
rect 39298 20204 39304 20216
rect 39356 20244 39362 20256
rect 39574 20244 39580 20256
rect 39356 20216 39580 20244
rect 39356 20204 39362 20216
rect 39574 20204 39580 20216
rect 39632 20204 39638 20256
rect 1104 20154 40572 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 40572 20154
rect 1104 20080 40572 20102
rect 3050 20000 3056 20052
rect 3108 20040 3114 20052
rect 3789 20043 3847 20049
rect 3789 20040 3801 20043
rect 3108 20012 3801 20040
rect 3108 20000 3114 20012
rect 3789 20009 3801 20012
rect 3835 20009 3847 20043
rect 3789 20003 3847 20009
rect 5810 20000 5816 20052
rect 5868 20040 5874 20052
rect 6089 20043 6147 20049
rect 6089 20040 6101 20043
rect 5868 20012 6101 20040
rect 5868 20000 5874 20012
rect 6089 20009 6101 20012
rect 6135 20009 6147 20043
rect 6089 20003 6147 20009
rect 6730 20000 6736 20052
rect 6788 20000 6794 20052
rect 7098 20000 7104 20052
rect 7156 20040 7162 20052
rect 7834 20040 7840 20052
rect 7156 20012 7840 20040
rect 7156 20000 7162 20012
rect 7834 20000 7840 20012
rect 7892 20000 7898 20052
rect 8018 20000 8024 20052
rect 8076 20000 8082 20052
rect 9306 20000 9312 20052
rect 9364 20000 9370 20052
rect 10137 20043 10195 20049
rect 10137 20009 10149 20043
rect 10183 20040 10195 20043
rect 10226 20040 10232 20052
rect 10183 20012 10232 20040
rect 10183 20009 10195 20012
rect 10137 20003 10195 20009
rect 10226 20000 10232 20012
rect 10284 20000 10290 20052
rect 13538 20000 13544 20052
rect 13596 20000 13602 20052
rect 13630 20000 13636 20052
rect 13688 20040 13694 20052
rect 13725 20043 13783 20049
rect 13725 20040 13737 20043
rect 13688 20012 13737 20040
rect 13688 20000 13694 20012
rect 13725 20009 13737 20012
rect 13771 20009 13783 20043
rect 13725 20003 13783 20009
rect 14182 20000 14188 20052
rect 14240 20040 14246 20052
rect 14369 20043 14427 20049
rect 14369 20040 14381 20043
rect 14240 20012 14381 20040
rect 14240 20000 14246 20012
rect 14369 20009 14381 20012
rect 14415 20009 14427 20043
rect 14369 20003 14427 20009
rect 14458 20000 14464 20052
rect 14516 20000 14522 20052
rect 15378 20040 15384 20052
rect 14752 20012 15384 20040
rect 5718 19932 5724 19984
rect 5776 19972 5782 19984
rect 6362 19972 6368 19984
rect 5776 19944 6368 19972
rect 5776 19932 5782 19944
rect 6362 19932 6368 19944
rect 6420 19932 6426 19984
rect 6454 19932 6460 19984
rect 6512 19972 6518 19984
rect 6825 19975 6883 19981
rect 6825 19972 6837 19975
rect 6512 19944 6837 19972
rect 6512 19932 6518 19944
rect 6825 19941 6837 19944
rect 6871 19941 6883 19975
rect 6825 19935 6883 19941
rect 7300 19944 10364 19972
rect 3602 19864 3608 19916
rect 3660 19904 3666 19916
rect 4341 19907 4399 19913
rect 4341 19904 4353 19907
rect 3660 19876 4353 19904
rect 3660 19864 3666 19876
rect 4341 19873 4353 19876
rect 4387 19873 4399 19907
rect 7098 19904 7104 19916
rect 4341 19867 4399 19873
rect 5092 19876 6500 19904
rect 3418 19796 3424 19848
rect 3476 19836 3482 19848
rect 5092 19845 5120 19876
rect 5077 19839 5135 19845
rect 5077 19836 5089 19839
rect 3476 19808 5089 19836
rect 3476 19796 3482 19808
rect 5077 19805 5089 19808
rect 5123 19805 5135 19839
rect 5077 19799 5135 19805
rect 5537 19839 5595 19845
rect 5537 19805 5549 19839
rect 5583 19836 5595 19839
rect 5626 19836 5632 19848
rect 5583 19808 5632 19836
rect 5583 19805 5595 19808
rect 5537 19799 5595 19805
rect 5626 19796 5632 19808
rect 5684 19796 5690 19848
rect 5718 19796 5724 19848
rect 5776 19796 5782 19848
rect 5905 19839 5963 19845
rect 5905 19805 5917 19839
rect 5951 19805 5963 19839
rect 5905 19799 5963 19805
rect 5813 19771 5871 19777
rect 5813 19737 5825 19771
rect 5859 19737 5871 19771
rect 5920 19768 5948 19799
rect 6178 19796 6184 19848
rect 6236 19796 6242 19848
rect 6362 19796 6368 19848
rect 6420 19796 6426 19848
rect 6472 19845 6500 19876
rect 7024 19876 7104 19904
rect 6457 19839 6515 19845
rect 6457 19805 6469 19839
rect 6503 19805 6515 19839
rect 6457 19799 6515 19805
rect 6549 19839 6607 19845
rect 6549 19805 6561 19839
rect 6595 19805 6607 19839
rect 6549 19799 6607 19805
rect 6564 19768 6592 19799
rect 6730 19796 6736 19848
rect 6788 19836 6794 19848
rect 7024 19845 7052 19876
rect 7098 19864 7104 19876
rect 7156 19864 7162 19916
rect 7300 19845 7328 19944
rect 8662 19904 8668 19916
rect 8348 19876 8668 19904
rect 7009 19839 7067 19845
rect 7009 19836 7021 19839
rect 6788 19808 7021 19836
rect 6788 19796 6794 19808
rect 7009 19805 7021 19808
rect 7055 19805 7067 19839
rect 7009 19799 7067 19805
rect 7285 19839 7343 19845
rect 7285 19805 7297 19839
rect 7331 19836 7343 19839
rect 7561 19839 7619 19845
rect 7561 19836 7573 19839
rect 7331 19808 7573 19836
rect 7331 19805 7343 19808
rect 7285 19799 7343 19805
rect 7561 19805 7573 19808
rect 7607 19805 7619 19839
rect 7561 19799 7619 19805
rect 6638 19768 6644 19780
rect 5920 19740 6644 19768
rect 5813 19731 5871 19737
rect 3878 19660 3884 19712
rect 3936 19700 3942 19712
rect 4525 19703 4583 19709
rect 4525 19700 4537 19703
rect 3936 19672 4537 19700
rect 3936 19660 3942 19672
rect 4525 19669 4537 19672
rect 4571 19669 4583 19703
rect 4525 19663 4583 19669
rect 5258 19660 5264 19712
rect 5316 19700 5322 19712
rect 5828 19700 5856 19731
rect 6638 19728 6644 19740
rect 6696 19768 6702 19780
rect 7300 19768 7328 19799
rect 7834 19796 7840 19848
rect 7892 19796 7898 19848
rect 6696 19740 7328 19768
rect 7653 19771 7711 19777
rect 6696 19728 6702 19740
rect 7653 19737 7665 19771
rect 7699 19768 7711 19771
rect 8348 19768 8376 19876
rect 8662 19864 8668 19876
rect 8720 19904 8726 19916
rect 8757 19907 8815 19913
rect 8757 19904 8769 19907
rect 8720 19876 8769 19904
rect 8720 19864 8726 19876
rect 8757 19873 8769 19876
rect 8803 19873 8815 19907
rect 8757 19867 8815 19873
rect 9766 19864 9772 19916
rect 9824 19864 9830 19916
rect 9858 19864 9864 19916
rect 9916 19864 9922 19916
rect 10336 19904 10364 19944
rect 10686 19932 10692 19984
rect 10744 19972 10750 19984
rect 10870 19972 10876 19984
rect 10744 19944 10876 19972
rect 10744 19932 10750 19944
rect 10870 19932 10876 19944
rect 10928 19932 10934 19984
rect 13173 19975 13231 19981
rect 13173 19941 13185 19975
rect 13219 19972 13231 19975
rect 13354 19972 13360 19984
rect 13219 19944 13360 19972
rect 13219 19941 13231 19944
rect 13173 19935 13231 19941
rect 13354 19932 13360 19944
rect 13412 19932 13418 19984
rect 14752 19972 14780 20012
rect 15378 20000 15384 20012
rect 15436 20000 15442 20052
rect 20073 20043 20131 20049
rect 20073 20009 20085 20043
rect 20119 20040 20131 20043
rect 20162 20040 20168 20052
rect 20119 20012 20168 20040
rect 20119 20009 20131 20012
rect 20073 20003 20131 20009
rect 20162 20000 20168 20012
rect 20220 20000 20226 20052
rect 20272 20012 21680 20040
rect 15470 19972 15476 19984
rect 14108 19944 14780 19972
rect 12526 19904 12532 19916
rect 10336 19876 12532 19904
rect 9677 19839 9735 19845
rect 9677 19805 9689 19839
rect 9723 19836 9735 19839
rect 9950 19836 9956 19848
rect 9723 19808 9956 19836
rect 9723 19805 9735 19808
rect 9677 19799 9735 19805
rect 9950 19796 9956 19808
rect 10008 19796 10014 19848
rect 10336 19845 10364 19876
rect 12526 19864 12532 19876
rect 12584 19864 12590 19916
rect 12710 19864 12716 19916
rect 12768 19904 12774 19916
rect 13265 19907 13323 19913
rect 13265 19904 13277 19907
rect 12768 19876 13277 19904
rect 12768 19864 12774 19876
rect 13265 19873 13277 19876
rect 13311 19873 13323 19907
rect 13265 19867 13323 19873
rect 10321 19839 10379 19845
rect 10321 19805 10333 19839
rect 10367 19805 10379 19839
rect 10321 19799 10379 19805
rect 10686 19796 10692 19848
rect 10744 19796 10750 19848
rect 12437 19839 12495 19845
rect 12437 19805 12449 19839
rect 12483 19836 12495 19839
rect 12618 19836 12624 19848
rect 12483 19808 12624 19836
rect 12483 19805 12495 19808
rect 12437 19799 12495 19805
rect 12618 19796 12624 19808
rect 12676 19796 12682 19848
rect 12805 19839 12863 19845
rect 12805 19805 12817 19839
rect 12851 19836 12863 19839
rect 12894 19836 12900 19848
rect 12851 19808 12900 19836
rect 12851 19805 12863 19808
rect 12805 19799 12863 19805
rect 12894 19796 12900 19808
rect 12952 19796 12958 19848
rect 12986 19796 12992 19848
rect 13044 19796 13050 19848
rect 14108 19845 14136 19944
rect 14200 19876 14504 19904
rect 14200 19845 14228 19876
rect 14093 19839 14151 19845
rect 14093 19805 14105 19839
rect 14139 19805 14151 19839
rect 14093 19799 14151 19805
rect 14185 19839 14243 19845
rect 14185 19805 14197 19839
rect 14231 19805 14243 19839
rect 14185 19799 14243 19805
rect 14476 19780 14504 19876
rect 14599 19839 14657 19845
rect 14599 19805 14611 19839
rect 14645 19836 14657 19839
rect 14752 19836 14780 19944
rect 15028 19944 15476 19972
rect 15028 19904 15056 19944
rect 15470 19932 15476 19944
rect 15528 19932 15534 19984
rect 17034 19932 17040 19984
rect 17092 19972 17098 19984
rect 20272 19972 20300 20012
rect 21174 19972 21180 19984
rect 17092 19944 20300 19972
rect 21008 19944 21180 19972
rect 17092 19932 17098 19944
rect 19702 19904 19708 19916
rect 14844 19876 15056 19904
rect 15488 19876 19708 19904
rect 14844 19845 14872 19876
rect 14645 19808 14780 19836
rect 14829 19839 14887 19845
rect 14645 19805 14657 19808
rect 14599 19799 14657 19805
rect 14829 19805 14841 19839
rect 14875 19805 14887 19839
rect 14829 19799 14887 19805
rect 14918 19796 14924 19848
rect 14976 19845 14982 19848
rect 14976 19839 15015 19845
rect 15003 19805 15015 19839
rect 14976 19799 15015 19805
rect 15105 19839 15163 19845
rect 15105 19805 15117 19839
rect 15151 19836 15163 19839
rect 15286 19836 15292 19848
rect 15151 19808 15292 19836
rect 15151 19805 15163 19808
rect 15105 19799 15163 19805
rect 14976 19796 14982 19799
rect 15286 19796 15292 19808
rect 15344 19796 15350 19848
rect 15378 19796 15384 19848
rect 15436 19796 15442 19848
rect 15488 19845 15516 19876
rect 19702 19864 19708 19876
rect 19760 19864 19766 19916
rect 21008 19913 21036 19944
rect 21174 19932 21180 19944
rect 21232 19932 21238 19984
rect 21266 19932 21272 19984
rect 21324 19932 21330 19984
rect 21358 19932 21364 19984
rect 21416 19932 21422 19984
rect 21652 19981 21680 20012
rect 22830 20000 22836 20052
rect 22888 20000 22894 20052
rect 23106 20000 23112 20052
rect 23164 20040 23170 20052
rect 25041 20043 25099 20049
rect 23164 20012 24440 20040
rect 23164 20000 23170 20012
rect 21637 19975 21695 19981
rect 21637 19941 21649 19975
rect 21683 19941 21695 19975
rect 21637 19935 21695 19941
rect 22094 19932 22100 19984
rect 22152 19972 22158 19984
rect 23198 19972 23204 19984
rect 22152 19944 23204 19972
rect 22152 19932 22158 19944
rect 23198 19932 23204 19944
rect 23256 19932 23262 19984
rect 24412 19972 24440 20012
rect 25041 20009 25053 20043
rect 25087 20040 25099 20043
rect 25130 20040 25136 20052
rect 25087 20012 25136 20040
rect 25087 20009 25099 20012
rect 25041 20003 25099 20009
rect 25130 20000 25136 20012
rect 25188 20000 25194 20052
rect 25314 20000 25320 20052
rect 25372 20000 25378 20052
rect 25406 20000 25412 20052
rect 25464 20040 25470 20052
rect 25501 20043 25559 20049
rect 25501 20040 25513 20043
rect 25464 20012 25513 20040
rect 25464 20000 25470 20012
rect 25501 20009 25513 20012
rect 25547 20009 25559 20043
rect 25501 20003 25559 20009
rect 26050 20000 26056 20052
rect 26108 20000 26114 20052
rect 26513 20043 26571 20049
rect 26513 20009 26525 20043
rect 26559 20040 26571 20043
rect 26694 20040 26700 20052
rect 26559 20012 26700 20040
rect 26559 20009 26571 20012
rect 26513 20003 26571 20009
rect 26694 20000 26700 20012
rect 26752 20000 26758 20052
rect 27706 20000 27712 20052
rect 27764 20040 27770 20052
rect 27893 20043 27951 20049
rect 27893 20040 27905 20043
rect 27764 20012 27905 20040
rect 27764 20000 27770 20012
rect 27893 20009 27905 20012
rect 27939 20009 27951 20043
rect 27893 20003 27951 20009
rect 25774 19972 25780 19984
rect 24412 19944 25780 19972
rect 20993 19907 21051 19913
rect 20993 19873 21005 19907
rect 21039 19873 21051 19907
rect 20993 19867 21051 19873
rect 21085 19907 21143 19913
rect 21085 19873 21097 19907
rect 21131 19904 21143 19907
rect 22830 19904 22836 19916
rect 21131 19876 22836 19904
rect 21131 19873 21143 19876
rect 21085 19867 21143 19873
rect 22830 19864 22836 19876
rect 22888 19864 22894 19916
rect 23293 19907 23351 19913
rect 23293 19873 23305 19907
rect 23339 19904 23351 19907
rect 23382 19904 23388 19916
rect 23339 19876 23388 19904
rect 23339 19873 23351 19876
rect 23293 19867 23351 19873
rect 23382 19864 23388 19876
rect 23440 19864 23446 19916
rect 15473 19839 15531 19845
rect 15473 19805 15485 19839
rect 15519 19805 15531 19839
rect 15473 19799 15531 19805
rect 7699 19740 8376 19768
rect 7699 19737 7711 19740
rect 7653 19731 7711 19737
rect 10410 19728 10416 19780
rect 10468 19728 10474 19780
rect 10505 19771 10563 19777
rect 10505 19737 10517 19771
rect 10551 19737 10563 19771
rect 10505 19731 10563 19737
rect 13725 19771 13783 19777
rect 13725 19737 13737 19771
rect 13771 19768 13783 19771
rect 13814 19768 13820 19780
rect 13771 19740 13820 19768
rect 13771 19737 13783 19740
rect 13725 19731 13783 19737
rect 5316 19672 5856 19700
rect 5316 19660 5322 19672
rect 7190 19660 7196 19712
rect 7248 19660 7254 19712
rect 8110 19660 8116 19712
rect 8168 19660 8174 19712
rect 10042 19660 10048 19712
rect 10100 19700 10106 19712
rect 10520 19700 10548 19731
rect 13814 19728 13820 19740
rect 13872 19728 13878 19780
rect 13921 19771 13979 19777
rect 13921 19737 13933 19771
rect 13967 19768 13979 19771
rect 13967 19740 14090 19768
rect 13967 19737 13979 19740
rect 13921 19731 13979 19737
rect 13538 19700 13544 19712
rect 10100 19672 13544 19700
rect 10100 19660 10106 19672
rect 13538 19660 13544 19672
rect 13596 19660 13602 19712
rect 14062 19700 14090 19740
rect 14366 19728 14372 19780
rect 14424 19728 14430 19780
rect 14458 19728 14464 19780
rect 14516 19768 14522 19780
rect 14737 19771 14795 19777
rect 14737 19768 14749 19771
rect 14516 19740 14749 19768
rect 14516 19728 14522 19740
rect 14737 19737 14749 19740
rect 14783 19768 14795 19771
rect 15488 19768 15516 19799
rect 15654 19796 15660 19848
rect 15712 19796 15718 19848
rect 15749 19839 15807 19845
rect 15749 19805 15761 19839
rect 15795 19805 15807 19839
rect 15749 19799 15807 19805
rect 14783 19740 15516 19768
rect 14783 19737 14795 19740
rect 14737 19731 14795 19737
rect 14274 19700 14280 19712
rect 14062 19672 14280 19700
rect 14274 19660 14280 19672
rect 14332 19660 14338 19712
rect 15010 19660 15016 19712
rect 15068 19700 15074 19712
rect 15197 19703 15255 19709
rect 15197 19700 15209 19703
rect 15068 19672 15209 19700
rect 15068 19660 15074 19672
rect 15197 19669 15209 19672
rect 15243 19669 15255 19703
rect 15197 19663 15255 19669
rect 15286 19660 15292 19712
rect 15344 19700 15350 19712
rect 15764 19700 15792 19799
rect 18690 19796 18696 19848
rect 18748 19836 18754 19848
rect 19518 19836 19524 19848
rect 18748 19808 19524 19836
rect 18748 19796 18754 19808
rect 19518 19796 19524 19808
rect 19576 19796 19582 19848
rect 20070 19796 20076 19848
rect 20128 19836 20134 19848
rect 20257 19839 20315 19845
rect 20257 19836 20269 19839
rect 20128 19808 20269 19836
rect 20128 19796 20134 19808
rect 20257 19805 20269 19808
rect 20303 19805 20315 19839
rect 20257 19799 20315 19805
rect 20349 19839 20407 19845
rect 20349 19805 20361 19839
rect 20395 19805 20407 19839
rect 20349 19799 20407 19805
rect 17586 19728 17592 19780
rect 17644 19768 17650 19780
rect 19334 19768 19340 19780
rect 17644 19740 19340 19768
rect 17644 19728 17650 19740
rect 19334 19728 19340 19740
rect 19392 19768 19398 19780
rect 19610 19768 19616 19780
rect 19392 19740 19616 19768
rect 19392 19728 19398 19740
rect 19610 19728 19616 19740
rect 19668 19728 19674 19780
rect 20364 19768 20392 19799
rect 20530 19796 20536 19848
rect 20588 19796 20594 19848
rect 20622 19796 20628 19848
rect 20680 19796 20686 19848
rect 20806 19796 20812 19848
rect 20864 19796 20870 19848
rect 20901 19839 20959 19845
rect 20901 19805 20913 19839
rect 20947 19805 20959 19839
rect 20901 19799 20959 19805
rect 20916 19768 20944 19799
rect 21266 19796 21272 19848
rect 21324 19836 21330 19848
rect 21545 19839 21603 19845
rect 21545 19836 21557 19839
rect 21324 19808 21557 19836
rect 21324 19796 21330 19808
rect 21545 19805 21557 19808
rect 21591 19805 21603 19839
rect 21545 19799 21603 19805
rect 21726 19796 21732 19848
rect 21784 19796 21790 19848
rect 21818 19796 21824 19848
rect 21876 19796 21882 19848
rect 22278 19836 22284 19848
rect 21928 19808 22284 19836
rect 21928 19768 21956 19808
rect 22278 19796 22284 19808
rect 22336 19796 22342 19848
rect 22738 19796 22744 19848
rect 22796 19836 22802 19848
rect 23017 19839 23075 19845
rect 23017 19836 23029 19839
rect 22796 19808 23029 19836
rect 22796 19796 22802 19808
rect 23017 19805 23029 19808
rect 23063 19836 23075 19839
rect 23106 19836 23112 19848
rect 23063 19808 23112 19836
rect 23063 19805 23075 19808
rect 23017 19799 23075 19805
rect 23106 19796 23112 19808
rect 23164 19796 23170 19848
rect 23566 19796 23572 19848
rect 23624 19836 23630 19848
rect 24412 19845 24440 19944
rect 25774 19932 25780 19944
rect 25832 19972 25838 19984
rect 26234 19972 26240 19984
rect 25832 19944 26240 19972
rect 25832 19932 25838 19944
rect 26234 19932 26240 19944
rect 26292 19932 26298 19984
rect 27801 19975 27859 19981
rect 27801 19941 27813 19975
rect 27847 19972 27859 19975
rect 28258 19972 28264 19984
rect 27847 19944 28264 19972
rect 27847 19941 27859 19944
rect 27801 19935 27859 19941
rect 28258 19932 28264 19944
rect 28316 19932 28322 19984
rect 29089 19975 29147 19981
rect 29089 19941 29101 19975
rect 29135 19972 29147 19975
rect 29914 19972 29920 19984
rect 29135 19944 29920 19972
rect 29135 19941 29147 19944
rect 29089 19935 29147 19941
rect 29914 19932 29920 19944
rect 29972 19932 29978 19984
rect 30098 19932 30104 19984
rect 30156 19932 30162 19984
rect 33686 19932 33692 19984
rect 33744 19972 33750 19984
rect 34422 19972 34428 19984
rect 33744 19944 34428 19972
rect 33744 19932 33750 19944
rect 34422 19932 34428 19944
rect 34480 19972 34486 19984
rect 34480 19944 39344 19972
rect 34480 19932 34486 19944
rect 24688 19876 24992 19904
rect 23753 19839 23811 19845
rect 23753 19836 23765 19839
rect 23624 19808 23765 19836
rect 23624 19796 23630 19808
rect 23753 19805 23765 19808
rect 23799 19805 23811 19839
rect 23753 19799 23811 19805
rect 24397 19839 24455 19845
rect 24397 19805 24409 19839
rect 24443 19805 24455 19839
rect 24397 19799 24455 19805
rect 24486 19796 24492 19848
rect 24544 19833 24550 19848
rect 24688 19845 24716 19876
rect 24581 19839 24639 19845
rect 24581 19833 24593 19839
rect 24544 19805 24593 19833
rect 24627 19805 24639 19839
rect 24544 19796 24550 19805
rect 24581 19799 24639 19805
rect 24673 19839 24731 19845
rect 24673 19805 24685 19839
rect 24719 19805 24731 19839
rect 24673 19799 24731 19805
rect 24765 19839 24823 19845
rect 24765 19805 24777 19839
rect 24811 19805 24823 19839
rect 24964 19836 24992 19876
rect 25038 19864 25044 19916
rect 25096 19904 25102 19916
rect 26421 19907 26479 19913
rect 25096 19876 25912 19904
rect 25096 19864 25102 19876
rect 24964 19808 25392 19836
rect 24765 19799 24823 19805
rect 20364 19740 21956 19768
rect 22186 19728 22192 19780
rect 22244 19768 22250 19780
rect 24512 19768 24540 19796
rect 24780 19768 24808 19799
rect 22244 19740 24540 19768
rect 24596 19740 24808 19768
rect 22244 19728 22250 19740
rect 24596 19712 24624 19740
rect 25130 19728 25136 19780
rect 25188 19728 25194 19780
rect 25364 19777 25392 19808
rect 25349 19771 25407 19777
rect 25349 19737 25361 19771
rect 25395 19768 25407 19771
rect 25498 19768 25504 19780
rect 25395 19740 25504 19768
rect 25395 19737 25407 19740
rect 25349 19731 25407 19737
rect 25498 19728 25504 19740
rect 25556 19728 25562 19780
rect 15344 19672 15792 19700
rect 15344 19660 15350 19672
rect 17402 19660 17408 19712
rect 17460 19700 17466 19712
rect 18874 19700 18880 19712
rect 17460 19672 18880 19700
rect 17460 19660 17466 19672
rect 18874 19660 18880 19672
rect 18932 19660 18938 19712
rect 22370 19660 22376 19712
rect 22428 19700 22434 19712
rect 23474 19700 23480 19712
rect 22428 19672 23480 19700
rect 22428 19660 22434 19672
rect 23474 19660 23480 19672
rect 23532 19700 23538 19712
rect 23569 19703 23627 19709
rect 23569 19700 23581 19703
rect 23532 19672 23581 19700
rect 23532 19660 23538 19672
rect 23569 19669 23581 19672
rect 23615 19669 23627 19703
rect 23569 19663 23627 19669
rect 23750 19660 23756 19712
rect 23808 19700 23814 19712
rect 24302 19700 24308 19712
rect 23808 19672 24308 19700
rect 23808 19660 23814 19672
rect 24302 19660 24308 19672
rect 24360 19660 24366 19712
rect 24578 19660 24584 19712
rect 24636 19660 24642 19712
rect 25884 19700 25912 19876
rect 26421 19873 26433 19907
rect 26467 19904 26479 19907
rect 28442 19904 28448 19916
rect 26467 19876 28448 19904
rect 26467 19873 26479 19876
rect 26421 19867 26479 19873
rect 28442 19864 28448 19876
rect 28500 19864 28506 19916
rect 29825 19907 29883 19913
rect 29825 19873 29837 19907
rect 29871 19904 29883 19907
rect 30116 19904 30144 19932
rect 31386 19904 31392 19916
rect 29871 19876 30144 19904
rect 31312 19876 31392 19904
rect 29871 19873 29883 19876
rect 29825 19867 29883 19873
rect 26237 19839 26295 19845
rect 26237 19805 26249 19839
rect 26283 19836 26295 19839
rect 26602 19836 26608 19848
rect 26283 19808 26608 19836
rect 26283 19805 26295 19808
rect 26237 19799 26295 19805
rect 26602 19796 26608 19808
rect 26660 19796 26666 19848
rect 27246 19796 27252 19848
rect 27304 19836 27310 19848
rect 27341 19839 27399 19845
rect 27341 19836 27353 19839
rect 27304 19808 27353 19836
rect 27304 19796 27310 19808
rect 27341 19805 27353 19808
rect 27387 19836 27399 19839
rect 27522 19836 27528 19848
rect 27387 19808 27528 19836
rect 27387 19805 27399 19808
rect 27341 19799 27399 19805
rect 27522 19796 27528 19808
rect 27580 19796 27586 19848
rect 27617 19839 27675 19845
rect 27617 19805 27629 19839
rect 27663 19805 27675 19839
rect 27617 19799 27675 19805
rect 26510 19728 26516 19780
rect 26568 19728 26574 19780
rect 27154 19728 27160 19780
rect 27212 19768 27218 19780
rect 27632 19768 27660 19799
rect 27890 19796 27896 19848
rect 27948 19836 27954 19848
rect 28261 19839 28319 19845
rect 28261 19836 28273 19839
rect 27948 19808 28273 19836
rect 27948 19796 27954 19808
rect 28261 19805 28273 19808
rect 28307 19805 28319 19839
rect 28261 19799 28319 19805
rect 28902 19796 28908 19848
rect 28960 19836 28966 19848
rect 29273 19839 29331 19845
rect 29273 19836 29285 19839
rect 28960 19808 29285 19836
rect 28960 19796 28966 19808
rect 29273 19805 29285 19808
rect 29319 19836 29331 19839
rect 30101 19839 30159 19845
rect 30101 19836 30113 19839
rect 29319 19808 30113 19836
rect 29319 19805 29331 19808
rect 29273 19799 29331 19805
rect 30101 19805 30113 19808
rect 30147 19805 30159 19839
rect 30101 19799 30159 19805
rect 31113 19839 31171 19845
rect 31113 19805 31125 19839
rect 31159 19836 31171 19839
rect 31202 19836 31208 19848
rect 31159 19808 31208 19836
rect 31159 19805 31171 19808
rect 31113 19799 31171 19805
rect 31202 19796 31208 19808
rect 31260 19796 31266 19848
rect 31312 19845 31340 19876
rect 31386 19864 31392 19876
rect 31444 19864 31450 19916
rect 33870 19864 33876 19916
rect 33928 19904 33934 19916
rect 35158 19904 35164 19916
rect 33928 19876 35164 19904
rect 33928 19864 33934 19876
rect 35158 19864 35164 19876
rect 35216 19864 35222 19916
rect 35342 19864 35348 19916
rect 35400 19904 35406 19916
rect 37918 19904 37924 19916
rect 35400 19876 37924 19904
rect 35400 19864 35406 19876
rect 37918 19864 37924 19876
rect 37976 19904 37982 19916
rect 39316 19913 39344 19944
rect 38933 19907 38991 19913
rect 38933 19904 38945 19907
rect 37976 19876 38945 19904
rect 37976 19864 37982 19876
rect 38933 19873 38945 19876
rect 38979 19873 38991 19907
rect 38933 19867 38991 19873
rect 39301 19907 39359 19913
rect 39301 19873 39313 19907
rect 39347 19873 39359 19907
rect 39301 19867 39359 19873
rect 31297 19839 31355 19845
rect 31297 19805 31309 19839
rect 31343 19805 31355 19839
rect 31297 19799 31355 19805
rect 31478 19796 31484 19848
rect 31536 19836 31542 19848
rect 31662 19836 31668 19848
rect 31536 19808 31668 19836
rect 31536 19796 31542 19808
rect 31662 19796 31668 19808
rect 31720 19796 31726 19848
rect 33042 19796 33048 19848
rect 33100 19836 33106 19848
rect 36446 19836 36452 19848
rect 33100 19808 36452 19836
rect 33100 19796 33106 19808
rect 36446 19796 36452 19808
rect 36504 19836 36510 19848
rect 36817 19839 36875 19845
rect 36817 19836 36829 19839
rect 36504 19808 36829 19836
rect 36504 19796 36510 19808
rect 36817 19805 36829 19808
rect 36863 19805 36875 19839
rect 36817 19799 36875 19805
rect 36906 19796 36912 19848
rect 36964 19796 36970 19848
rect 37274 19796 37280 19848
rect 37332 19845 37338 19848
rect 37332 19836 37340 19845
rect 38010 19836 38016 19848
rect 37332 19808 38016 19836
rect 37332 19799 37340 19808
rect 37332 19796 37338 19799
rect 38010 19796 38016 19808
rect 38068 19796 38074 19848
rect 38841 19839 38899 19845
rect 38841 19805 38853 19839
rect 38887 19805 38899 19839
rect 38841 19799 38899 19805
rect 39117 19839 39175 19845
rect 39117 19805 39129 19839
rect 39163 19836 39175 19839
rect 39206 19836 39212 19848
rect 39163 19808 39212 19836
rect 39163 19805 39175 19808
rect 39117 19799 39175 19805
rect 27212 19740 27660 19768
rect 27212 19728 27218 19740
rect 27706 19728 27712 19780
rect 27764 19768 27770 19780
rect 27982 19768 27988 19780
rect 27764 19740 27988 19768
rect 27764 19728 27770 19740
rect 27982 19728 27988 19740
rect 28040 19768 28046 19780
rect 28077 19771 28135 19777
rect 28077 19768 28089 19771
rect 28040 19740 28089 19768
rect 28040 19728 28046 19740
rect 28077 19737 28089 19740
rect 28123 19737 28135 19771
rect 28077 19731 28135 19737
rect 30466 19728 30472 19780
rect 30524 19768 30530 19780
rect 31389 19771 31447 19777
rect 31389 19768 31401 19771
rect 30524 19740 31401 19768
rect 30524 19728 30530 19740
rect 31389 19737 31401 19740
rect 31435 19737 31447 19771
rect 31389 19731 31447 19737
rect 33318 19728 33324 19780
rect 33376 19768 33382 19780
rect 36170 19768 36176 19780
rect 33376 19740 36176 19768
rect 33376 19728 33382 19740
rect 36170 19728 36176 19740
rect 36228 19728 36234 19780
rect 36354 19728 36360 19780
rect 36412 19768 36418 19780
rect 37093 19771 37151 19777
rect 37093 19768 37105 19771
rect 36412 19740 37105 19768
rect 36412 19728 36418 19740
rect 37093 19737 37105 19740
rect 37139 19737 37151 19771
rect 37093 19731 37151 19737
rect 37182 19728 37188 19780
rect 37240 19728 37246 19780
rect 38102 19768 38108 19780
rect 37384 19740 38108 19768
rect 37384 19712 37412 19740
rect 38102 19728 38108 19740
rect 38160 19768 38166 19780
rect 38565 19771 38623 19777
rect 38565 19768 38577 19771
rect 38160 19740 38577 19768
rect 38160 19728 38166 19740
rect 38565 19737 38577 19740
rect 38611 19737 38623 19771
rect 38856 19768 38884 19799
rect 39206 19796 39212 19808
rect 39264 19796 39270 19848
rect 39666 19768 39672 19780
rect 38856 19740 39672 19768
rect 38565 19731 38623 19737
rect 39666 19728 39672 19740
rect 39724 19728 39730 19780
rect 27433 19703 27491 19709
rect 27433 19700 27445 19703
rect 25884 19672 27445 19700
rect 27433 19669 27445 19672
rect 27479 19669 27491 19703
rect 27433 19663 27491 19669
rect 28718 19660 28724 19712
rect 28776 19700 28782 19712
rect 31570 19700 31576 19712
rect 28776 19672 31576 19700
rect 28776 19660 28782 19672
rect 31570 19660 31576 19672
rect 31628 19660 31634 19712
rect 31665 19703 31723 19709
rect 31665 19669 31677 19703
rect 31711 19700 31723 19703
rect 32398 19700 32404 19712
rect 31711 19672 32404 19700
rect 31711 19669 31723 19672
rect 31665 19663 31723 19669
rect 32398 19660 32404 19672
rect 32456 19660 32462 19712
rect 33686 19660 33692 19712
rect 33744 19700 33750 19712
rect 33870 19700 33876 19712
rect 33744 19672 33876 19700
rect 33744 19660 33750 19672
rect 33870 19660 33876 19672
rect 33928 19660 33934 19712
rect 37366 19660 37372 19712
rect 37424 19660 37430 19712
rect 37458 19660 37464 19712
rect 37516 19660 37522 19712
rect 1104 19610 40572 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 40572 19610
rect 1104 19536 40572 19558
rect 3418 19456 3424 19508
rect 3476 19456 3482 19508
rect 3878 19456 3884 19508
rect 3936 19456 3942 19508
rect 4798 19456 4804 19508
rect 4856 19496 4862 19508
rect 5166 19496 5172 19508
rect 4856 19468 5172 19496
rect 4856 19456 4862 19468
rect 5166 19456 5172 19468
rect 5224 19496 5230 19508
rect 6822 19496 6828 19508
rect 5224 19468 6828 19496
rect 5224 19456 5230 19468
rect 6822 19456 6828 19468
rect 6880 19496 6886 19508
rect 8570 19496 8576 19508
rect 6880 19468 8576 19496
rect 6880 19456 6886 19468
rect 3510 19388 3516 19440
rect 3568 19428 3574 19440
rect 3973 19431 4031 19437
rect 3973 19428 3985 19431
rect 3568 19400 3985 19428
rect 3568 19388 3574 19400
rect 3973 19397 3985 19400
rect 4019 19428 4031 19431
rect 5718 19428 5724 19440
rect 4019 19400 5724 19428
rect 4019 19397 4031 19400
rect 3973 19391 4031 19397
rect 5718 19388 5724 19400
rect 5776 19388 5782 19440
rect 6733 19431 6791 19437
rect 6733 19428 6745 19431
rect 5828 19400 6745 19428
rect 3050 19320 3056 19372
rect 3108 19320 3114 19372
rect 5534 19320 5540 19372
rect 5592 19360 5598 19372
rect 5828 19369 5856 19400
rect 6733 19397 6745 19400
rect 6779 19397 6791 19431
rect 6733 19391 6791 19397
rect 5813 19363 5871 19369
rect 5813 19360 5825 19363
rect 5592 19332 5825 19360
rect 5592 19320 5598 19332
rect 5813 19329 5825 19332
rect 5859 19329 5871 19363
rect 6549 19363 6607 19369
rect 6549 19360 6561 19363
rect 6527 19332 6561 19360
rect 5813 19323 5871 19329
rect 6549 19329 6561 19332
rect 6595 19329 6607 19363
rect 6549 19323 6607 19329
rect 1578 19252 1584 19304
rect 1636 19292 1642 19304
rect 1673 19295 1731 19301
rect 1673 19292 1685 19295
rect 1636 19264 1685 19292
rect 1636 19252 1642 19264
rect 1673 19261 1685 19264
rect 1719 19261 1731 19295
rect 1673 19255 1731 19261
rect 1949 19295 2007 19301
rect 1949 19261 1961 19295
rect 1995 19292 2007 19295
rect 1995 19264 3556 19292
rect 1995 19261 2007 19264
rect 1949 19255 2007 19261
rect 3528 19233 3556 19264
rect 4062 19252 4068 19304
rect 4120 19252 4126 19304
rect 4614 19252 4620 19304
rect 4672 19252 4678 19304
rect 4890 19252 4896 19304
rect 4948 19292 4954 19304
rect 5442 19292 5448 19304
rect 4948 19264 5448 19292
rect 4948 19252 4954 19264
rect 5442 19252 5448 19264
rect 5500 19252 5506 19304
rect 5902 19252 5908 19304
rect 5960 19292 5966 19304
rect 6365 19295 6423 19301
rect 6365 19292 6377 19295
rect 5960 19264 6377 19292
rect 5960 19252 5966 19264
rect 6365 19261 6377 19264
rect 6411 19261 6423 19295
rect 6564 19292 6592 19323
rect 6638 19320 6644 19372
rect 6696 19360 6702 19372
rect 6932 19369 6960 19468
rect 8570 19456 8576 19468
rect 8628 19456 8634 19508
rect 8662 19456 8668 19508
rect 8720 19456 8726 19508
rect 10410 19456 10416 19508
rect 10468 19496 10474 19508
rect 10505 19499 10563 19505
rect 10505 19496 10517 19499
rect 10468 19468 10517 19496
rect 10468 19456 10474 19468
rect 10505 19465 10517 19468
rect 10551 19465 10563 19499
rect 10505 19459 10563 19465
rect 7466 19388 7472 19440
rect 7524 19428 7530 19440
rect 9490 19428 9496 19440
rect 7524 19400 7682 19428
rect 8418 19400 9496 19428
rect 7524 19388 7530 19400
rect 9490 19388 9496 19400
rect 9548 19388 9554 19440
rect 6825 19363 6883 19369
rect 6825 19360 6837 19363
rect 6696 19332 6837 19360
rect 6696 19320 6702 19332
rect 6825 19329 6837 19332
rect 6871 19329 6883 19363
rect 6825 19323 6883 19329
rect 6917 19363 6975 19369
rect 6917 19329 6929 19363
rect 6963 19329 6975 19363
rect 6917 19323 6975 19329
rect 8570 19320 8576 19372
rect 8628 19360 8634 19372
rect 8757 19363 8815 19369
rect 8757 19360 8769 19363
rect 8628 19332 8769 19360
rect 8628 19320 8634 19332
rect 8757 19329 8769 19332
rect 8803 19329 8815 19363
rect 10520 19360 10548 19459
rect 12526 19456 12532 19508
rect 12584 19496 12590 19508
rect 13725 19499 13783 19505
rect 13725 19496 13737 19499
rect 12584 19468 13737 19496
rect 12584 19456 12590 19468
rect 13725 19465 13737 19468
rect 13771 19465 13783 19499
rect 13725 19459 13783 19465
rect 14274 19456 14280 19508
rect 14332 19456 14338 19508
rect 15010 19496 15016 19508
rect 14384 19468 15016 19496
rect 14384 19428 14412 19468
rect 15010 19456 15016 19468
rect 15068 19456 15074 19508
rect 15197 19499 15255 19505
rect 15197 19465 15209 19499
rect 15243 19496 15255 19499
rect 15286 19496 15292 19508
rect 15243 19468 15292 19496
rect 15243 19465 15255 19468
rect 15197 19459 15255 19465
rect 15212 19428 15240 19459
rect 15286 19456 15292 19468
rect 15344 19456 15350 19508
rect 15562 19456 15568 19508
rect 15620 19496 15626 19508
rect 15657 19499 15715 19505
rect 15657 19496 15669 19499
rect 15620 19468 15669 19496
rect 15620 19456 15626 19468
rect 15657 19465 15669 19468
rect 15703 19465 15715 19499
rect 15657 19459 15715 19465
rect 17126 19456 17132 19508
rect 17184 19456 17190 19508
rect 17221 19499 17279 19505
rect 17221 19465 17233 19499
rect 17267 19496 17279 19499
rect 17402 19496 17408 19508
rect 17267 19468 17408 19496
rect 17267 19465 17279 19468
rect 17221 19459 17279 19465
rect 17402 19456 17408 19468
rect 17460 19456 17466 19508
rect 18417 19499 18475 19505
rect 18417 19496 18429 19499
rect 17696 19468 18429 19496
rect 13832 19400 14412 19428
rect 14476 19400 15240 19428
rect 13832 19369 13860 19400
rect 13817 19363 13875 19369
rect 10520 19332 11192 19360
rect 8757 19323 8815 19329
rect 6730 19292 6736 19304
rect 6564 19264 6736 19292
rect 6365 19255 6423 19261
rect 6730 19252 6736 19264
rect 6788 19252 6794 19304
rect 7193 19295 7251 19301
rect 7193 19261 7205 19295
rect 7239 19292 7251 19295
rect 7650 19292 7656 19304
rect 7239 19264 7656 19292
rect 7239 19261 7251 19264
rect 7193 19255 7251 19261
rect 7650 19252 7656 19264
rect 7708 19252 7714 19304
rect 9033 19295 9091 19301
rect 9033 19261 9045 19295
rect 9079 19292 9091 19295
rect 9490 19292 9496 19304
rect 9079 19264 9496 19292
rect 9079 19261 9091 19264
rect 9033 19255 9091 19261
rect 9490 19252 9496 19264
rect 9548 19252 9554 19304
rect 11164 19301 11192 19332
rect 13817 19329 13829 19363
rect 13863 19329 13875 19363
rect 13817 19323 13875 19329
rect 14001 19363 14059 19369
rect 14001 19329 14013 19363
rect 14047 19360 14059 19363
rect 14090 19360 14096 19372
rect 14047 19332 14096 19360
rect 14047 19329 14059 19332
rect 14001 19323 14059 19329
rect 14090 19320 14096 19332
rect 14148 19320 14154 19372
rect 14366 19320 14372 19372
rect 14424 19320 14430 19372
rect 14476 19369 14504 19400
rect 15746 19388 15752 19440
rect 15804 19428 15810 19440
rect 17696 19437 17724 19468
rect 18417 19465 18429 19468
rect 18463 19496 18475 19499
rect 18463 19468 19012 19496
rect 18463 19465 18475 19468
rect 18417 19459 18475 19465
rect 17681 19431 17739 19437
rect 15804 19400 17448 19428
rect 15804 19388 15810 19400
rect 14461 19363 14519 19369
rect 14461 19329 14473 19363
rect 14507 19329 14519 19363
rect 14645 19363 14703 19369
rect 14645 19360 14657 19363
rect 14461 19323 14519 19329
rect 14568 19332 14657 19360
rect 11149 19295 11207 19301
rect 11149 19261 11161 19295
rect 11195 19261 11207 19295
rect 14384 19292 14412 19320
rect 14568 19292 14596 19332
rect 14645 19329 14657 19332
rect 14691 19329 14703 19363
rect 14645 19323 14703 19329
rect 14737 19363 14795 19369
rect 14737 19329 14749 19363
rect 14783 19360 14795 19363
rect 15286 19360 15292 19372
rect 14783 19332 15292 19360
rect 14783 19329 14795 19332
rect 14737 19323 14795 19329
rect 15286 19320 15292 19332
rect 15344 19320 15350 19372
rect 15381 19363 15439 19369
rect 15381 19329 15393 19363
rect 15427 19360 15439 19363
rect 15838 19360 15844 19372
rect 15427 19332 15844 19360
rect 15427 19329 15439 19332
rect 15381 19323 15439 19329
rect 15838 19320 15844 19332
rect 15896 19360 15902 19372
rect 15933 19363 15991 19369
rect 15933 19360 15945 19363
rect 15896 19332 15945 19360
rect 15896 19320 15902 19332
rect 15933 19329 15945 19332
rect 15979 19329 15991 19363
rect 15933 19323 15991 19329
rect 16206 19320 16212 19372
rect 16264 19320 16270 19372
rect 16390 19320 16396 19372
rect 16448 19320 16454 19372
rect 17420 19369 17448 19400
rect 17681 19397 17693 19431
rect 17727 19397 17739 19431
rect 17681 19391 17739 19397
rect 17957 19431 18015 19437
rect 17957 19397 17969 19431
rect 18003 19428 18015 19431
rect 18046 19428 18052 19440
rect 18003 19400 18052 19428
rect 18003 19397 18015 19400
rect 17957 19391 18015 19397
rect 18046 19388 18052 19400
rect 18104 19388 18110 19440
rect 18233 19431 18291 19437
rect 18233 19397 18245 19431
rect 18279 19428 18291 19431
rect 18690 19428 18696 19440
rect 18279 19400 18696 19428
rect 18279 19397 18291 19400
rect 18233 19391 18291 19397
rect 18690 19388 18696 19400
rect 18748 19388 18754 19440
rect 17586 19369 17592 19372
rect 17037 19363 17095 19369
rect 17037 19329 17049 19363
rect 17083 19329 17095 19363
rect 17037 19323 17095 19329
rect 17405 19363 17463 19369
rect 17405 19329 17417 19363
rect 17451 19329 17463 19363
rect 17584 19360 17592 19369
rect 17547 19332 17592 19360
rect 17405 19323 17463 19329
rect 17584 19323 17592 19332
rect 14384 19264 14596 19292
rect 15565 19295 15623 19301
rect 11149 19255 11207 19261
rect 15565 19261 15577 19295
rect 15611 19292 15623 19295
rect 15657 19295 15715 19301
rect 15657 19292 15669 19295
rect 15611 19264 15669 19292
rect 15611 19261 15623 19264
rect 15565 19255 15623 19261
rect 15657 19261 15669 19264
rect 15703 19292 15715 19295
rect 16758 19292 16764 19304
rect 15703 19264 16764 19292
rect 15703 19261 15715 19264
rect 15657 19255 15715 19261
rect 16758 19252 16764 19264
rect 16816 19252 16822 19304
rect 17052 19292 17080 19323
rect 17586 19320 17592 19323
rect 17644 19320 17650 19372
rect 17770 19320 17776 19372
rect 17828 19320 17834 19372
rect 18322 19320 18328 19372
rect 18380 19320 18386 19372
rect 18506 19320 18512 19372
rect 18564 19320 18570 19372
rect 18984 19360 19012 19468
rect 20806 19456 20812 19508
rect 20864 19496 20870 19508
rect 21358 19496 21364 19508
rect 20864 19468 21364 19496
rect 20864 19456 20870 19468
rect 21358 19456 21364 19468
rect 21416 19456 21422 19508
rect 21634 19456 21640 19508
rect 21692 19496 21698 19508
rect 21818 19496 21824 19508
rect 21692 19468 21824 19496
rect 21692 19456 21698 19468
rect 21818 19456 21824 19468
rect 21876 19456 21882 19508
rect 21910 19456 21916 19508
rect 21968 19496 21974 19508
rect 22005 19499 22063 19505
rect 22005 19496 22017 19499
rect 21968 19468 22017 19496
rect 21968 19456 21974 19468
rect 22005 19465 22017 19468
rect 22051 19496 22063 19499
rect 22370 19496 22376 19508
rect 22051 19468 22376 19496
rect 22051 19465 22063 19468
rect 22005 19459 22063 19465
rect 22370 19456 22376 19468
rect 22428 19456 22434 19508
rect 23290 19456 23296 19508
rect 23348 19496 23354 19508
rect 23385 19499 23443 19505
rect 23385 19496 23397 19499
rect 23348 19468 23397 19496
rect 23348 19456 23354 19468
rect 23385 19465 23397 19468
rect 23431 19465 23443 19499
rect 23385 19459 23443 19465
rect 24029 19499 24087 19505
rect 24029 19465 24041 19499
rect 24075 19465 24087 19499
rect 24029 19459 24087 19465
rect 22922 19428 22928 19440
rect 19168 19400 22048 19428
rect 19168 19360 19196 19400
rect 18984 19332 19196 19360
rect 19242 19320 19248 19372
rect 19300 19360 19306 19372
rect 21266 19360 21272 19372
rect 19300 19332 21272 19360
rect 19300 19320 19306 19332
rect 21266 19320 21272 19332
rect 21324 19320 21330 19372
rect 21821 19363 21879 19369
rect 21821 19329 21833 19363
rect 21867 19358 21879 19363
rect 21867 19329 21956 19358
rect 21821 19323 21956 19329
rect 17865 19295 17923 19301
rect 17865 19292 17877 19295
rect 17052 19264 17877 19292
rect 17865 19261 17877 19264
rect 17911 19261 17923 19295
rect 17865 19255 17923 19261
rect 3513 19227 3571 19233
rect 3513 19193 3525 19227
rect 3559 19193 3571 19227
rect 4632 19224 4660 19252
rect 4982 19224 4988 19236
rect 4632 19196 4988 19224
rect 3513 19187 3571 19193
rect 4982 19184 4988 19196
rect 5040 19184 5046 19236
rect 14182 19184 14188 19236
rect 14240 19224 14246 19236
rect 14734 19224 14740 19236
rect 14240 19196 14740 19224
rect 14240 19184 14246 19196
rect 14734 19184 14740 19196
rect 14792 19184 14798 19236
rect 15841 19227 15899 19233
rect 15841 19193 15853 19227
rect 15887 19224 15899 19227
rect 15887 19196 16804 19224
rect 15887 19193 15899 19196
rect 15841 19187 15899 19193
rect 4341 19159 4399 19165
rect 4341 19125 4353 19159
rect 4387 19156 4399 19159
rect 4614 19156 4620 19168
rect 4387 19128 4620 19156
rect 4387 19125 4399 19128
rect 4341 19119 4399 19125
rect 4614 19116 4620 19128
rect 4672 19116 4678 19168
rect 4706 19116 4712 19168
rect 4764 19156 4770 19168
rect 5169 19159 5227 19165
rect 5169 19156 5181 19159
rect 4764 19128 5181 19156
rect 4764 19116 4770 19128
rect 5169 19125 5181 19128
rect 5215 19125 5227 19159
rect 5169 19119 5227 19125
rect 10594 19116 10600 19168
rect 10652 19116 10658 19168
rect 15930 19116 15936 19168
rect 15988 19156 15994 19168
rect 16393 19159 16451 19165
rect 16393 19156 16405 19159
rect 15988 19128 16405 19156
rect 15988 19116 15994 19128
rect 16393 19125 16405 19128
rect 16439 19125 16451 19159
rect 16776 19156 16804 19196
rect 16850 19184 16856 19236
rect 16908 19184 16914 19236
rect 18233 19227 18291 19233
rect 18233 19193 18245 19227
rect 18279 19224 18291 19227
rect 18340 19224 18368 19320
rect 21836 19306 21956 19323
rect 21634 19252 21640 19304
rect 21692 19292 21698 19304
rect 21836 19292 21864 19306
rect 21692 19264 21864 19292
rect 22020 19292 22048 19400
rect 22112 19400 22928 19428
rect 22112 19369 22140 19400
rect 22922 19388 22928 19400
rect 22980 19388 22986 19440
rect 23474 19388 23480 19440
rect 23532 19428 23538 19440
rect 23532 19400 23888 19428
rect 23532 19388 23538 19400
rect 22097 19363 22155 19369
rect 22097 19329 22109 19363
rect 22143 19329 22155 19363
rect 22097 19323 22155 19329
rect 22186 19320 22192 19372
rect 22244 19320 22250 19372
rect 22830 19320 22836 19372
rect 22888 19360 22894 19372
rect 23382 19360 23388 19372
rect 22888 19332 23388 19360
rect 22888 19320 22894 19332
rect 23382 19320 23388 19332
rect 23440 19320 23446 19372
rect 23566 19320 23572 19372
rect 23624 19320 23630 19372
rect 23860 19369 23888 19400
rect 23845 19363 23903 19369
rect 23845 19329 23857 19363
rect 23891 19329 23903 19363
rect 23845 19323 23903 19329
rect 22204 19292 22232 19320
rect 22020 19264 22232 19292
rect 21692 19252 21698 19264
rect 23750 19252 23756 19304
rect 23808 19292 23814 19304
rect 24044 19292 24072 19459
rect 25498 19456 25504 19508
rect 25556 19496 25562 19508
rect 27246 19496 27252 19508
rect 25556 19468 27252 19496
rect 25556 19456 25562 19468
rect 27246 19456 27252 19468
rect 27304 19456 27310 19508
rect 27338 19456 27344 19508
rect 27396 19496 27402 19508
rect 27433 19499 27491 19505
rect 27433 19496 27445 19499
rect 27396 19468 27445 19496
rect 27396 19456 27402 19468
rect 27433 19465 27445 19468
rect 27479 19465 27491 19499
rect 28905 19499 28963 19505
rect 28905 19496 28917 19499
rect 27433 19459 27491 19465
rect 27540 19468 28917 19496
rect 24486 19388 24492 19440
rect 24544 19428 24550 19440
rect 27540 19428 27568 19468
rect 28905 19465 28917 19468
rect 28951 19496 28963 19499
rect 28994 19496 29000 19508
rect 28951 19468 29000 19496
rect 28951 19465 28963 19468
rect 28905 19459 28963 19465
rect 28994 19456 29000 19468
rect 29052 19456 29058 19508
rect 30282 19456 30288 19508
rect 30340 19456 30346 19508
rect 31018 19456 31024 19508
rect 31076 19496 31082 19508
rect 31076 19468 31616 19496
rect 31076 19456 31082 19468
rect 27614 19437 27620 19440
rect 24544 19400 27568 19428
rect 27601 19431 27620 19437
rect 24544 19388 24550 19400
rect 27601 19397 27613 19431
rect 27601 19391 27620 19397
rect 27614 19388 27620 19391
rect 27672 19388 27678 19440
rect 27798 19388 27804 19440
rect 27856 19428 27862 19440
rect 31588 19437 31616 19468
rect 31662 19456 31668 19508
rect 31720 19496 31726 19508
rect 31720 19468 34744 19496
rect 31720 19456 31726 19468
rect 31573 19431 31631 19437
rect 27856 19400 30052 19428
rect 27856 19388 27862 19400
rect 30024 19372 30052 19400
rect 31343 19397 31401 19403
rect 25130 19320 25136 19372
rect 25188 19360 25194 19372
rect 25406 19360 25412 19372
rect 25188 19332 25412 19360
rect 25188 19320 25194 19332
rect 25406 19320 25412 19332
rect 25464 19360 25470 19372
rect 26326 19360 26332 19372
rect 25464 19332 26332 19360
rect 25464 19320 25470 19332
rect 26326 19320 26332 19332
rect 26384 19360 26390 19372
rect 28718 19360 28724 19372
rect 26384 19332 28724 19360
rect 26384 19320 26390 19332
rect 28718 19320 28724 19332
rect 28776 19320 28782 19372
rect 29273 19363 29331 19369
rect 29273 19329 29285 19363
rect 29319 19360 29331 19363
rect 29362 19360 29368 19372
rect 29319 19332 29368 19360
rect 29319 19329 29331 19332
rect 29273 19323 29331 19329
rect 29362 19320 29368 19332
rect 29420 19320 29426 19372
rect 29454 19320 29460 19372
rect 29512 19320 29518 19372
rect 29549 19363 29607 19369
rect 29549 19329 29561 19363
rect 29595 19360 29607 19363
rect 29914 19360 29920 19372
rect 29595 19332 29920 19360
rect 29595 19329 29607 19332
rect 29549 19323 29607 19329
rect 29914 19320 29920 19332
rect 29972 19320 29978 19372
rect 30006 19320 30012 19372
rect 30064 19360 30070 19372
rect 30469 19363 30527 19369
rect 30064 19332 30328 19360
rect 30064 19320 30070 19332
rect 23808 19264 24072 19292
rect 23808 19252 23814 19264
rect 29086 19252 29092 19304
rect 29144 19252 29150 19304
rect 29472 19292 29500 19320
rect 30098 19292 30104 19304
rect 29472 19264 30104 19292
rect 30098 19252 30104 19264
rect 30156 19252 30162 19304
rect 30190 19252 30196 19304
rect 30248 19252 30254 19304
rect 30300 19292 30328 19332
rect 30469 19329 30481 19363
rect 30515 19360 30527 19363
rect 30834 19360 30840 19372
rect 30515 19332 30840 19360
rect 30515 19329 30527 19332
rect 30469 19323 30527 19329
rect 30834 19320 30840 19332
rect 30892 19360 30898 19372
rect 31018 19360 31024 19372
rect 30892 19332 31024 19360
rect 30892 19320 30898 19332
rect 31018 19320 31024 19332
rect 31076 19320 31082 19372
rect 31343 19363 31355 19397
rect 31389 19363 31401 19397
rect 31573 19397 31585 19431
rect 31619 19397 31631 19431
rect 31573 19391 31631 19397
rect 32582 19388 32588 19440
rect 32640 19428 32646 19440
rect 33318 19428 33324 19440
rect 32640 19400 33324 19428
rect 32640 19388 32646 19400
rect 33318 19388 33324 19400
rect 33376 19388 33382 19440
rect 33962 19437 33968 19440
rect 33939 19431 33968 19437
rect 33939 19397 33951 19431
rect 33939 19391 33968 19397
rect 33962 19388 33968 19391
rect 34020 19388 34026 19440
rect 34146 19388 34152 19440
rect 34204 19388 34210 19440
rect 34517 19431 34575 19437
rect 34517 19397 34529 19431
rect 34563 19428 34575 19431
rect 34606 19428 34612 19440
rect 34563 19400 34612 19428
rect 34563 19397 34575 19400
rect 34517 19391 34575 19397
rect 34606 19388 34612 19400
rect 34664 19388 34670 19440
rect 31343 19360 31401 19363
rect 31343 19357 34008 19360
rect 31358 19332 34008 19357
rect 30653 19295 30711 19301
rect 30653 19292 30665 19295
rect 30300 19264 30665 19292
rect 30653 19261 30665 19264
rect 30699 19261 30711 19295
rect 33781 19295 33839 19301
rect 33781 19292 33793 19295
rect 30653 19255 30711 19261
rect 30760 19264 33793 19292
rect 18279 19196 18368 19224
rect 18279 19193 18291 19196
rect 18233 19187 18291 19193
rect 21818 19184 21824 19236
rect 21876 19184 21882 19236
rect 27706 19184 27712 19236
rect 27764 19224 27770 19236
rect 27764 19196 29040 19224
rect 27764 19184 27770 19196
rect 18322 19156 18328 19168
rect 16776 19128 18328 19156
rect 16393 19119 16451 19125
rect 18322 19116 18328 19128
rect 18380 19116 18386 19168
rect 27246 19116 27252 19168
rect 27304 19156 27310 19168
rect 27617 19159 27675 19165
rect 27617 19156 27629 19159
rect 27304 19128 27629 19156
rect 27304 19116 27310 19128
rect 27617 19125 27629 19128
rect 27663 19156 27675 19159
rect 28258 19156 28264 19168
rect 27663 19128 28264 19156
rect 27663 19125 27675 19128
rect 27617 19119 27675 19125
rect 28258 19116 28264 19128
rect 28316 19116 28322 19168
rect 29012 19156 29040 19196
rect 29270 19184 29276 19236
rect 29328 19224 29334 19236
rect 29365 19227 29423 19233
rect 29365 19224 29377 19227
rect 29328 19196 29377 19224
rect 29328 19184 29334 19196
rect 29365 19193 29377 19196
rect 29411 19193 29423 19227
rect 29365 19187 29423 19193
rect 29457 19227 29515 19233
rect 29457 19193 29469 19227
rect 29503 19224 29515 19227
rect 29638 19224 29644 19236
rect 29503 19196 29644 19224
rect 29503 19193 29515 19196
rect 29457 19187 29515 19193
rect 29638 19184 29644 19196
rect 29696 19224 29702 19236
rect 30760 19224 30788 19264
rect 33781 19261 33793 19264
rect 33827 19261 33839 19295
rect 33980 19292 34008 19332
rect 34054 19320 34060 19372
rect 34112 19320 34118 19372
rect 34238 19360 34244 19372
rect 34164 19332 34244 19360
rect 34164 19292 34192 19332
rect 34238 19320 34244 19332
rect 34296 19320 34302 19372
rect 34716 19369 34744 19468
rect 34790 19456 34796 19508
rect 34848 19496 34854 19508
rect 35161 19499 35219 19505
rect 35161 19496 35173 19499
rect 34848 19468 35173 19496
rect 34848 19456 34854 19468
rect 35161 19465 35173 19468
rect 35207 19465 35219 19499
rect 35161 19459 35219 19465
rect 35437 19499 35495 19505
rect 35437 19465 35449 19499
rect 35483 19496 35495 19499
rect 35526 19496 35532 19508
rect 35483 19468 35532 19496
rect 35483 19465 35495 19468
rect 35437 19459 35495 19465
rect 35526 19456 35532 19468
rect 35584 19456 35590 19508
rect 35802 19456 35808 19508
rect 35860 19496 35866 19508
rect 36725 19499 36783 19505
rect 35860 19468 36676 19496
rect 35860 19456 35866 19468
rect 36265 19431 36323 19437
rect 36265 19428 36277 19431
rect 34808 19400 36277 19428
rect 34425 19363 34483 19369
rect 34425 19329 34437 19363
rect 34471 19360 34483 19363
rect 34701 19363 34759 19369
rect 34471 19332 34652 19360
rect 34471 19329 34483 19332
rect 34425 19323 34483 19329
rect 33980 19264 34192 19292
rect 34624 19292 34652 19332
rect 34701 19329 34713 19363
rect 34747 19329 34759 19363
rect 34701 19323 34759 19329
rect 34808 19292 34836 19400
rect 36265 19397 36277 19400
rect 36311 19428 36323 19431
rect 36354 19428 36360 19440
rect 36311 19400 36360 19428
rect 36311 19397 36323 19400
rect 36265 19391 36323 19397
rect 36354 19388 36360 19400
rect 36412 19388 36418 19440
rect 34974 19320 34980 19372
rect 35032 19320 35038 19372
rect 35158 19320 35164 19372
rect 35216 19360 35222 19372
rect 35216 19332 35388 19360
rect 35216 19320 35222 19332
rect 34624 19264 34836 19292
rect 33781 19255 33839 19261
rect 34882 19252 34888 19304
rect 34940 19252 34946 19304
rect 35360 19292 35388 19332
rect 35434 19320 35440 19372
rect 35492 19360 35498 19372
rect 35621 19363 35679 19369
rect 35621 19360 35633 19363
rect 35492 19332 35633 19360
rect 35492 19320 35498 19332
rect 35621 19329 35633 19332
rect 35667 19329 35679 19363
rect 35621 19323 35679 19329
rect 35713 19363 35771 19369
rect 35713 19329 35725 19363
rect 35759 19329 35771 19363
rect 35713 19323 35771 19329
rect 35728 19292 35756 19323
rect 35802 19320 35808 19372
rect 35860 19320 35866 19372
rect 35989 19363 36047 19369
rect 35989 19329 36001 19363
rect 36035 19360 36047 19363
rect 36170 19360 36176 19372
rect 36035 19332 36176 19360
rect 36035 19329 36047 19332
rect 35989 19323 36047 19329
rect 36170 19320 36176 19332
rect 36228 19320 36234 19372
rect 36446 19320 36452 19372
rect 36504 19320 36510 19372
rect 36541 19363 36599 19369
rect 36541 19329 36553 19363
rect 36587 19329 36599 19363
rect 36648 19360 36676 19468
rect 36725 19465 36737 19499
rect 36771 19496 36783 19499
rect 37182 19496 37188 19508
rect 36771 19468 37188 19496
rect 36771 19465 36783 19468
rect 36725 19459 36783 19465
rect 37182 19456 37188 19468
rect 37240 19456 37246 19508
rect 38102 19456 38108 19508
rect 38160 19496 38166 19508
rect 38648 19499 38706 19505
rect 38160 19468 38516 19496
rect 38160 19456 38166 19468
rect 38488 19428 38516 19468
rect 38648 19465 38660 19499
rect 38694 19496 38706 19499
rect 39022 19496 39028 19508
rect 38694 19468 39028 19496
rect 38694 19465 38706 19468
rect 38648 19459 38706 19465
rect 39022 19456 39028 19468
rect 39080 19496 39086 19508
rect 39482 19496 39488 19508
rect 39080 19468 39488 19496
rect 39080 19456 39086 19468
rect 39482 19456 39488 19468
rect 39540 19456 39546 19508
rect 38488 19400 39068 19428
rect 39040 19369 39068 19400
rect 38381 19363 38439 19369
rect 38381 19360 38393 19363
rect 36648 19332 38393 19360
rect 36541 19323 36599 19329
rect 38381 19329 38393 19332
rect 38427 19360 38439 19363
rect 39025 19363 39083 19369
rect 38427 19332 38700 19360
rect 38427 19329 38439 19332
rect 38381 19323 38439 19329
rect 35360 19264 35756 19292
rect 29696 19196 30788 19224
rect 29696 19184 29702 19196
rect 30834 19184 30840 19236
rect 30892 19224 30898 19236
rect 30892 19196 31340 19224
rect 30892 19184 30898 19196
rect 29733 19159 29791 19165
rect 29733 19156 29745 19159
rect 29012 19128 29745 19156
rect 29733 19125 29745 19128
rect 29779 19125 29791 19159
rect 29733 19119 29791 19125
rect 29914 19116 29920 19168
rect 29972 19156 29978 19168
rect 30098 19156 30104 19168
rect 29972 19128 30104 19156
rect 29972 19116 29978 19128
rect 30098 19116 30104 19128
rect 30156 19116 30162 19168
rect 31202 19116 31208 19168
rect 31260 19116 31266 19168
rect 31312 19156 31340 19196
rect 34054 19184 34060 19236
rect 34112 19224 34118 19236
rect 34422 19224 34428 19236
rect 34112 19196 34428 19224
rect 34112 19184 34118 19196
rect 34422 19184 34428 19196
rect 34480 19184 34486 19236
rect 36170 19184 36176 19236
rect 36228 19224 36234 19236
rect 36556 19224 36584 19323
rect 38672 19292 38700 19332
rect 39025 19329 39037 19363
rect 39071 19329 39083 19363
rect 39025 19323 39083 19329
rect 39206 19292 39212 19304
rect 38672 19264 39212 19292
rect 39206 19252 39212 19264
rect 39264 19252 39270 19304
rect 36228 19196 36584 19224
rect 36228 19184 36234 19196
rect 31389 19159 31447 19165
rect 31389 19156 31401 19159
rect 31312 19128 31401 19156
rect 31389 19125 31401 19128
rect 31435 19125 31447 19159
rect 31389 19119 31447 19125
rect 33962 19116 33968 19168
rect 34020 19156 34026 19168
rect 35802 19156 35808 19168
rect 34020 19128 35808 19156
rect 34020 19116 34026 19128
rect 35802 19116 35808 19128
rect 35860 19116 35866 19168
rect 35894 19116 35900 19168
rect 35952 19156 35958 19168
rect 36265 19159 36323 19165
rect 36265 19156 36277 19159
rect 35952 19128 36277 19156
rect 35952 19116 35958 19128
rect 36265 19125 36277 19128
rect 36311 19125 36323 19159
rect 36265 19119 36323 19125
rect 36538 19116 36544 19168
rect 36596 19156 36602 19168
rect 36814 19156 36820 19168
rect 36596 19128 36820 19156
rect 36596 19116 36602 19128
rect 36814 19116 36820 19128
rect 36872 19116 36878 19168
rect 38657 19159 38715 19165
rect 38657 19125 38669 19159
rect 38703 19156 38715 19159
rect 38746 19156 38752 19168
rect 38703 19128 38752 19156
rect 38703 19125 38715 19128
rect 38657 19119 38715 19125
rect 38746 19116 38752 19128
rect 38804 19116 38810 19168
rect 1104 19066 40572 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 40572 19066
rect 1104 18992 40572 19014
rect 3329 18955 3387 18961
rect 3329 18921 3341 18955
rect 3375 18952 3387 18955
rect 4890 18952 4896 18964
rect 3375 18924 4896 18952
rect 3375 18921 3387 18924
rect 3329 18915 3387 18921
rect 4890 18912 4896 18924
rect 4948 18912 4954 18964
rect 5074 18912 5080 18964
rect 5132 18952 5138 18964
rect 5132 18924 7052 18952
rect 5132 18912 5138 18924
rect 3786 18844 3792 18896
rect 3844 18884 3850 18896
rect 3844 18856 5304 18884
rect 3844 18844 3850 18856
rect 1578 18776 1584 18828
rect 1636 18776 1642 18828
rect 3050 18776 3056 18828
rect 3108 18776 3114 18828
rect 4062 18776 4068 18828
rect 4120 18816 4126 18828
rect 4430 18816 4436 18828
rect 4120 18788 4436 18816
rect 4120 18776 4126 18788
rect 4430 18776 4436 18788
rect 4488 18816 4494 18828
rect 4893 18819 4951 18825
rect 4893 18816 4905 18819
rect 4488 18788 4905 18816
rect 4488 18776 4494 18788
rect 4893 18785 4905 18788
rect 4939 18816 4951 18819
rect 5074 18816 5080 18828
rect 4939 18788 5080 18816
rect 4939 18785 4951 18788
rect 4893 18779 4951 18785
rect 5074 18776 5080 18788
rect 5132 18776 5138 18828
rect 5166 18776 5172 18828
rect 5224 18776 5230 18828
rect 5276 18816 5304 18856
rect 7024 18828 7052 18924
rect 7650 18912 7656 18964
rect 7708 18912 7714 18964
rect 9490 18912 9496 18964
rect 9548 18912 9554 18964
rect 12618 18912 12624 18964
rect 12676 18912 12682 18964
rect 15838 18912 15844 18964
rect 15896 18912 15902 18964
rect 20622 18912 20628 18964
rect 20680 18952 20686 18964
rect 20809 18955 20867 18961
rect 20809 18952 20821 18955
rect 20680 18924 20821 18952
rect 20680 18912 20686 18924
rect 20809 18921 20821 18924
rect 20855 18921 20867 18955
rect 20809 18915 20867 18921
rect 21634 18912 21640 18964
rect 21692 18912 21698 18964
rect 23382 18912 23388 18964
rect 23440 18952 23446 18964
rect 24673 18955 24731 18961
rect 24673 18952 24685 18955
rect 23440 18924 24685 18952
rect 23440 18912 23446 18924
rect 24673 18921 24685 18924
rect 24719 18921 24731 18955
rect 24673 18915 24731 18921
rect 20254 18844 20260 18896
rect 20312 18884 20318 18896
rect 20441 18887 20499 18893
rect 20441 18884 20453 18887
rect 20312 18856 20453 18884
rect 20312 18844 20318 18856
rect 20441 18853 20453 18856
rect 20487 18853 20499 18887
rect 23106 18884 23112 18896
rect 20441 18847 20499 18853
rect 20640 18856 23112 18884
rect 5276 18788 6592 18816
rect 1854 18640 1860 18692
rect 1912 18640 1918 18692
rect 3068 18680 3096 18776
rect 4706 18708 4712 18760
rect 4764 18708 4770 18760
rect 4801 18751 4859 18757
rect 4801 18717 4813 18751
rect 4847 18748 4859 18751
rect 4982 18748 4988 18760
rect 4847 18720 4988 18748
rect 4847 18717 4859 18720
rect 4801 18711 4859 18717
rect 4982 18708 4988 18720
rect 5040 18708 5046 18760
rect 6564 18734 6592 18788
rect 7006 18776 7012 18828
rect 7064 18816 7070 18828
rect 8297 18819 8355 18825
rect 8297 18816 8309 18819
rect 7064 18788 8309 18816
rect 7064 18776 7070 18788
rect 8297 18785 8309 18788
rect 8343 18816 8355 18819
rect 10137 18819 10195 18825
rect 10137 18816 10149 18819
rect 8343 18788 10149 18816
rect 8343 18785 8355 18788
rect 8297 18779 8355 18785
rect 10137 18785 10149 18788
rect 10183 18816 10195 18819
rect 11146 18816 11152 18828
rect 10183 18788 11152 18816
rect 10183 18785 10195 18788
rect 10137 18779 10195 18785
rect 11146 18776 11152 18788
rect 11204 18776 11210 18828
rect 11238 18776 11244 18828
rect 11296 18816 11302 18828
rect 11296 18788 17264 18816
rect 11296 18776 11302 18788
rect 8021 18751 8079 18757
rect 8021 18717 8033 18751
rect 8067 18748 8079 18751
rect 8110 18748 8116 18760
rect 8067 18720 8116 18748
rect 8067 18717 8079 18720
rect 8021 18711 8079 18717
rect 8110 18708 8116 18720
rect 8168 18708 8174 18760
rect 8754 18708 8760 18760
rect 8812 18748 8818 18760
rect 9217 18751 9275 18757
rect 9217 18748 9229 18751
rect 8812 18720 9229 18748
rect 8812 18708 8818 18720
rect 9217 18717 9229 18720
rect 9263 18717 9275 18751
rect 9217 18711 9275 18717
rect 9398 18708 9404 18760
rect 9456 18708 9462 18760
rect 9861 18751 9919 18757
rect 9861 18717 9873 18751
rect 9907 18748 9919 18751
rect 10594 18748 10600 18760
rect 9907 18720 10600 18748
rect 9907 18717 9919 18720
rect 9861 18711 9919 18717
rect 10594 18708 10600 18720
rect 10652 18708 10658 18760
rect 10873 18751 10931 18757
rect 10873 18717 10885 18751
rect 10919 18717 10931 18751
rect 10873 18711 10931 18717
rect 3068 18666 3188 18680
rect 3082 18652 3188 18666
rect 3160 18612 3188 18652
rect 3234 18640 3240 18692
rect 3292 18680 3298 18692
rect 3292 18652 4936 18680
rect 3292 18640 3298 18652
rect 3786 18612 3792 18624
rect 3160 18584 3792 18612
rect 3786 18572 3792 18584
rect 3844 18572 3850 18624
rect 4062 18572 4068 18624
rect 4120 18612 4126 18624
rect 4341 18615 4399 18621
rect 4341 18612 4353 18615
rect 4120 18584 4353 18612
rect 4120 18572 4126 18584
rect 4341 18581 4353 18584
rect 4387 18581 4399 18615
rect 4908 18612 4936 18652
rect 5442 18640 5448 18692
rect 5500 18640 5506 18692
rect 10888 18680 10916 18711
rect 12250 18708 12256 18760
rect 12308 18750 12314 18760
rect 12308 18748 12434 18750
rect 12308 18722 12572 18748
rect 12308 18708 12314 18722
rect 12406 18720 12572 18722
rect 6748 18652 10916 18680
rect 6748 18612 6776 18652
rect 11146 18640 11152 18692
rect 11204 18640 11210 18692
rect 12544 18680 12572 18720
rect 12618 18708 12624 18760
rect 12676 18748 12682 18760
rect 13265 18751 13323 18757
rect 13265 18748 13277 18751
rect 12676 18720 13277 18748
rect 12676 18708 12682 18720
rect 13265 18717 13277 18720
rect 13311 18717 13323 18751
rect 13265 18711 13323 18717
rect 15930 18708 15936 18760
rect 15988 18708 15994 18760
rect 14090 18680 14096 18692
rect 12544 18652 14096 18680
rect 14090 18640 14096 18652
rect 14148 18640 14154 18692
rect 17236 18680 17264 18788
rect 20346 18708 20352 18760
rect 20404 18708 20410 18760
rect 20640 18757 20668 18856
rect 23106 18844 23112 18856
rect 23164 18884 23170 18896
rect 23750 18884 23756 18896
rect 23164 18856 23756 18884
rect 23164 18844 23170 18856
rect 23750 18844 23756 18856
rect 23808 18844 23814 18896
rect 24688 18884 24716 18915
rect 24946 18912 24952 18964
rect 25004 18952 25010 18964
rect 25133 18955 25191 18961
rect 25133 18952 25145 18955
rect 25004 18924 25145 18952
rect 25004 18912 25010 18924
rect 25133 18921 25145 18924
rect 25179 18921 25191 18955
rect 25133 18915 25191 18921
rect 26145 18955 26203 18961
rect 26145 18921 26157 18955
rect 26191 18952 26203 18955
rect 26510 18952 26516 18964
rect 26191 18924 26516 18952
rect 26191 18921 26203 18924
rect 26145 18915 26203 18921
rect 26510 18912 26516 18924
rect 26568 18912 26574 18964
rect 26786 18912 26792 18964
rect 26844 18952 26850 18964
rect 26881 18955 26939 18961
rect 26881 18952 26893 18955
rect 26844 18924 26893 18952
rect 26844 18912 26850 18924
rect 26881 18921 26893 18924
rect 26927 18921 26939 18955
rect 26881 18915 26939 18921
rect 27065 18955 27123 18961
rect 27065 18921 27077 18955
rect 27111 18921 27123 18955
rect 27065 18915 27123 18921
rect 25222 18884 25228 18896
rect 24688 18856 25228 18884
rect 25222 18844 25228 18856
rect 25280 18844 25286 18896
rect 26234 18844 26240 18896
rect 26292 18884 26298 18896
rect 26804 18884 26832 18912
rect 26292 18856 26832 18884
rect 27080 18884 27108 18915
rect 27430 18912 27436 18964
rect 27488 18912 27494 18964
rect 27614 18912 27620 18964
rect 27672 18912 27678 18964
rect 28718 18912 28724 18964
rect 28776 18952 28782 18964
rect 29733 18955 29791 18961
rect 29733 18952 29745 18955
rect 28776 18924 29745 18952
rect 28776 18912 28782 18924
rect 29733 18921 29745 18924
rect 29779 18921 29791 18955
rect 29733 18915 29791 18921
rect 30558 18912 30564 18964
rect 30616 18952 30622 18964
rect 32766 18952 32772 18964
rect 30616 18924 32772 18952
rect 30616 18912 30622 18924
rect 32766 18912 32772 18924
rect 32824 18912 32830 18964
rect 35526 18912 35532 18964
rect 35584 18952 35590 18964
rect 36538 18952 36544 18964
rect 35584 18924 36544 18952
rect 35584 18912 35590 18924
rect 36538 18912 36544 18924
rect 36596 18912 36602 18964
rect 27798 18884 27804 18896
rect 27080 18856 27804 18884
rect 26292 18844 26298 18856
rect 27798 18844 27804 18856
rect 27856 18844 27862 18896
rect 28166 18844 28172 18896
rect 28224 18844 28230 18896
rect 29270 18844 29276 18896
rect 29328 18844 29334 18896
rect 31018 18844 31024 18896
rect 31076 18884 31082 18896
rect 31662 18884 31668 18896
rect 31076 18856 31668 18884
rect 31076 18844 31082 18856
rect 31662 18844 31668 18856
rect 31720 18844 31726 18896
rect 34606 18844 34612 18896
rect 34664 18884 34670 18896
rect 35986 18884 35992 18896
rect 34664 18856 35992 18884
rect 34664 18844 34670 18856
rect 35986 18844 35992 18856
rect 36044 18844 36050 18896
rect 21266 18776 21272 18828
rect 21324 18816 21330 18828
rect 21324 18788 22048 18816
rect 21324 18776 21330 18788
rect 22020 18760 22048 18788
rect 24578 18776 24584 18828
rect 24636 18816 24642 18828
rect 30926 18816 30932 18828
rect 24636 18788 26096 18816
rect 24636 18776 24642 18788
rect 20625 18751 20683 18757
rect 20625 18717 20637 18751
rect 20671 18717 20683 18751
rect 20625 18711 20683 18717
rect 20714 18708 20720 18760
rect 20772 18748 20778 18760
rect 20901 18751 20959 18757
rect 20901 18748 20913 18751
rect 20772 18720 20913 18748
rect 20772 18708 20778 18720
rect 20901 18717 20913 18720
rect 20947 18717 20959 18751
rect 20901 18711 20959 18717
rect 21085 18751 21143 18757
rect 21085 18717 21097 18751
rect 21131 18748 21143 18751
rect 21634 18748 21640 18760
rect 21131 18720 21640 18748
rect 21131 18717 21143 18720
rect 21085 18711 21143 18717
rect 21634 18708 21640 18720
rect 21692 18708 21698 18760
rect 21818 18708 21824 18760
rect 21876 18748 21882 18760
rect 21913 18751 21971 18757
rect 21913 18748 21925 18751
rect 21876 18720 21925 18748
rect 21876 18708 21882 18720
rect 21913 18717 21925 18720
rect 21959 18717 21971 18751
rect 21913 18711 21971 18717
rect 22002 18708 22008 18760
rect 22060 18708 22066 18760
rect 22097 18751 22155 18757
rect 22097 18717 22109 18751
rect 22143 18717 22155 18751
rect 22097 18711 22155 18717
rect 22281 18751 22339 18757
rect 22281 18717 22293 18751
rect 22327 18748 22339 18751
rect 23198 18748 23204 18760
rect 22327 18720 23204 18748
rect 22327 18717 22339 18720
rect 22281 18711 22339 18717
rect 19702 18680 19708 18692
rect 17236 18652 19708 18680
rect 19702 18640 19708 18652
rect 19760 18640 19766 18692
rect 4908 18584 6776 18612
rect 6917 18615 6975 18621
rect 4341 18575 4399 18581
rect 6917 18581 6929 18615
rect 6963 18612 6975 18615
rect 7190 18612 7196 18624
rect 6963 18584 7196 18612
rect 6963 18581 6975 18584
rect 6917 18575 6975 18581
rect 7190 18572 7196 18584
rect 7248 18612 7254 18624
rect 7742 18612 7748 18624
rect 7248 18584 7748 18612
rect 7248 18572 7254 18584
rect 7742 18572 7748 18584
rect 7800 18572 7806 18624
rect 8110 18572 8116 18624
rect 8168 18572 8174 18624
rect 9309 18615 9367 18621
rect 9309 18581 9321 18615
rect 9355 18612 9367 18615
rect 9858 18612 9864 18624
rect 9355 18584 9864 18612
rect 9355 18581 9367 18584
rect 9309 18575 9367 18581
rect 9858 18572 9864 18584
rect 9916 18572 9922 18624
rect 9950 18572 9956 18624
rect 10008 18572 10014 18624
rect 10042 18572 10048 18624
rect 10100 18612 10106 18624
rect 12618 18612 12624 18624
rect 10100 18584 12624 18612
rect 10100 18572 10106 18584
rect 12618 18572 12624 18584
rect 12676 18572 12682 18624
rect 12710 18572 12716 18624
rect 12768 18572 12774 18624
rect 17954 18572 17960 18624
rect 18012 18612 18018 18624
rect 21269 18615 21327 18621
rect 21269 18612 21281 18615
rect 18012 18584 21281 18612
rect 18012 18572 18018 18584
rect 21269 18581 21281 18584
rect 21315 18581 21327 18615
rect 21269 18575 21327 18581
rect 21634 18572 21640 18624
rect 21692 18612 21698 18624
rect 22112 18612 22140 18711
rect 23198 18708 23204 18720
rect 23256 18748 23262 18760
rect 24394 18748 24400 18760
rect 23256 18720 24400 18748
rect 23256 18708 23262 18720
rect 24394 18708 24400 18720
rect 24452 18748 24458 18760
rect 24452 18720 24900 18748
rect 24452 18708 24458 18720
rect 24872 18689 24900 18720
rect 24946 18708 24952 18760
rect 25004 18748 25010 18760
rect 25685 18751 25743 18757
rect 25685 18748 25697 18751
rect 25004 18720 25697 18748
rect 25004 18708 25010 18720
rect 25685 18717 25697 18720
rect 25731 18717 25743 18751
rect 25685 18711 25743 18717
rect 25774 18708 25780 18760
rect 25832 18708 25838 18760
rect 25869 18751 25927 18757
rect 25869 18717 25881 18751
rect 25915 18717 25927 18751
rect 25869 18711 25927 18717
rect 24857 18683 24915 18689
rect 24857 18649 24869 18683
rect 24903 18649 24915 18683
rect 25317 18683 25375 18689
rect 24857 18643 24915 18649
rect 24964 18652 25268 18680
rect 21692 18584 22140 18612
rect 21692 18572 21698 18584
rect 22186 18572 22192 18624
rect 22244 18612 22250 18624
rect 24489 18615 24547 18621
rect 24489 18612 24501 18615
rect 22244 18584 24501 18612
rect 22244 18572 22250 18584
rect 24489 18581 24501 18584
rect 24535 18581 24547 18615
rect 24489 18575 24547 18581
rect 24578 18572 24584 18624
rect 24636 18612 24642 18624
rect 24964 18621 24992 18652
rect 25130 18621 25136 18624
rect 24673 18615 24731 18621
rect 24673 18612 24685 18615
rect 24636 18584 24685 18612
rect 24636 18572 24642 18584
rect 24673 18581 24685 18584
rect 24719 18581 24731 18615
rect 24673 18575 24731 18581
rect 24949 18615 25007 18621
rect 24949 18581 24961 18615
rect 24995 18581 25007 18615
rect 24949 18575 25007 18581
rect 25117 18615 25136 18621
rect 25117 18581 25129 18615
rect 25117 18575 25136 18581
rect 25130 18572 25136 18575
rect 25188 18572 25194 18624
rect 25240 18612 25268 18652
rect 25317 18649 25329 18683
rect 25363 18680 25375 18683
rect 25406 18680 25412 18692
rect 25363 18652 25412 18680
rect 25363 18649 25375 18652
rect 25317 18643 25375 18649
rect 25406 18640 25412 18652
rect 25464 18640 25470 18692
rect 25884 18680 25912 18711
rect 25958 18708 25964 18760
rect 26016 18708 26022 18760
rect 26068 18748 26096 18788
rect 27816 18788 30932 18816
rect 27614 18748 27620 18760
rect 26068 18720 27082 18748
rect 27019 18717 27082 18720
rect 27019 18683 27031 18717
rect 27065 18686 27082 18717
rect 27264 18720 27620 18748
rect 27264 18689 27292 18720
rect 27614 18708 27620 18720
rect 27672 18708 27678 18760
rect 27816 18689 27844 18788
rect 30926 18776 30932 18788
rect 30984 18776 30990 18828
rect 34422 18816 34428 18828
rect 31036 18788 34428 18816
rect 27890 18708 27896 18760
rect 27948 18748 27954 18760
rect 28537 18751 28595 18757
rect 28537 18748 28549 18751
rect 27948 18720 28549 18748
rect 27948 18708 27954 18720
rect 28537 18717 28549 18720
rect 28583 18748 28595 18751
rect 28718 18748 28724 18760
rect 28583 18720 28724 18748
rect 28583 18717 28595 18720
rect 28537 18711 28595 18717
rect 28718 18708 28724 18720
rect 28776 18708 28782 18760
rect 28994 18708 29000 18760
rect 29052 18748 29058 18760
rect 29089 18751 29147 18757
rect 29089 18748 29101 18751
rect 29052 18720 29101 18748
rect 29052 18708 29058 18720
rect 29089 18717 29101 18720
rect 29135 18717 29147 18751
rect 29089 18711 29147 18717
rect 29362 18708 29368 18760
rect 29420 18708 29426 18760
rect 29914 18748 29920 18760
rect 29656 18720 29920 18748
rect 27065 18683 27077 18686
rect 25884 18652 26004 18680
rect 27019 18677 27077 18683
rect 27249 18683 27307 18689
rect 25976 18624 26004 18652
rect 27249 18649 27261 18683
rect 27295 18649 27307 18683
rect 27249 18643 27307 18649
rect 27801 18683 27859 18689
rect 27801 18649 27813 18683
rect 27847 18649 27859 18683
rect 27801 18643 27859 18649
rect 28350 18640 28356 18692
rect 28408 18640 28414 18692
rect 28626 18640 28632 18692
rect 28684 18680 28690 18692
rect 29656 18689 29684 18720
rect 29914 18708 29920 18720
rect 29972 18708 29978 18760
rect 30193 18751 30251 18757
rect 30193 18717 30205 18751
rect 30239 18717 30251 18751
rect 30193 18711 30251 18717
rect 28905 18683 28963 18689
rect 28905 18680 28917 18683
rect 28684 18652 28917 18680
rect 28684 18640 28690 18652
rect 28905 18649 28917 18652
rect 28951 18649 28963 18683
rect 28905 18643 28963 18649
rect 29641 18683 29699 18689
rect 29641 18649 29653 18683
rect 29687 18649 29699 18683
rect 30208 18680 30236 18711
rect 30282 18708 30288 18760
rect 30340 18708 30346 18760
rect 31036 18757 31064 18788
rect 34422 18776 34428 18788
rect 34480 18816 34486 18828
rect 35069 18819 35127 18825
rect 35069 18816 35081 18819
rect 34480 18788 35081 18816
rect 34480 18776 34486 18788
rect 35069 18785 35081 18788
rect 35115 18785 35127 18819
rect 35069 18779 35127 18785
rect 35728 18788 36032 18816
rect 31021 18751 31079 18757
rect 31021 18717 31033 18751
rect 31067 18717 31079 18751
rect 31021 18711 31079 18717
rect 31202 18708 31208 18760
rect 31260 18708 31266 18760
rect 31389 18751 31447 18757
rect 31389 18717 31401 18751
rect 31435 18748 31447 18751
rect 31478 18748 31484 18760
rect 31435 18720 31484 18748
rect 31435 18717 31447 18720
rect 31389 18711 31447 18717
rect 31478 18708 31484 18720
rect 31536 18708 31542 18760
rect 31665 18751 31723 18757
rect 31665 18717 31677 18751
rect 31711 18748 31723 18751
rect 31754 18748 31760 18760
rect 31711 18720 31760 18748
rect 31711 18717 31723 18720
rect 31665 18711 31723 18717
rect 31754 18708 31760 18720
rect 31812 18708 31818 18760
rect 34698 18708 34704 18760
rect 34756 18748 34762 18760
rect 34885 18751 34943 18757
rect 34885 18748 34897 18751
rect 34756 18720 34897 18748
rect 34756 18708 34762 18720
rect 34885 18717 34897 18720
rect 34931 18717 34943 18751
rect 34885 18711 34943 18717
rect 35342 18708 35348 18760
rect 35400 18748 35406 18760
rect 35621 18751 35679 18757
rect 35621 18748 35633 18751
rect 35400 18720 35633 18748
rect 35400 18708 35406 18720
rect 35621 18717 35633 18720
rect 35667 18717 35679 18751
rect 35621 18711 35679 18717
rect 30926 18680 30932 18692
rect 30208 18652 30932 18680
rect 29641 18643 29699 18649
rect 30926 18640 30932 18652
rect 30984 18640 30990 18692
rect 31297 18683 31355 18689
rect 31297 18649 31309 18683
rect 31343 18649 31355 18683
rect 31846 18680 31852 18692
rect 31297 18643 31355 18649
rect 31726 18652 31852 18680
rect 25682 18612 25688 18624
rect 25240 18584 25688 18612
rect 25682 18572 25688 18584
rect 25740 18572 25746 18624
rect 25958 18572 25964 18624
rect 26016 18572 26022 18624
rect 27430 18572 27436 18624
rect 27488 18612 27494 18624
rect 27591 18615 27649 18621
rect 27591 18612 27603 18615
rect 27488 18584 27603 18612
rect 27488 18572 27494 18584
rect 27591 18581 27603 18584
rect 27637 18581 27649 18615
rect 27591 18575 27649 18581
rect 27982 18572 27988 18624
rect 28040 18612 28046 18624
rect 28721 18615 28779 18621
rect 28721 18612 28733 18615
rect 28040 18584 28733 18612
rect 28040 18572 28046 18584
rect 28721 18581 28733 18584
rect 28767 18581 28779 18615
rect 28721 18575 28779 18581
rect 28810 18572 28816 18624
rect 28868 18612 28874 18624
rect 29270 18612 29276 18624
rect 28868 18584 29276 18612
rect 28868 18572 28874 18584
rect 29270 18572 29276 18584
rect 29328 18572 29334 18624
rect 29914 18572 29920 18624
rect 29972 18612 29978 18624
rect 30190 18612 30196 18624
rect 29972 18584 30196 18612
rect 29972 18572 29978 18584
rect 30190 18572 30196 18584
rect 30248 18612 30254 18624
rect 30469 18615 30527 18621
rect 30469 18612 30481 18615
rect 30248 18584 30481 18612
rect 30248 18572 30254 18584
rect 30469 18581 30481 18584
rect 30515 18612 30527 18615
rect 31312 18612 31340 18643
rect 30515 18584 31340 18612
rect 31573 18615 31631 18621
rect 30515 18581 30527 18584
rect 30469 18575 30527 18581
rect 31573 18581 31585 18615
rect 31619 18612 31631 18615
rect 31726 18612 31754 18652
rect 31846 18640 31852 18652
rect 31904 18640 31910 18692
rect 32858 18640 32864 18692
rect 32916 18680 32922 18692
rect 35728 18680 35756 18788
rect 35802 18708 35808 18760
rect 35860 18708 35866 18760
rect 35894 18708 35900 18760
rect 35952 18708 35958 18760
rect 36004 18757 36032 18788
rect 38930 18776 38936 18828
rect 38988 18816 38994 18828
rect 39301 18819 39359 18825
rect 39301 18816 39313 18819
rect 38988 18788 39313 18816
rect 38988 18776 38994 18788
rect 39301 18785 39313 18788
rect 39347 18785 39359 18819
rect 39301 18779 39359 18785
rect 35989 18751 36047 18757
rect 35989 18717 36001 18751
rect 36035 18717 36047 18751
rect 35989 18711 36047 18717
rect 39025 18751 39083 18757
rect 39025 18717 39037 18751
rect 39071 18748 39083 18751
rect 39114 18748 39120 18760
rect 39071 18720 39120 18748
rect 39071 18717 39083 18720
rect 39025 18711 39083 18717
rect 39114 18708 39120 18720
rect 39172 18708 39178 18760
rect 39206 18708 39212 18760
rect 39264 18708 39270 18760
rect 32916 18652 35756 18680
rect 32916 18640 32922 18652
rect 31619 18584 31754 18612
rect 32033 18615 32091 18621
rect 31619 18581 31631 18584
rect 31573 18575 31631 18581
rect 32033 18581 32045 18615
rect 32079 18612 32091 18615
rect 32214 18612 32220 18624
rect 32079 18584 32220 18612
rect 32079 18581 32091 18584
rect 32033 18575 32091 18581
rect 32214 18572 32220 18584
rect 32272 18572 32278 18624
rect 34606 18572 34612 18624
rect 34664 18612 34670 18624
rect 34701 18615 34759 18621
rect 34701 18612 34713 18615
rect 34664 18584 34713 18612
rect 34664 18572 34670 18584
rect 34701 18581 34713 18584
rect 34747 18581 34759 18615
rect 34701 18575 34759 18581
rect 36170 18572 36176 18624
rect 36228 18572 36234 18624
rect 38562 18572 38568 18624
rect 38620 18612 38626 18624
rect 38841 18615 38899 18621
rect 38841 18612 38853 18615
rect 38620 18584 38853 18612
rect 38620 18572 38626 18584
rect 38841 18581 38853 18584
rect 38887 18581 38899 18615
rect 38841 18575 38899 18581
rect 1104 18522 40572 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 40572 18522
rect 1104 18448 40572 18470
rect 1854 18368 1860 18420
rect 1912 18408 1918 18420
rect 2685 18411 2743 18417
rect 2685 18408 2697 18411
rect 1912 18380 2697 18408
rect 1912 18368 1918 18380
rect 2685 18377 2697 18380
rect 2731 18377 2743 18411
rect 2685 18371 2743 18377
rect 3145 18411 3203 18417
rect 3145 18377 3157 18411
rect 3191 18408 3203 18411
rect 3326 18408 3332 18420
rect 3191 18380 3332 18408
rect 3191 18377 3203 18380
rect 3145 18371 3203 18377
rect 3326 18368 3332 18380
rect 3384 18408 3390 18420
rect 3694 18408 3700 18420
rect 3384 18380 3700 18408
rect 3384 18368 3390 18380
rect 3694 18368 3700 18380
rect 3752 18368 3758 18420
rect 4798 18408 4804 18420
rect 3896 18380 4804 18408
rect 2498 18300 2504 18352
rect 2556 18340 2562 18352
rect 3896 18340 3924 18380
rect 4798 18368 4804 18380
rect 4856 18368 4862 18420
rect 5442 18368 5448 18420
rect 5500 18408 5506 18420
rect 6365 18411 6423 18417
rect 6365 18408 6377 18411
rect 5500 18380 6377 18408
rect 5500 18368 5506 18380
rect 6365 18377 6377 18380
rect 6411 18377 6423 18411
rect 6365 18371 6423 18377
rect 8110 18368 8116 18420
rect 8168 18408 8174 18420
rect 10042 18408 10048 18420
rect 8168 18380 10048 18408
rect 8168 18368 8174 18380
rect 10042 18368 10048 18380
rect 10100 18368 10106 18420
rect 11146 18368 11152 18420
rect 11204 18408 11210 18420
rect 11701 18411 11759 18417
rect 11701 18408 11713 18411
rect 11204 18380 11713 18408
rect 11204 18368 11210 18380
rect 11701 18377 11713 18380
rect 11747 18377 11759 18411
rect 11701 18371 11759 18377
rect 12069 18411 12127 18417
rect 12069 18377 12081 18411
rect 12115 18408 12127 18411
rect 12710 18408 12716 18420
rect 12115 18380 12716 18408
rect 12115 18377 12127 18380
rect 12069 18371 12127 18377
rect 12710 18368 12716 18380
rect 12768 18368 12774 18420
rect 14182 18368 14188 18420
rect 14240 18408 14246 18420
rect 14277 18411 14335 18417
rect 14277 18408 14289 18411
rect 14240 18380 14289 18408
rect 14240 18368 14246 18380
rect 14277 18377 14289 18380
rect 14323 18377 14335 18411
rect 14277 18371 14335 18377
rect 15933 18411 15991 18417
rect 15933 18377 15945 18411
rect 15979 18408 15991 18411
rect 16022 18408 16028 18420
rect 15979 18380 16028 18408
rect 15979 18377 15991 18380
rect 15933 18371 15991 18377
rect 16022 18368 16028 18380
rect 16080 18368 16086 18420
rect 16758 18368 16764 18420
rect 16816 18368 16822 18420
rect 20254 18368 20260 18420
rect 20312 18408 20318 18420
rect 26789 18411 26847 18417
rect 20312 18380 25728 18408
rect 20312 18368 20318 18380
rect 2556 18312 3924 18340
rect 2556 18300 2562 18312
rect 3804 18281 3832 18312
rect 4062 18300 4068 18352
rect 4120 18300 4126 18352
rect 4154 18300 4160 18352
rect 4212 18340 4218 18352
rect 4212 18312 4554 18340
rect 4212 18300 4218 18312
rect 5350 18300 5356 18352
rect 5408 18340 5414 18352
rect 6825 18343 6883 18349
rect 6825 18340 6837 18343
rect 5408 18312 6837 18340
rect 5408 18300 5414 18312
rect 6825 18309 6837 18312
rect 6871 18340 6883 18343
rect 7834 18340 7840 18352
rect 6871 18312 7840 18340
rect 6871 18309 6883 18312
rect 6825 18303 6883 18309
rect 7834 18300 7840 18312
rect 7892 18300 7898 18352
rect 12161 18343 12219 18349
rect 12161 18309 12173 18343
rect 12207 18340 12219 18343
rect 12802 18340 12808 18352
rect 12207 18312 12808 18340
rect 12207 18309 12219 18312
rect 12161 18303 12219 18309
rect 12802 18300 12808 18312
rect 12860 18300 12866 18352
rect 14090 18340 14096 18352
rect 14030 18312 14096 18340
rect 14090 18300 14096 18312
rect 14148 18340 14154 18352
rect 16298 18340 16304 18352
rect 14148 18312 16304 18340
rect 14148 18300 14154 18312
rect 16298 18300 16304 18312
rect 16356 18300 16362 18352
rect 3053 18275 3111 18281
rect 3053 18241 3065 18275
rect 3099 18272 3111 18275
rect 3789 18275 3847 18281
rect 3099 18244 3740 18272
rect 3099 18241 3111 18244
rect 3053 18235 3111 18241
rect 3329 18207 3387 18213
rect 3329 18173 3341 18207
rect 3375 18204 3387 18207
rect 3712 18204 3740 18244
rect 3789 18241 3801 18275
rect 3835 18241 3847 18275
rect 3789 18235 3847 18241
rect 6733 18275 6791 18281
rect 6733 18241 6745 18275
rect 6779 18272 6791 18275
rect 7193 18275 7251 18281
rect 7193 18272 7205 18275
rect 6779 18244 7205 18272
rect 6779 18241 6791 18244
rect 6733 18235 6791 18241
rect 7193 18241 7205 18244
rect 7239 18241 7251 18275
rect 7193 18235 7251 18241
rect 7742 18232 7748 18284
rect 7800 18232 7806 18284
rect 15562 18232 15568 18284
rect 15620 18232 15626 18284
rect 15930 18232 15936 18284
rect 15988 18272 15994 18284
rect 16117 18275 16175 18281
rect 16117 18272 16129 18275
rect 15988 18244 16129 18272
rect 15988 18232 15994 18244
rect 16117 18241 16129 18244
rect 16163 18241 16175 18275
rect 16117 18235 16175 18241
rect 16393 18275 16451 18281
rect 16393 18241 16405 18275
rect 16439 18272 16451 18275
rect 16776 18272 16804 18368
rect 22278 18340 22284 18352
rect 22112 18312 22284 18340
rect 16439 18244 16804 18272
rect 17037 18275 17095 18281
rect 16439 18241 16451 18244
rect 16393 18235 16451 18241
rect 17037 18241 17049 18275
rect 17083 18272 17095 18275
rect 21818 18272 21824 18284
rect 17083 18244 21824 18272
rect 17083 18241 17095 18244
rect 17037 18235 17095 18241
rect 21818 18232 21824 18244
rect 21876 18232 21882 18284
rect 22112 18281 22140 18312
rect 22278 18300 22284 18312
rect 22336 18300 22342 18352
rect 22097 18275 22155 18281
rect 22097 18241 22109 18275
rect 22143 18241 22155 18275
rect 22097 18235 22155 18241
rect 22186 18232 22192 18284
rect 22244 18232 22250 18284
rect 22370 18232 22376 18284
rect 22428 18232 22434 18284
rect 22465 18275 22523 18281
rect 22465 18241 22477 18275
rect 22511 18241 22523 18275
rect 22465 18235 22523 18241
rect 4614 18204 4620 18216
rect 3375 18176 3648 18204
rect 3712 18176 4620 18204
rect 3375 18173 3387 18176
rect 3329 18167 3387 18173
rect 3620 18068 3648 18176
rect 4614 18164 4620 18176
rect 4672 18164 4678 18216
rect 5534 18164 5540 18216
rect 5592 18164 5598 18216
rect 7006 18164 7012 18216
rect 7064 18164 7070 18216
rect 11054 18164 11060 18216
rect 11112 18204 11118 18216
rect 12250 18204 12256 18216
rect 11112 18176 12256 18204
rect 11112 18164 11118 18176
rect 12250 18164 12256 18176
rect 12308 18164 12314 18216
rect 12529 18207 12587 18213
rect 12529 18173 12541 18207
rect 12575 18173 12587 18207
rect 12529 18167 12587 18173
rect 5442 18096 5448 18148
rect 5500 18136 5506 18148
rect 7466 18136 7472 18148
rect 5500 18108 7472 18136
rect 5500 18096 5506 18108
rect 7466 18096 7472 18108
rect 7524 18096 7530 18148
rect 7558 18096 7564 18148
rect 7616 18136 7622 18148
rect 12434 18136 12440 18148
rect 7616 18108 12440 18136
rect 7616 18096 7622 18108
rect 12434 18096 12440 18108
rect 12492 18096 12498 18148
rect 4430 18068 4436 18080
rect 3620 18040 4436 18068
rect 4430 18028 4436 18040
rect 4488 18028 4494 18080
rect 4706 18028 4712 18080
rect 4764 18068 4770 18080
rect 9214 18068 9220 18080
rect 4764 18040 9220 18068
rect 4764 18028 4770 18040
rect 9214 18028 9220 18040
rect 9272 18028 9278 18080
rect 12544 18068 12572 18167
rect 12802 18164 12808 18216
rect 12860 18164 12866 18216
rect 13262 18164 13268 18216
rect 13320 18204 13326 18216
rect 15381 18207 15439 18213
rect 15381 18204 15393 18207
rect 13320 18176 15393 18204
rect 13320 18164 13326 18176
rect 15381 18173 15393 18176
rect 15427 18173 15439 18207
rect 15381 18167 15439 18173
rect 15841 18207 15899 18213
rect 15841 18173 15853 18207
rect 15887 18204 15899 18207
rect 16209 18207 16267 18213
rect 16209 18204 16221 18207
rect 15887 18176 16221 18204
rect 15887 18173 15899 18176
rect 15841 18167 15899 18173
rect 16209 18173 16221 18176
rect 16255 18204 16267 18207
rect 18138 18204 18144 18216
rect 16255 18176 18144 18204
rect 16255 18173 16267 18176
rect 16209 18167 16267 18173
rect 18138 18164 18144 18176
rect 18196 18164 18202 18216
rect 15470 18136 15476 18148
rect 14200 18108 15476 18136
rect 14200 18068 14228 18108
rect 15470 18096 15476 18108
rect 15528 18096 15534 18148
rect 16301 18139 16359 18145
rect 16301 18105 16313 18139
rect 16347 18136 16359 18139
rect 16574 18136 16580 18148
rect 16347 18108 16580 18136
rect 16347 18105 16359 18108
rect 16301 18099 16359 18105
rect 16574 18096 16580 18108
rect 16632 18096 16638 18148
rect 12544 18040 14228 18068
rect 15746 18028 15752 18080
rect 15804 18028 15810 18080
rect 18598 18028 18604 18080
rect 18656 18068 18662 18080
rect 22204 18068 22232 18232
rect 22480 18204 22508 18235
rect 23934 18232 23940 18284
rect 23992 18272 23998 18284
rect 24397 18275 24455 18281
rect 24397 18272 24409 18275
rect 23992 18244 24409 18272
rect 23992 18232 23998 18244
rect 24397 18241 24409 18244
rect 24443 18241 24455 18275
rect 24397 18235 24455 18241
rect 24670 18232 24676 18284
rect 24728 18232 24734 18284
rect 24118 18204 24124 18216
rect 22480 18176 24124 18204
rect 24118 18164 24124 18176
rect 24176 18164 24182 18216
rect 24489 18207 24547 18213
rect 24489 18173 24501 18207
rect 24535 18204 24547 18207
rect 24762 18204 24768 18216
rect 24535 18176 24768 18204
rect 24535 18173 24547 18176
rect 24489 18167 24547 18173
rect 24762 18164 24768 18176
rect 24820 18164 24826 18216
rect 25700 18204 25728 18380
rect 26789 18377 26801 18411
rect 26835 18408 26847 18411
rect 27154 18408 27160 18420
rect 26835 18380 27160 18408
rect 26835 18377 26847 18380
rect 26789 18371 26847 18377
rect 27154 18368 27160 18380
rect 27212 18368 27218 18420
rect 27430 18368 27436 18420
rect 27488 18408 27494 18420
rect 31570 18408 31576 18420
rect 27488 18380 31576 18408
rect 27488 18368 27494 18380
rect 31570 18368 31576 18380
rect 31628 18368 31634 18420
rect 31726 18380 32444 18408
rect 25774 18300 25780 18352
rect 25832 18340 25838 18352
rect 27893 18343 27951 18349
rect 25832 18312 26372 18340
rect 25832 18300 25838 18312
rect 26050 18232 26056 18284
rect 26108 18272 26114 18284
rect 26344 18281 26372 18312
rect 27893 18309 27905 18343
rect 27939 18340 27951 18343
rect 28166 18340 28172 18352
rect 27939 18312 28172 18340
rect 27939 18309 27951 18312
rect 27893 18303 27951 18309
rect 28166 18300 28172 18312
rect 28224 18300 28230 18352
rect 31726 18340 31754 18380
rect 29932 18312 31754 18340
rect 26145 18275 26203 18281
rect 26145 18272 26157 18275
rect 26108 18244 26157 18272
rect 26108 18232 26114 18244
rect 26145 18241 26157 18244
rect 26191 18241 26203 18275
rect 26145 18235 26203 18241
rect 26329 18275 26387 18281
rect 26329 18241 26341 18275
rect 26375 18241 26387 18275
rect 26329 18235 26387 18241
rect 26421 18275 26479 18281
rect 26421 18241 26433 18275
rect 26467 18241 26479 18275
rect 26421 18235 26479 18241
rect 26436 18204 26464 18235
rect 26510 18232 26516 18284
rect 26568 18232 26574 18284
rect 27062 18232 27068 18284
rect 27120 18272 27126 18284
rect 27157 18275 27215 18281
rect 27157 18272 27169 18275
rect 27120 18244 27169 18272
rect 27120 18232 27126 18244
rect 27157 18241 27169 18244
rect 27203 18241 27215 18275
rect 27157 18235 27215 18241
rect 27341 18275 27399 18281
rect 27341 18241 27353 18275
rect 27387 18272 27399 18275
rect 27706 18272 27712 18284
rect 27387 18244 27712 18272
rect 27387 18241 27399 18244
rect 27341 18235 27399 18241
rect 27706 18232 27712 18244
rect 27764 18232 27770 18284
rect 27982 18232 27988 18284
rect 28040 18272 28046 18284
rect 28077 18275 28135 18281
rect 28077 18272 28089 18275
rect 28040 18244 28089 18272
rect 28040 18232 28046 18244
rect 28077 18241 28089 18244
rect 28123 18241 28135 18275
rect 28077 18235 28135 18241
rect 26786 18204 26792 18216
rect 25700 18176 26372 18204
rect 26436 18176 26792 18204
rect 24581 18139 24639 18145
rect 24581 18105 24593 18139
rect 24627 18136 24639 18139
rect 26234 18136 26240 18148
rect 24627 18108 26240 18136
rect 24627 18105 24639 18108
rect 24581 18099 24639 18105
rect 26234 18096 26240 18108
rect 26292 18096 26298 18148
rect 26344 18136 26372 18176
rect 26786 18164 26792 18176
rect 26844 18164 26850 18216
rect 27246 18164 27252 18216
rect 27304 18204 27310 18216
rect 29932 18204 29960 18312
rect 31846 18300 31852 18352
rect 31904 18340 31910 18352
rect 32309 18343 32367 18349
rect 32309 18340 32321 18343
rect 31904 18312 32321 18340
rect 31904 18300 31910 18312
rect 32309 18309 32321 18312
rect 32355 18309 32367 18343
rect 32416 18340 32444 18380
rect 33594 18340 33600 18352
rect 32416 18312 33600 18340
rect 32309 18303 32367 18309
rect 33594 18300 33600 18312
rect 33652 18340 33658 18352
rect 34422 18340 34428 18352
rect 33652 18312 34428 18340
rect 33652 18300 33658 18312
rect 34422 18300 34428 18312
rect 34480 18300 34486 18352
rect 30561 18275 30619 18281
rect 30561 18241 30573 18275
rect 30607 18272 30619 18275
rect 32125 18275 32183 18281
rect 30607 18244 32076 18272
rect 30607 18241 30619 18244
rect 30561 18235 30619 18241
rect 27304 18176 29960 18204
rect 27304 18164 27310 18176
rect 30006 18164 30012 18216
rect 30064 18204 30070 18216
rect 30745 18207 30803 18213
rect 30745 18204 30757 18207
rect 30064 18176 30757 18204
rect 30064 18164 30070 18176
rect 30745 18173 30757 18176
rect 30791 18173 30803 18207
rect 32048 18204 32076 18244
rect 32125 18241 32137 18275
rect 32171 18272 32183 18275
rect 32398 18272 32404 18284
rect 32171 18244 32404 18272
rect 32171 18241 32183 18244
rect 32125 18235 32183 18241
rect 32398 18232 32404 18244
rect 32456 18232 32462 18284
rect 33778 18232 33784 18284
rect 33836 18272 33842 18284
rect 35434 18272 35440 18284
rect 33836 18244 35440 18272
rect 33836 18232 33842 18244
rect 35434 18232 35440 18244
rect 35492 18232 35498 18284
rect 36446 18232 36452 18284
rect 36504 18272 36510 18284
rect 38010 18272 38016 18284
rect 36504 18244 38016 18272
rect 36504 18232 36510 18244
rect 38010 18232 38016 18244
rect 38068 18272 38074 18284
rect 38197 18275 38255 18281
rect 38197 18272 38209 18275
rect 38068 18244 38209 18272
rect 38068 18232 38074 18244
rect 38197 18241 38209 18244
rect 38243 18241 38255 18275
rect 38197 18235 38255 18241
rect 38286 18232 38292 18284
rect 38344 18272 38350 18284
rect 38381 18275 38439 18281
rect 38381 18272 38393 18275
rect 38344 18244 38393 18272
rect 38344 18232 38350 18244
rect 38381 18241 38393 18244
rect 38427 18241 38439 18275
rect 38381 18235 38439 18241
rect 38562 18232 38568 18284
rect 38620 18232 38626 18284
rect 34514 18204 34520 18216
rect 32048 18176 34520 18204
rect 30745 18167 30803 18173
rect 34514 18164 34520 18176
rect 34572 18164 34578 18216
rect 36170 18164 36176 18216
rect 36228 18204 36234 18216
rect 38473 18207 38531 18213
rect 38473 18204 38485 18207
rect 36228 18176 38485 18204
rect 36228 18164 36234 18176
rect 38473 18173 38485 18176
rect 38519 18173 38531 18207
rect 38473 18167 38531 18173
rect 39301 18207 39359 18213
rect 39301 18173 39313 18207
rect 39347 18204 39359 18207
rect 39390 18204 39396 18216
rect 39347 18176 39396 18204
rect 39347 18173 39359 18176
rect 39301 18167 39359 18173
rect 39390 18164 39396 18176
rect 39448 18164 39454 18216
rect 39666 18164 39672 18216
rect 39724 18164 39730 18216
rect 29362 18136 29368 18148
rect 26344 18108 29368 18136
rect 29362 18096 29368 18108
rect 29420 18136 29426 18148
rect 30377 18139 30435 18145
rect 30377 18136 30389 18139
rect 29420 18108 30389 18136
rect 29420 18096 29426 18108
rect 30377 18105 30389 18108
rect 30423 18136 30435 18139
rect 33134 18136 33140 18148
rect 30423 18108 33140 18136
rect 30423 18105 30435 18108
rect 30377 18099 30435 18105
rect 33134 18096 33140 18108
rect 33192 18096 33198 18148
rect 34054 18136 34060 18148
rect 33862 18108 34060 18136
rect 18656 18040 22232 18068
rect 18656 18028 18662 18040
rect 22370 18028 22376 18080
rect 22428 18068 22434 18080
rect 22649 18071 22707 18077
rect 22649 18068 22661 18071
rect 22428 18040 22661 18068
rect 22428 18028 22434 18040
rect 22649 18037 22661 18040
rect 22695 18037 22707 18071
rect 22649 18031 22707 18037
rect 23842 18028 23848 18080
rect 23900 18068 23906 18080
rect 24213 18071 24271 18077
rect 24213 18068 24225 18071
rect 23900 18040 24225 18068
rect 23900 18028 23906 18040
rect 24213 18037 24225 18040
rect 24259 18037 24271 18071
rect 24213 18031 24271 18037
rect 26418 18028 26424 18080
rect 26476 18068 26482 18080
rect 26970 18068 26976 18080
rect 26476 18040 26976 18068
rect 26476 18028 26482 18040
rect 26970 18028 26976 18040
rect 27028 18028 27034 18080
rect 27614 18028 27620 18080
rect 27672 18068 27678 18080
rect 27801 18071 27859 18077
rect 27801 18068 27813 18071
rect 27672 18040 27813 18068
rect 27672 18028 27678 18040
rect 27801 18037 27813 18040
rect 27847 18068 27859 18071
rect 27982 18068 27988 18080
rect 27847 18040 27988 18068
rect 27847 18037 27859 18040
rect 27801 18031 27859 18037
rect 27982 18028 27988 18040
rect 28040 18028 28046 18080
rect 31478 18028 31484 18080
rect 31536 18068 31542 18080
rect 32122 18068 32128 18080
rect 31536 18040 32128 18068
rect 31536 18028 31542 18040
rect 32122 18028 32128 18040
rect 32180 18028 32186 18080
rect 32493 18071 32551 18077
rect 32493 18037 32505 18071
rect 32539 18068 32551 18071
rect 33862 18068 33890 18108
rect 34054 18096 34060 18108
rect 34112 18096 34118 18148
rect 37458 18096 37464 18148
rect 37516 18136 37522 18148
rect 38562 18136 38568 18148
rect 37516 18108 38568 18136
rect 37516 18096 37522 18108
rect 38562 18096 38568 18108
rect 38620 18136 38626 18148
rect 38657 18139 38715 18145
rect 38657 18136 38669 18139
rect 38620 18108 38669 18136
rect 38620 18096 38626 18108
rect 38657 18105 38669 18108
rect 38703 18105 38715 18139
rect 38657 18099 38715 18105
rect 32539 18040 33890 18068
rect 32539 18037 32551 18040
rect 32493 18031 32551 18037
rect 38746 18028 38752 18080
rect 38804 18068 38810 18080
rect 38933 18071 38991 18077
rect 38933 18068 38945 18071
rect 38804 18040 38945 18068
rect 38804 18028 38810 18040
rect 38933 18037 38945 18040
rect 38979 18037 38991 18071
rect 38933 18031 38991 18037
rect 1104 17978 40572 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 40572 17978
rect 1104 17904 40572 17926
rect 12802 17824 12808 17876
rect 12860 17824 12866 17876
rect 13446 17824 13452 17876
rect 13504 17864 13510 17876
rect 13504 17836 16528 17864
rect 13504 17824 13510 17836
rect 9582 17756 9588 17808
rect 9640 17796 9646 17808
rect 16500 17796 16528 17836
rect 16574 17824 16580 17876
rect 16632 17824 16638 17876
rect 17034 17824 17040 17876
rect 17092 17824 17098 17876
rect 18046 17824 18052 17876
rect 18104 17864 18110 17876
rect 18417 17867 18475 17873
rect 18417 17864 18429 17867
rect 18104 17836 18429 17864
rect 18104 17824 18110 17836
rect 18417 17833 18429 17836
rect 18463 17833 18475 17867
rect 18417 17827 18475 17833
rect 18892 17836 19932 17864
rect 18892 17796 18920 17836
rect 9640 17768 13492 17796
rect 16500 17768 18920 17796
rect 9640 17756 9646 17768
rect 4433 17731 4491 17737
rect 4433 17697 4445 17731
rect 4479 17728 4491 17731
rect 4614 17728 4620 17740
rect 4479 17700 4620 17728
rect 4479 17697 4491 17700
rect 4433 17691 4491 17697
rect 4614 17688 4620 17700
rect 4672 17688 4678 17740
rect 5258 17688 5264 17740
rect 5316 17688 5322 17740
rect 8018 17688 8024 17740
rect 8076 17728 8082 17740
rect 9401 17731 9459 17737
rect 9401 17728 9413 17731
rect 8076 17700 9413 17728
rect 8076 17688 8082 17700
rect 9401 17697 9413 17700
rect 9447 17728 9459 17731
rect 9447 17700 9904 17728
rect 9447 17697 9459 17700
rect 9401 17691 9459 17697
rect 7282 17620 7288 17672
rect 7340 17660 7346 17672
rect 7377 17663 7435 17669
rect 7377 17660 7389 17663
rect 7340 17632 7389 17660
rect 7340 17620 7346 17632
rect 7377 17629 7389 17632
rect 7423 17629 7435 17663
rect 7377 17623 7435 17629
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17629 8631 17663
rect 8573 17623 8631 17629
rect 3142 17552 3148 17604
rect 3200 17592 3206 17604
rect 4157 17595 4215 17601
rect 3200 17564 3924 17592
rect 3200 17552 3206 17564
rect 2774 17484 2780 17536
rect 2832 17524 2838 17536
rect 3789 17527 3847 17533
rect 3789 17524 3801 17527
rect 2832 17496 3801 17524
rect 2832 17484 2838 17496
rect 3789 17493 3801 17496
rect 3835 17493 3847 17527
rect 3896 17524 3924 17564
rect 4157 17561 4169 17595
rect 4203 17592 4215 17595
rect 4617 17595 4675 17601
rect 4617 17592 4629 17595
rect 4203 17564 4629 17592
rect 4203 17561 4215 17564
rect 4157 17555 4215 17561
rect 4617 17561 4629 17564
rect 4663 17561 4675 17595
rect 4617 17555 4675 17561
rect 7193 17595 7251 17601
rect 7193 17561 7205 17595
rect 7239 17592 7251 17595
rect 7466 17592 7472 17604
rect 7239 17564 7472 17592
rect 7239 17561 7251 17564
rect 7193 17555 7251 17561
rect 7466 17552 7472 17564
rect 7524 17592 7530 17604
rect 8588 17592 8616 17623
rect 8754 17620 8760 17672
rect 8812 17620 8818 17672
rect 9214 17620 9220 17672
rect 9272 17620 9278 17672
rect 9674 17620 9680 17672
rect 9732 17620 9738 17672
rect 9876 17669 9904 17700
rect 10870 17688 10876 17740
rect 10928 17728 10934 17740
rect 12802 17728 12808 17740
rect 10928 17700 12808 17728
rect 10928 17688 10934 17700
rect 12802 17688 12808 17700
rect 12860 17688 12866 17740
rect 13464 17737 13492 17768
rect 18966 17756 18972 17808
rect 19024 17796 19030 17808
rect 19794 17796 19800 17808
rect 19024 17768 19800 17796
rect 19024 17756 19030 17768
rect 19794 17756 19800 17768
rect 19852 17756 19858 17808
rect 13449 17731 13507 17737
rect 13449 17697 13461 17731
rect 13495 17728 13507 17731
rect 19334 17728 19340 17740
rect 13495 17700 19340 17728
rect 13495 17697 13507 17700
rect 13449 17691 13507 17697
rect 19334 17688 19340 17700
rect 19392 17688 19398 17740
rect 19904 17728 19932 17836
rect 23474 17824 23480 17876
rect 23532 17864 23538 17876
rect 23750 17864 23756 17876
rect 23532 17836 23756 17864
rect 23532 17824 23538 17836
rect 23750 17824 23756 17836
rect 23808 17824 23814 17876
rect 24857 17867 24915 17873
rect 24857 17833 24869 17867
rect 24903 17864 24915 17867
rect 26418 17864 26424 17876
rect 24903 17836 26424 17864
rect 24903 17833 24915 17836
rect 24857 17827 24915 17833
rect 26418 17824 26424 17836
rect 26476 17824 26482 17876
rect 26513 17867 26571 17873
rect 26513 17833 26525 17867
rect 26559 17864 26571 17867
rect 26602 17864 26608 17876
rect 26559 17836 26608 17864
rect 26559 17833 26571 17836
rect 26513 17827 26571 17833
rect 26602 17824 26608 17836
rect 26660 17824 26666 17876
rect 28534 17864 28540 17876
rect 28460 17836 28540 17864
rect 22186 17756 22192 17808
rect 22244 17796 22250 17808
rect 22925 17799 22983 17805
rect 22925 17796 22937 17799
rect 22244 17768 22937 17796
rect 22244 17756 22250 17768
rect 22848 17737 22876 17768
rect 22925 17765 22937 17768
rect 22971 17765 22983 17799
rect 28460 17796 28488 17836
rect 28534 17824 28540 17836
rect 28592 17824 28598 17876
rect 28810 17824 28816 17876
rect 28868 17864 28874 17876
rect 32766 17864 32772 17876
rect 28868 17836 32772 17864
rect 28868 17824 28874 17836
rect 32766 17824 32772 17836
rect 32824 17824 32830 17876
rect 32953 17867 33011 17873
rect 32953 17833 32965 17867
rect 32999 17833 33011 17867
rect 32953 17827 33011 17833
rect 22925 17759 22983 17765
rect 24964 17768 28488 17796
rect 21637 17731 21695 17737
rect 21637 17728 21649 17731
rect 19904 17700 21649 17728
rect 21637 17697 21649 17700
rect 21683 17697 21695 17731
rect 21637 17691 21695 17697
rect 22833 17731 22891 17737
rect 22833 17697 22845 17731
rect 22879 17697 22891 17731
rect 24302 17728 24308 17740
rect 22833 17691 22891 17697
rect 23124 17700 24308 17728
rect 9861 17663 9919 17669
rect 9861 17629 9873 17663
rect 9907 17629 9919 17663
rect 9861 17623 9919 17629
rect 9950 17620 9956 17672
rect 10008 17660 10014 17672
rect 10965 17663 11023 17669
rect 10965 17660 10977 17663
rect 10008 17632 10977 17660
rect 10008 17620 10014 17632
rect 10965 17629 10977 17632
rect 11011 17629 11023 17663
rect 10965 17623 11023 17629
rect 11149 17663 11207 17669
rect 11149 17629 11161 17663
rect 11195 17660 11207 17663
rect 13262 17660 13268 17672
rect 11195 17632 13268 17660
rect 11195 17629 11207 17632
rect 11149 17623 11207 17629
rect 13262 17620 13268 17632
rect 13320 17620 13326 17672
rect 16761 17663 16819 17669
rect 16761 17629 16773 17663
rect 16807 17629 16819 17663
rect 16761 17623 16819 17629
rect 16853 17663 16911 17669
rect 16853 17629 16865 17663
rect 16899 17660 16911 17663
rect 16942 17660 16948 17672
rect 16899 17632 16948 17660
rect 16899 17629 16911 17632
rect 16853 17623 16911 17629
rect 7524 17564 9444 17592
rect 7524 17552 7530 17564
rect 9416 17536 9444 17564
rect 12894 17552 12900 17604
rect 12952 17592 12958 17604
rect 13173 17595 13231 17601
rect 13173 17592 13185 17595
rect 12952 17564 13185 17592
rect 12952 17552 12958 17564
rect 13173 17561 13185 17564
rect 13219 17561 13231 17595
rect 13173 17555 13231 17561
rect 4249 17527 4307 17533
rect 4249 17524 4261 17527
rect 3896 17496 4261 17524
rect 3789 17487 3847 17493
rect 4249 17493 4261 17496
rect 4295 17524 4307 17527
rect 5350 17524 5356 17536
rect 4295 17496 5356 17524
rect 4295 17493 4307 17496
rect 4249 17487 4307 17493
rect 5350 17484 5356 17496
rect 5408 17484 5414 17536
rect 7009 17527 7067 17533
rect 7009 17493 7021 17527
rect 7055 17524 7067 17527
rect 7282 17524 7288 17536
rect 7055 17496 7288 17524
rect 7055 17493 7067 17496
rect 7009 17487 7067 17493
rect 7282 17484 7288 17496
rect 7340 17484 7346 17536
rect 8662 17484 8668 17536
rect 8720 17484 8726 17536
rect 8846 17484 8852 17536
rect 8904 17524 8910 17536
rect 9033 17527 9091 17533
rect 9033 17524 9045 17527
rect 8904 17496 9045 17524
rect 8904 17484 8910 17496
rect 9033 17493 9045 17496
rect 9079 17493 9091 17527
rect 9033 17487 9091 17493
rect 9398 17484 9404 17536
rect 9456 17484 9462 17536
rect 9861 17527 9919 17533
rect 9861 17493 9873 17527
rect 9907 17524 9919 17527
rect 10042 17524 10048 17536
rect 9907 17496 10048 17524
rect 9907 17493 9919 17496
rect 9861 17487 9919 17493
rect 10042 17484 10048 17496
rect 10100 17484 10106 17536
rect 11146 17484 11152 17536
rect 11204 17484 11210 17536
rect 13265 17527 13323 17533
rect 13265 17493 13277 17527
rect 13311 17524 13323 17527
rect 14182 17524 14188 17536
rect 13311 17496 14188 17524
rect 13311 17493 13323 17496
rect 13265 17487 13323 17493
rect 14182 17484 14188 17496
rect 14240 17484 14246 17536
rect 16776 17524 16804 17623
rect 16942 17620 16948 17632
rect 17000 17620 17006 17672
rect 18230 17620 18236 17672
rect 18288 17620 18294 17672
rect 18509 17663 18567 17669
rect 18509 17629 18521 17663
rect 18555 17660 18567 17663
rect 20806 17660 20812 17672
rect 18555 17632 20812 17660
rect 18555 17629 18567 17632
rect 18509 17623 18567 17629
rect 20806 17620 20812 17632
rect 20864 17620 20870 17672
rect 21818 17620 21824 17672
rect 21876 17660 21882 17672
rect 22189 17663 22247 17669
rect 22189 17660 22201 17663
rect 21876 17632 22201 17660
rect 21876 17620 21882 17632
rect 22189 17629 22201 17632
rect 22235 17629 22247 17663
rect 22189 17623 22247 17629
rect 22370 17620 22376 17672
rect 22428 17620 22434 17672
rect 22646 17620 22652 17672
rect 22704 17620 22710 17672
rect 23124 17669 23152 17700
rect 24302 17688 24308 17700
rect 24360 17688 24366 17740
rect 24964 17737 24992 17768
rect 24949 17731 25007 17737
rect 24949 17697 24961 17731
rect 24995 17697 25007 17731
rect 24949 17691 25007 17697
rect 26421 17731 26479 17737
rect 26421 17697 26433 17731
rect 26467 17728 26479 17731
rect 28353 17731 28411 17737
rect 28353 17728 28365 17731
rect 26467 17700 28365 17728
rect 26467 17697 26479 17700
rect 26421 17691 26479 17697
rect 28353 17697 28365 17700
rect 28399 17697 28411 17731
rect 28828 17728 28856 17824
rect 30926 17756 30932 17808
rect 30984 17796 30990 17808
rect 31294 17796 31300 17808
rect 30984 17768 31300 17796
rect 30984 17756 30990 17768
rect 31294 17756 31300 17768
rect 31352 17756 31358 17808
rect 31665 17799 31723 17805
rect 31665 17765 31677 17799
rect 31711 17765 31723 17799
rect 32968 17796 32996 17827
rect 34054 17824 34060 17876
rect 34112 17824 34118 17876
rect 38565 17867 38623 17873
rect 38565 17833 38577 17867
rect 38611 17864 38623 17867
rect 39850 17864 39856 17876
rect 38611 17836 39856 17864
rect 38611 17833 38623 17836
rect 38565 17827 38623 17833
rect 39850 17824 39856 17836
rect 39908 17824 39914 17876
rect 33502 17796 33508 17808
rect 32968 17768 33508 17796
rect 31665 17759 31723 17765
rect 31680 17728 31708 17759
rect 33502 17756 33508 17768
rect 33560 17796 33566 17808
rect 33560 17768 34192 17796
rect 33560 17756 33566 17768
rect 28353 17691 28411 17697
rect 28552 17700 28856 17728
rect 31128 17700 31616 17728
rect 31680 17700 32812 17728
rect 28552 17672 28580 17700
rect 23109 17663 23167 17669
rect 23109 17629 23121 17663
rect 23155 17629 23167 17663
rect 23109 17623 23167 17629
rect 23382 17620 23388 17672
rect 23440 17660 23446 17672
rect 23477 17663 23535 17669
rect 23477 17660 23489 17663
rect 23440 17632 23489 17660
rect 23440 17620 23446 17632
rect 23477 17629 23489 17632
rect 23523 17629 23535 17663
rect 23477 17623 23535 17629
rect 23750 17620 23756 17672
rect 23808 17660 23814 17672
rect 24210 17660 24216 17672
rect 23808 17632 24216 17660
rect 23808 17620 23814 17632
rect 24210 17620 24216 17632
rect 24268 17660 24274 17672
rect 24673 17663 24731 17669
rect 24673 17660 24685 17663
rect 24268 17632 24685 17660
rect 24268 17620 24274 17632
rect 24673 17629 24685 17632
rect 24719 17629 24731 17663
rect 24673 17623 24731 17629
rect 26513 17663 26571 17669
rect 26513 17629 26525 17663
rect 26559 17660 26571 17663
rect 26878 17660 26884 17672
rect 26559 17632 26884 17660
rect 26559 17629 26571 17632
rect 26513 17623 26571 17629
rect 26878 17620 26884 17632
rect 26936 17620 26942 17672
rect 28534 17620 28540 17672
rect 28592 17620 28598 17672
rect 28629 17663 28687 17669
rect 28629 17629 28641 17663
rect 28675 17660 28687 17663
rect 28718 17660 28724 17672
rect 28675 17632 28724 17660
rect 28675 17629 28687 17632
rect 28629 17623 28687 17629
rect 28718 17620 28724 17632
rect 28776 17620 28782 17672
rect 28810 17620 28816 17672
rect 28868 17620 28874 17672
rect 28905 17663 28963 17669
rect 28905 17629 28917 17663
rect 28951 17660 28963 17663
rect 29270 17660 29276 17672
rect 28951 17632 29276 17660
rect 28951 17629 28963 17632
rect 28905 17623 28963 17629
rect 29270 17620 29276 17632
rect 29328 17620 29334 17672
rect 31018 17620 31024 17672
rect 31076 17660 31082 17672
rect 31128 17669 31156 17700
rect 31113 17663 31171 17669
rect 31113 17660 31125 17663
rect 31076 17632 31125 17660
rect 31076 17620 31082 17632
rect 31113 17629 31125 17632
rect 31159 17629 31171 17663
rect 31113 17623 31171 17629
rect 31478 17620 31484 17672
rect 31536 17620 31542 17672
rect 17034 17552 17040 17604
rect 17092 17552 17098 17604
rect 18598 17552 18604 17604
rect 18656 17592 18662 17604
rect 19242 17592 19248 17604
rect 18656 17564 19248 17592
rect 18656 17552 18662 17564
rect 19242 17552 19248 17564
rect 19300 17552 19306 17604
rect 23201 17595 23259 17601
rect 23201 17561 23213 17595
rect 23247 17561 23259 17595
rect 23201 17555 23259 17561
rect 23293 17595 23351 17601
rect 23293 17561 23305 17595
rect 23339 17592 23351 17595
rect 23658 17592 23664 17604
rect 23339 17564 23664 17592
rect 23339 17561 23351 17564
rect 23293 17555 23351 17561
rect 18046 17524 18052 17536
rect 16776 17496 18052 17524
rect 18046 17484 18052 17496
rect 18104 17484 18110 17536
rect 18414 17484 18420 17536
rect 18472 17524 18478 17536
rect 19150 17524 19156 17536
rect 18472 17496 19156 17524
rect 18472 17484 18478 17496
rect 19150 17484 19156 17496
rect 19208 17484 19214 17536
rect 23216 17524 23244 17555
rect 23658 17552 23664 17564
rect 23716 17552 23722 17604
rect 24394 17552 24400 17604
rect 24452 17592 24458 17604
rect 26237 17595 26295 17601
rect 26237 17592 26249 17595
rect 24452 17564 26249 17592
rect 24452 17552 24458 17564
rect 26237 17561 26249 17564
rect 26283 17561 26295 17595
rect 26237 17555 26295 17561
rect 27706 17552 27712 17604
rect 27764 17592 27770 17604
rect 28442 17592 28448 17604
rect 27764 17564 28448 17592
rect 27764 17552 27770 17564
rect 28442 17552 28448 17564
rect 28500 17592 28506 17604
rect 29086 17592 29092 17604
rect 28500 17564 29092 17592
rect 28500 17552 28506 17564
rect 29086 17552 29092 17564
rect 29144 17552 29150 17604
rect 31294 17552 31300 17604
rect 31352 17552 31358 17604
rect 31389 17595 31447 17601
rect 31389 17561 31401 17595
rect 31435 17592 31447 17595
rect 31588 17592 31616 17700
rect 31846 17620 31852 17672
rect 31904 17620 31910 17672
rect 32122 17620 32128 17672
rect 32180 17660 32186 17672
rect 32309 17663 32367 17669
rect 32309 17660 32321 17663
rect 32180 17632 32321 17660
rect 32180 17620 32186 17632
rect 32309 17629 32321 17632
rect 32355 17629 32367 17663
rect 32309 17623 32367 17629
rect 32493 17663 32551 17669
rect 32493 17629 32505 17663
rect 32539 17660 32551 17663
rect 32674 17660 32680 17672
rect 32539 17632 32680 17660
rect 32539 17629 32551 17632
rect 32493 17623 32551 17629
rect 32674 17620 32680 17632
rect 32732 17620 32738 17672
rect 32784 17669 32812 17700
rect 33042 17688 33048 17740
rect 33100 17728 33106 17740
rect 34164 17728 34192 17768
rect 36538 17756 36544 17808
rect 36596 17796 36602 17808
rect 38286 17796 38292 17808
rect 36596 17768 38292 17796
rect 36596 17756 36602 17768
rect 38286 17756 38292 17768
rect 38344 17756 38350 17808
rect 37090 17728 37096 17740
rect 33100 17700 33916 17728
rect 34164 17700 34284 17728
rect 33100 17688 33106 17700
rect 32769 17663 32827 17669
rect 32769 17629 32781 17663
rect 32815 17629 32827 17663
rect 32769 17623 32827 17629
rect 32950 17620 32956 17672
rect 33008 17620 33014 17672
rect 33318 17620 33324 17672
rect 33376 17620 33382 17672
rect 33689 17663 33747 17669
rect 33689 17629 33701 17663
rect 33735 17660 33747 17663
rect 33778 17660 33784 17672
rect 33735 17632 33784 17660
rect 33735 17629 33747 17632
rect 33689 17623 33747 17629
rect 33778 17620 33784 17632
rect 33836 17620 33842 17672
rect 33888 17670 33916 17700
rect 33888 17669 33982 17670
rect 33888 17663 34023 17669
rect 33888 17642 33977 17663
rect 33954 17632 33977 17642
rect 33965 17629 33977 17632
rect 34011 17629 34023 17663
rect 33965 17623 34023 17629
rect 34146 17620 34152 17672
rect 34204 17620 34210 17672
rect 34256 17669 34284 17700
rect 36464 17700 37096 17728
rect 34241 17663 34299 17669
rect 34241 17629 34253 17663
rect 34287 17629 34299 17663
rect 34241 17623 34299 17629
rect 34422 17620 34428 17672
rect 34480 17660 34486 17672
rect 34480 17632 34652 17660
rect 34480 17620 34486 17632
rect 32401 17595 32459 17601
rect 32401 17592 32413 17595
rect 31435 17564 31469 17592
rect 31588 17564 32413 17592
rect 31435 17561 31447 17564
rect 31389 17555 31447 17561
rect 32401 17561 32413 17564
rect 32447 17561 32459 17595
rect 32401 17555 32459 17561
rect 23474 17524 23480 17536
rect 23216 17496 23480 17524
rect 23474 17484 23480 17496
rect 23532 17484 23538 17536
rect 24210 17484 24216 17536
rect 24268 17524 24274 17536
rect 24489 17527 24547 17533
rect 24489 17524 24501 17527
rect 24268 17496 24501 17524
rect 24268 17484 24274 17496
rect 24489 17493 24501 17496
rect 24535 17493 24547 17527
rect 24489 17487 24547 17493
rect 26697 17527 26755 17533
rect 26697 17493 26709 17527
rect 26743 17524 26755 17527
rect 27154 17524 27160 17536
rect 26743 17496 27160 17524
rect 26743 17493 26755 17496
rect 26697 17487 26755 17493
rect 27154 17484 27160 17496
rect 27212 17484 27218 17536
rect 27246 17484 27252 17536
rect 27304 17524 27310 17536
rect 31404 17524 31432 17555
rect 33502 17552 33508 17604
rect 33560 17552 33566 17604
rect 33594 17552 33600 17604
rect 33652 17552 33658 17604
rect 34624 17592 34652 17632
rect 36078 17620 36084 17672
rect 36136 17620 36142 17672
rect 36170 17620 36176 17672
rect 36228 17660 36234 17672
rect 36464 17660 36492 17700
rect 37090 17688 37096 17700
rect 37148 17688 37154 17740
rect 38562 17688 38568 17740
rect 38620 17688 38626 17740
rect 36228 17632 36492 17660
rect 36228 17620 36234 17632
rect 36538 17620 36544 17672
rect 36596 17669 36602 17672
rect 36596 17660 36604 17669
rect 38381 17663 38439 17669
rect 38381 17660 38393 17663
rect 36596 17632 36641 17660
rect 36740 17632 38393 17660
rect 36596 17623 36604 17632
rect 36596 17620 36602 17623
rect 36357 17595 36415 17601
rect 36357 17592 36369 17595
rect 34624 17564 36369 17592
rect 36357 17561 36369 17564
rect 36403 17561 36415 17595
rect 36357 17555 36415 17561
rect 36449 17595 36507 17601
rect 36449 17561 36461 17595
rect 36495 17561 36507 17595
rect 36449 17555 36507 17561
rect 31941 17527 31999 17533
rect 31941 17524 31953 17527
rect 27304 17496 31953 17524
rect 27304 17484 27310 17496
rect 31941 17493 31953 17496
rect 31987 17493 31999 17527
rect 31941 17487 31999 17493
rect 32950 17484 32956 17536
rect 33008 17524 33014 17536
rect 33137 17527 33195 17533
rect 33137 17524 33149 17527
rect 33008 17496 33149 17524
rect 33008 17484 33014 17496
rect 33137 17493 33149 17496
rect 33183 17493 33195 17527
rect 33137 17487 33195 17493
rect 33873 17527 33931 17533
rect 33873 17493 33885 17527
rect 33919 17524 33931 17527
rect 34146 17524 34152 17536
rect 33919 17496 34152 17524
rect 33919 17493 33931 17496
rect 33873 17487 33931 17493
rect 34146 17484 34152 17496
rect 34204 17484 34210 17536
rect 34422 17484 34428 17536
rect 34480 17484 34486 17536
rect 34882 17484 34888 17536
rect 34940 17524 34946 17536
rect 36464 17524 36492 17555
rect 36740 17533 36768 17632
rect 38381 17629 38393 17632
rect 38427 17660 38439 17663
rect 38470 17660 38476 17672
rect 38427 17632 38476 17660
rect 38427 17629 38439 17632
rect 38381 17623 38439 17629
rect 38470 17620 38476 17632
rect 38528 17620 38534 17672
rect 37366 17552 37372 17604
rect 37424 17592 37430 17604
rect 38657 17595 38715 17601
rect 38657 17592 38669 17595
rect 37424 17564 38669 17592
rect 37424 17552 37430 17564
rect 38657 17561 38669 17564
rect 38703 17561 38715 17595
rect 38657 17555 38715 17561
rect 34940 17496 36492 17524
rect 36725 17527 36783 17533
rect 34940 17484 34946 17496
rect 36725 17493 36737 17527
rect 36771 17493 36783 17527
rect 36725 17487 36783 17493
rect 38102 17484 38108 17536
rect 38160 17524 38166 17536
rect 38197 17527 38255 17533
rect 38197 17524 38209 17527
rect 38160 17496 38209 17524
rect 38160 17484 38166 17496
rect 38197 17493 38209 17496
rect 38243 17493 38255 17527
rect 38197 17487 38255 17493
rect 1104 17434 40572 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 40572 17434
rect 1104 17360 40572 17382
rect 4249 17323 4307 17329
rect 4249 17289 4261 17323
rect 4295 17320 4307 17323
rect 5258 17320 5264 17332
rect 4295 17292 5264 17320
rect 4295 17289 4307 17292
rect 4249 17283 4307 17289
rect 5258 17280 5264 17292
rect 5316 17280 5322 17332
rect 5350 17280 5356 17332
rect 5408 17320 5414 17332
rect 10965 17323 11023 17329
rect 5408 17292 8156 17320
rect 5408 17280 5414 17292
rect 2774 17212 2780 17264
rect 2832 17212 2838 17264
rect 3786 17212 3792 17264
rect 3844 17212 3850 17264
rect 6546 17212 6552 17264
rect 6604 17252 6610 17264
rect 7374 17252 7380 17264
rect 6604 17224 7380 17252
rect 6604 17212 6610 17224
rect 7374 17212 7380 17224
rect 7432 17212 7438 17264
rect 7834 17252 7840 17264
rect 7576 17224 7840 17252
rect 2498 17144 2504 17196
rect 2556 17144 2562 17196
rect 6914 17144 6920 17196
rect 6972 17184 6978 17196
rect 7101 17187 7159 17193
rect 7101 17184 7113 17187
rect 6972 17156 7113 17184
rect 6972 17144 6978 17156
rect 7101 17153 7113 17156
rect 7147 17153 7159 17187
rect 7101 17147 7159 17153
rect 7285 17187 7343 17193
rect 7285 17153 7297 17187
rect 7331 17184 7343 17187
rect 7466 17184 7472 17196
rect 7331 17156 7472 17184
rect 7331 17153 7343 17156
rect 7285 17147 7343 17153
rect 7466 17144 7472 17156
rect 7524 17144 7530 17196
rect 7576 17193 7604 17224
rect 7834 17212 7840 17224
rect 7892 17212 7898 17264
rect 7561 17187 7619 17193
rect 7561 17153 7573 17187
rect 7607 17153 7619 17187
rect 7561 17147 7619 17153
rect 7745 17187 7803 17193
rect 7745 17153 7757 17187
rect 7791 17184 7803 17187
rect 7929 17187 7987 17193
rect 7929 17184 7941 17187
rect 7791 17156 7941 17184
rect 7791 17153 7803 17156
rect 7745 17147 7803 17153
rect 7929 17153 7941 17156
rect 7975 17184 7987 17187
rect 8018 17184 8024 17196
rect 7975 17156 8024 17184
rect 7975 17153 7987 17156
rect 7929 17147 7987 17153
rect 8018 17144 8024 17156
rect 8076 17144 8082 17196
rect 8128 17193 8156 17292
rect 10965 17289 10977 17323
rect 11011 17320 11023 17323
rect 11238 17320 11244 17332
rect 11011 17292 11244 17320
rect 11011 17289 11023 17292
rect 10965 17283 11023 17289
rect 11238 17280 11244 17292
rect 11296 17280 11302 17332
rect 17402 17280 17408 17332
rect 17460 17320 17466 17332
rect 18414 17320 18420 17332
rect 17460 17292 18420 17320
rect 17460 17280 17466 17292
rect 18414 17280 18420 17292
rect 18472 17280 18478 17332
rect 18506 17280 18512 17332
rect 18564 17320 18570 17332
rect 20622 17320 20628 17332
rect 18564 17292 20628 17320
rect 18564 17280 18570 17292
rect 20622 17280 20628 17292
rect 20680 17280 20686 17332
rect 24394 17280 24400 17332
rect 24452 17280 24458 17332
rect 27246 17320 27252 17332
rect 24596 17292 27252 17320
rect 9398 17212 9404 17264
rect 9456 17252 9462 17264
rect 9769 17255 9827 17261
rect 9769 17252 9781 17255
rect 9456 17224 9781 17252
rect 9456 17212 9462 17224
rect 9769 17221 9781 17224
rect 9815 17252 9827 17255
rect 10873 17255 10931 17261
rect 9815 17224 10640 17252
rect 9815 17221 9827 17224
rect 9769 17215 9827 17221
rect 8113 17187 8171 17193
rect 8113 17153 8125 17187
rect 8159 17153 8171 17187
rect 8113 17147 8171 17153
rect 8662 17144 8668 17196
rect 8720 17184 8726 17196
rect 9585 17187 9643 17193
rect 9585 17184 9597 17187
rect 8720 17156 9597 17184
rect 8720 17144 8726 17156
rect 9585 17153 9597 17156
rect 9631 17153 9643 17187
rect 9585 17147 9643 17153
rect 9861 17187 9919 17193
rect 9861 17153 9873 17187
rect 9907 17184 9919 17187
rect 10612 17184 10640 17224
rect 10873 17221 10885 17255
rect 10919 17252 10931 17255
rect 11054 17252 11060 17264
rect 10919 17224 11060 17252
rect 10919 17221 10931 17224
rect 10873 17215 10931 17221
rect 11054 17212 11060 17224
rect 11112 17212 11118 17264
rect 14001 17255 14059 17261
rect 14001 17221 14013 17255
rect 14047 17252 14059 17255
rect 14642 17252 14648 17264
rect 14047 17224 14648 17252
rect 14047 17221 14059 17224
rect 14001 17215 14059 17221
rect 14642 17212 14648 17224
rect 14700 17212 14706 17264
rect 17770 17252 17776 17264
rect 16960 17224 17776 17252
rect 11793 17187 11851 17193
rect 9907 17156 10548 17184
rect 10612 17156 11192 17184
rect 9907 17153 9919 17156
rect 9861 17147 9919 17153
rect 5442 17076 5448 17128
rect 5500 17116 5506 17128
rect 5994 17116 6000 17128
rect 5500 17088 6000 17116
rect 5500 17076 5506 17088
rect 5994 17076 6000 17088
rect 6052 17076 6058 17128
rect 7193 17119 7251 17125
rect 7193 17085 7205 17119
rect 7239 17116 7251 17119
rect 7650 17116 7656 17128
rect 7239 17088 7656 17116
rect 7239 17085 7251 17088
rect 7193 17079 7251 17085
rect 7650 17076 7656 17088
rect 7708 17076 7714 17128
rect 10520 17057 10548 17156
rect 11057 17119 11115 17125
rect 11057 17085 11069 17119
rect 11103 17085 11115 17119
rect 11164 17116 11192 17156
rect 11793 17153 11805 17187
rect 11839 17184 11851 17187
rect 12526 17184 12532 17196
rect 11839 17156 12532 17184
rect 11839 17153 11851 17156
rect 11793 17147 11851 17153
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 13817 17187 13875 17193
rect 13817 17153 13829 17187
rect 13863 17184 13875 17187
rect 16850 17184 16856 17196
rect 13863 17156 16856 17184
rect 13863 17153 13875 17156
rect 13817 17147 13875 17153
rect 11882 17116 11888 17128
rect 11164 17088 11888 17116
rect 11057 17079 11115 17085
rect 10505 17051 10563 17057
rect 10505 17017 10517 17051
rect 10551 17017 10563 17051
rect 10505 17011 10563 17017
rect 10870 17008 10876 17060
rect 10928 17048 10934 17060
rect 11072 17048 11100 17079
rect 11882 17076 11888 17088
rect 11940 17116 11946 17128
rect 13832 17116 13860 17147
rect 16850 17144 16856 17156
rect 16908 17144 16914 17196
rect 16960 17193 16988 17224
rect 17770 17212 17776 17224
rect 17828 17212 17834 17264
rect 18598 17212 18604 17264
rect 18656 17212 18662 17264
rect 18690 17212 18696 17264
rect 18748 17252 18754 17264
rect 19029 17255 19087 17261
rect 19029 17252 19041 17255
rect 18748 17224 19041 17252
rect 18748 17212 18754 17224
rect 19029 17221 19041 17224
rect 19075 17221 19087 17255
rect 19029 17215 19087 17221
rect 19242 17212 19248 17264
rect 19300 17212 19306 17264
rect 19610 17212 19616 17264
rect 19668 17212 19674 17264
rect 23937 17255 23995 17261
rect 23937 17221 23949 17255
rect 23983 17252 23995 17255
rect 24489 17255 24547 17261
rect 24489 17252 24501 17255
rect 23983 17224 24501 17252
rect 23983 17221 23995 17224
rect 23937 17215 23995 17221
rect 24489 17221 24501 17224
rect 24535 17221 24547 17255
rect 24489 17215 24547 17221
rect 16945 17187 17003 17193
rect 16945 17153 16957 17187
rect 16991 17153 17003 17187
rect 16945 17147 17003 17153
rect 17034 17144 17040 17196
rect 17092 17144 17098 17196
rect 17313 17187 17371 17193
rect 17313 17153 17325 17187
rect 17359 17184 17371 17187
rect 18230 17184 18236 17196
rect 17359 17156 18236 17184
rect 17359 17153 17371 17156
rect 17313 17147 17371 17153
rect 18230 17144 18236 17156
rect 18288 17184 18294 17196
rect 18616 17184 18644 17212
rect 18288 17156 18644 17184
rect 18785 17187 18843 17193
rect 18288 17144 18294 17156
rect 18785 17153 18797 17187
rect 18831 17184 18843 17187
rect 19426 17184 19432 17196
rect 18831 17156 19432 17184
rect 18831 17153 18843 17156
rect 18785 17147 18843 17153
rect 19426 17144 19432 17156
rect 19484 17144 19490 17196
rect 19705 17187 19763 17193
rect 19705 17153 19717 17187
rect 19751 17153 19763 17187
rect 19705 17147 19763 17153
rect 11940 17088 13860 17116
rect 17052 17116 17080 17144
rect 19720 17116 19748 17147
rect 19794 17144 19800 17196
rect 19852 17184 19858 17196
rect 19852 17156 24164 17184
rect 19852 17144 19858 17156
rect 20162 17116 20168 17128
rect 17052 17088 18920 17116
rect 11940 17076 11946 17088
rect 18892 17057 18920 17088
rect 18984 17088 20168 17116
rect 10928 17020 11100 17048
rect 17221 17051 17279 17057
rect 10928 17008 10934 17020
rect 17221 17017 17233 17051
rect 17267 17048 17279 17051
rect 18877 17051 18935 17057
rect 17267 17020 18828 17048
rect 17267 17017 17279 17020
rect 17221 17011 17279 17017
rect 7374 16940 7380 16992
rect 7432 16940 7438 16992
rect 7558 16940 7564 16992
rect 7616 16980 7622 16992
rect 8021 16983 8079 16989
rect 8021 16980 8033 16983
rect 7616 16952 8033 16980
rect 7616 16940 7622 16952
rect 8021 16949 8033 16952
rect 8067 16980 8079 16983
rect 8110 16980 8116 16992
rect 8067 16952 8116 16980
rect 8067 16949 8079 16952
rect 8021 16943 8079 16949
rect 8110 16940 8116 16952
rect 8168 16940 8174 16992
rect 9401 16983 9459 16989
rect 9401 16949 9413 16983
rect 9447 16980 9459 16983
rect 9582 16980 9588 16992
rect 9447 16952 9588 16980
rect 9447 16949 9459 16952
rect 9401 16943 9459 16949
rect 9582 16940 9588 16952
rect 9640 16940 9646 16992
rect 11885 16983 11943 16989
rect 11885 16949 11897 16983
rect 11931 16980 11943 16983
rect 11974 16980 11980 16992
rect 11931 16952 11980 16980
rect 11931 16949 11943 16952
rect 11885 16943 11943 16949
rect 11974 16940 11980 16952
rect 12032 16940 12038 16992
rect 13630 16940 13636 16992
rect 13688 16940 13694 16992
rect 16761 16983 16819 16989
rect 16761 16949 16773 16983
rect 16807 16980 16819 16983
rect 16942 16980 16948 16992
rect 16807 16952 16948 16980
rect 16807 16949 16819 16952
rect 16761 16943 16819 16949
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 18800 16980 18828 17020
rect 18877 17017 18889 17051
rect 18923 17017 18935 17051
rect 18877 17011 18935 17017
rect 18984 16980 19012 17088
rect 20162 17076 20168 17088
rect 20220 17116 20226 17128
rect 22922 17116 22928 17128
rect 20220 17088 22928 17116
rect 20220 17076 20226 17088
rect 22922 17076 22928 17088
rect 22980 17076 22986 17128
rect 23290 17076 23296 17128
rect 23348 17116 23354 17128
rect 24029 17119 24087 17125
rect 24029 17116 24041 17119
rect 23348 17088 24041 17116
rect 23348 17076 23354 17088
rect 24029 17085 24041 17088
rect 24075 17085 24087 17119
rect 24136 17116 24164 17156
rect 24210 17144 24216 17196
rect 24268 17144 24274 17196
rect 24596 17116 24624 17292
rect 27246 17280 27252 17292
rect 27304 17280 27310 17332
rect 27338 17280 27344 17332
rect 27396 17320 27402 17332
rect 27396 17292 28764 17320
rect 27396 17280 27402 17292
rect 25130 17212 25136 17264
rect 25188 17252 25194 17264
rect 28736 17261 28764 17292
rect 28810 17280 28816 17332
rect 28868 17320 28874 17332
rect 28997 17323 29055 17329
rect 28997 17320 29009 17323
rect 28868 17292 29009 17320
rect 28868 17280 28874 17292
rect 28997 17289 29009 17292
rect 29043 17289 29055 17323
rect 28997 17283 29055 17289
rect 33502 17280 33508 17332
rect 33560 17320 33566 17332
rect 33781 17323 33839 17329
rect 33781 17320 33793 17323
rect 33560 17292 33793 17320
rect 33560 17280 33566 17292
rect 33781 17289 33793 17292
rect 33827 17289 33839 17323
rect 33781 17283 33839 17289
rect 38378 17280 38384 17332
rect 38436 17280 38442 17332
rect 28721 17255 28779 17261
rect 25188 17224 27292 17252
rect 25188 17212 25194 17224
rect 24670 17144 24676 17196
rect 24728 17144 24734 17196
rect 25590 17144 25596 17196
rect 25648 17184 25654 17196
rect 25648 17156 27108 17184
rect 25648 17144 25654 17156
rect 24136 17088 24624 17116
rect 24949 17119 25007 17125
rect 24029 17079 24087 17085
rect 24949 17085 24961 17119
rect 24995 17116 25007 17119
rect 25038 17116 25044 17128
rect 24995 17088 25044 17116
rect 24995 17085 25007 17088
rect 24949 17079 25007 17085
rect 20622 17008 20628 17060
rect 20680 17048 20686 17060
rect 24964 17048 24992 17079
rect 25038 17076 25044 17088
rect 25096 17076 25102 17128
rect 26973 17119 27031 17125
rect 26973 17085 26985 17119
rect 27019 17085 27031 17119
rect 27080 17116 27108 17156
rect 27154 17144 27160 17196
rect 27212 17144 27218 17196
rect 27264 17184 27292 17224
rect 27586 17224 28672 17252
rect 27586 17184 27614 17224
rect 27264 17156 27614 17184
rect 28166 17144 28172 17196
rect 28224 17184 28230 17196
rect 28644 17193 28672 17224
rect 28721 17221 28733 17255
rect 28767 17221 28779 17255
rect 28721 17215 28779 17221
rect 32674 17212 32680 17264
rect 32732 17252 32738 17264
rect 32732 17224 33916 17252
rect 32732 17212 32738 17224
rect 28342 17187 28400 17193
rect 28342 17184 28354 17187
rect 28224 17156 28354 17184
rect 28224 17144 28230 17156
rect 28342 17153 28354 17156
rect 28388 17153 28400 17187
rect 28473 17187 28531 17193
rect 28473 17184 28485 17187
rect 28342 17147 28400 17153
rect 28460 17153 28485 17184
rect 28519 17153 28531 17187
rect 28460 17147 28531 17153
rect 28629 17187 28687 17193
rect 28629 17153 28641 17187
rect 28675 17153 28687 17187
rect 28837 17187 28895 17193
rect 28837 17184 28849 17187
rect 28629 17147 28687 17153
rect 28736 17156 28849 17184
rect 27433 17119 27491 17125
rect 27433 17116 27445 17119
rect 27080 17088 27445 17116
rect 26973 17079 27031 17085
rect 27433 17085 27445 17088
rect 27479 17085 27491 17119
rect 27433 17079 27491 17085
rect 27985 17119 28043 17125
rect 27985 17085 27997 17119
rect 28031 17085 28043 17119
rect 27985 17079 28043 17085
rect 25222 17048 25228 17060
rect 20680 17020 24992 17048
rect 25056 17020 25228 17048
rect 20680 17008 20686 17020
rect 18800 16952 19012 16980
rect 19061 16983 19119 16989
rect 19061 16949 19073 16983
rect 19107 16980 19119 16983
rect 19150 16980 19156 16992
rect 19107 16952 19156 16980
rect 19107 16949 19119 16952
rect 19061 16943 19119 16949
rect 19150 16940 19156 16952
rect 19208 16940 19214 16992
rect 19978 16940 19984 16992
rect 20036 16940 20042 16992
rect 22830 16940 22836 16992
rect 22888 16980 22894 16992
rect 23937 16983 23995 16989
rect 23937 16980 23949 16983
rect 22888 16952 23949 16980
rect 22888 16940 22894 16952
rect 23937 16949 23949 16952
rect 23983 16949 23995 16983
rect 23937 16943 23995 16949
rect 24854 16940 24860 16992
rect 24912 16980 24918 16992
rect 25056 16980 25084 17020
rect 25222 17008 25228 17020
rect 25280 17008 25286 17060
rect 26988 17048 27016 17079
rect 27798 17048 27804 17060
rect 26988 17020 27804 17048
rect 27798 17008 27804 17020
rect 27856 17008 27862 17060
rect 24912 16952 25084 16980
rect 28000 16980 28028 17079
rect 28460 17048 28488 17147
rect 28736 17128 28764 17156
rect 28837 17153 28849 17156
rect 28883 17153 28895 17187
rect 28837 17147 28895 17153
rect 30101 17187 30159 17193
rect 30101 17153 30113 17187
rect 30147 17153 30159 17187
rect 30101 17147 30159 17153
rect 30285 17187 30343 17193
rect 30285 17153 30297 17187
rect 30331 17184 30343 17187
rect 31938 17184 31944 17196
rect 30331 17156 31944 17184
rect 30331 17153 30343 17156
rect 30285 17147 30343 17153
rect 28718 17076 28724 17128
rect 28776 17076 28782 17128
rect 28994 17048 29000 17060
rect 28460 17020 29000 17048
rect 28994 17008 29000 17020
rect 29052 17048 29058 17060
rect 30116 17048 30144 17147
rect 31938 17144 31944 17156
rect 31996 17144 32002 17196
rect 32582 17144 32588 17196
rect 32640 17184 32646 17196
rect 33594 17184 33600 17196
rect 32640 17156 33600 17184
rect 32640 17144 32646 17156
rect 33594 17144 33600 17156
rect 33652 17144 33658 17196
rect 33888 17193 33916 17224
rect 34422 17212 34428 17264
rect 34480 17252 34486 17264
rect 37921 17255 37979 17261
rect 37921 17252 37933 17255
rect 34480 17224 37933 17252
rect 34480 17212 34486 17224
rect 37921 17221 37933 17224
rect 37967 17221 37979 17255
rect 37921 17215 37979 17221
rect 33689 17187 33747 17193
rect 33689 17153 33701 17187
rect 33735 17153 33747 17187
rect 33689 17147 33747 17153
rect 33873 17187 33931 17193
rect 33873 17153 33885 17187
rect 33919 17153 33931 17187
rect 33873 17147 33931 17153
rect 30374 17076 30380 17128
rect 30432 17076 30438 17128
rect 33704 17116 33732 17147
rect 34790 17144 34796 17196
rect 34848 17184 34854 17196
rect 35250 17193 35256 17196
rect 35069 17187 35127 17193
rect 35069 17184 35081 17187
rect 34848 17156 35081 17184
rect 34848 17144 34854 17156
rect 35069 17153 35081 17156
rect 35115 17153 35127 17187
rect 35069 17147 35127 17153
rect 35217 17187 35256 17193
rect 35217 17153 35229 17187
rect 35217 17147 35256 17153
rect 35250 17144 35256 17147
rect 35308 17144 35314 17196
rect 35342 17144 35348 17196
rect 35400 17144 35406 17196
rect 35437 17187 35495 17193
rect 35437 17153 35449 17187
rect 35483 17153 35495 17187
rect 35437 17147 35495 17153
rect 35575 17187 35633 17193
rect 35575 17153 35587 17187
rect 35621 17153 35633 17187
rect 35575 17147 35633 17153
rect 35897 17187 35955 17193
rect 35897 17153 35909 17187
rect 35943 17184 35955 17187
rect 35986 17184 35992 17196
rect 35943 17156 35992 17184
rect 35943 17153 35955 17156
rect 35897 17147 35955 17153
rect 33612 17088 33732 17116
rect 33612 17060 33640 17088
rect 29052 17020 30144 17048
rect 29052 17008 29058 17020
rect 33594 17008 33600 17060
rect 33652 17008 33658 17060
rect 35342 17008 35348 17060
rect 35400 17048 35406 17060
rect 35452 17048 35480 17147
rect 35590 17116 35618 17147
rect 35986 17144 35992 17156
rect 36044 17144 36050 17196
rect 38102 17144 38108 17196
rect 38160 17144 38166 17196
rect 38197 17187 38255 17193
rect 38197 17153 38209 17187
rect 38243 17153 38255 17187
rect 38197 17147 38255 17153
rect 36446 17116 36452 17128
rect 35590 17088 36452 17116
rect 36446 17076 36452 17088
rect 36504 17076 36510 17128
rect 37090 17076 37096 17128
rect 37148 17116 37154 17128
rect 38212 17116 38240 17147
rect 37148 17088 38240 17116
rect 37148 17076 37154 17088
rect 36081 17051 36139 17057
rect 36081 17048 36093 17051
rect 35400 17020 36093 17048
rect 35400 17008 35406 17020
rect 36081 17017 36093 17020
rect 36127 17017 36139 17051
rect 36081 17011 36139 17017
rect 28350 16980 28356 16992
rect 28000 16952 28356 16980
rect 24912 16940 24918 16952
rect 28350 16940 28356 16952
rect 28408 16940 28414 16992
rect 29270 16940 29276 16992
rect 29328 16980 29334 16992
rect 29917 16983 29975 16989
rect 29917 16980 29929 16983
rect 29328 16952 29929 16980
rect 29328 16940 29334 16952
rect 29917 16949 29929 16952
rect 29963 16949 29975 16983
rect 29917 16943 29975 16949
rect 35434 16940 35440 16992
rect 35492 16980 35498 16992
rect 35713 16983 35771 16989
rect 35713 16980 35725 16983
rect 35492 16952 35725 16980
rect 35492 16940 35498 16952
rect 35713 16949 35725 16952
rect 35759 16949 35771 16983
rect 35713 16943 35771 16949
rect 37918 16940 37924 16992
rect 37976 16940 37982 16992
rect 1104 16890 40572 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 40572 16890
rect 1104 16816 40572 16838
rect 6546 16736 6552 16788
rect 6604 16736 6610 16788
rect 6914 16736 6920 16788
rect 6972 16776 6978 16788
rect 7282 16776 7288 16788
rect 6972 16748 7288 16776
rect 6972 16736 6978 16748
rect 7282 16736 7288 16748
rect 7340 16736 7346 16788
rect 7650 16736 7656 16788
rect 7708 16776 7714 16788
rect 7837 16779 7895 16785
rect 7837 16776 7849 16779
rect 7708 16748 7849 16776
rect 7708 16736 7714 16748
rect 7837 16745 7849 16748
rect 7883 16745 7895 16779
rect 7837 16739 7895 16745
rect 7006 16668 7012 16720
rect 7064 16668 7070 16720
rect 7101 16711 7159 16717
rect 7101 16677 7113 16711
rect 7147 16677 7159 16711
rect 7101 16671 7159 16677
rect 4798 16600 4804 16652
rect 4856 16600 4862 16652
rect 5077 16643 5135 16649
rect 5077 16609 5089 16643
rect 5123 16640 5135 16643
rect 6086 16640 6092 16652
rect 5123 16612 6092 16640
rect 5123 16609 5135 16612
rect 5077 16603 5135 16609
rect 6086 16600 6092 16612
rect 6144 16600 6150 16652
rect 6822 16600 6828 16652
rect 6880 16640 6886 16652
rect 7116 16640 7144 16671
rect 6880 16612 7144 16640
rect 6880 16600 6886 16612
rect 7558 16600 7564 16652
rect 7616 16640 7622 16652
rect 7653 16643 7711 16649
rect 7653 16640 7665 16643
rect 7616 16612 7665 16640
rect 7616 16600 7622 16612
rect 7653 16609 7665 16612
rect 7699 16609 7711 16643
rect 7852 16640 7880 16739
rect 8202 16736 8208 16788
rect 8260 16736 8266 16788
rect 12342 16736 12348 16788
rect 12400 16776 12406 16788
rect 12989 16779 13047 16785
rect 12989 16776 13001 16779
rect 12400 16748 13001 16776
rect 12400 16736 12406 16748
rect 12989 16745 13001 16748
rect 13035 16745 13047 16779
rect 12989 16739 13047 16745
rect 16390 16736 16396 16788
rect 16448 16776 16454 16788
rect 19058 16776 19064 16788
rect 16448 16748 19064 16776
rect 16448 16736 16454 16748
rect 19058 16736 19064 16748
rect 19116 16736 19122 16788
rect 21177 16779 21235 16785
rect 21177 16745 21189 16779
rect 21223 16776 21235 16779
rect 21269 16779 21327 16785
rect 21269 16776 21281 16779
rect 21223 16748 21281 16776
rect 21223 16745 21235 16748
rect 21177 16739 21235 16745
rect 21269 16745 21281 16748
rect 21315 16745 21327 16779
rect 22281 16779 22339 16785
rect 22281 16776 22293 16779
rect 21269 16739 21327 16745
rect 21376 16748 22293 16776
rect 7926 16668 7932 16720
rect 7984 16708 7990 16720
rect 12158 16708 12164 16720
rect 7984 16680 9444 16708
rect 7984 16668 7990 16680
rect 7852 16612 8064 16640
rect 7653 16603 7711 16609
rect 6733 16575 6791 16581
rect 6733 16541 6745 16575
rect 6779 16572 6791 16575
rect 7282 16572 7288 16584
rect 6779 16544 7288 16572
rect 6779 16541 6791 16544
rect 6733 16535 6791 16541
rect 7282 16532 7288 16544
rect 7340 16532 7346 16584
rect 8036 16581 8064 16612
rect 8110 16600 8116 16652
rect 8168 16600 8174 16652
rect 9416 16649 9444 16680
rect 11348 16680 12164 16708
rect 9401 16643 9459 16649
rect 9401 16609 9413 16643
rect 9447 16609 9459 16643
rect 9401 16603 9459 16609
rect 9490 16600 9496 16652
rect 9548 16600 9554 16652
rect 10502 16600 10508 16652
rect 10560 16600 10566 16652
rect 11348 16649 11376 16680
rect 12158 16668 12164 16680
rect 12216 16668 12222 16720
rect 17402 16708 17408 16720
rect 12268 16680 13032 16708
rect 11333 16643 11391 16649
rect 11333 16609 11345 16643
rect 11379 16609 11391 16643
rect 11333 16603 11391 16609
rect 11698 16600 11704 16652
rect 11756 16600 11762 16652
rect 12268 16640 12296 16680
rect 13004 16652 13032 16680
rect 16868 16680 17408 16708
rect 11900 16612 12296 16640
rect 7929 16575 7987 16581
rect 7929 16541 7941 16575
rect 7975 16541 7987 16575
rect 7929 16535 7987 16541
rect 8021 16575 8079 16581
rect 8021 16541 8033 16575
rect 8067 16541 8079 16575
rect 8021 16535 8079 16541
rect 10229 16575 10287 16581
rect 10229 16541 10241 16575
rect 10275 16572 10287 16575
rect 11149 16575 11207 16581
rect 11149 16572 11161 16575
rect 10275 16544 11161 16572
rect 10275 16541 10287 16544
rect 10229 16535 10287 16541
rect 11149 16541 11161 16544
rect 11195 16572 11207 16575
rect 11238 16572 11244 16584
rect 11195 16544 11244 16572
rect 11195 16541 11207 16544
rect 11149 16535 11207 16541
rect 3786 16464 3792 16516
rect 3844 16504 3850 16516
rect 6825 16507 6883 16513
rect 3844 16476 5566 16504
rect 3844 16464 3850 16476
rect 6825 16473 6837 16507
rect 6871 16504 6883 16507
rect 6914 16504 6920 16516
rect 6871 16476 6920 16504
rect 6871 16473 6883 16476
rect 6825 16467 6883 16473
rect 6914 16464 6920 16476
rect 6972 16464 6978 16516
rect 7009 16507 7067 16513
rect 7009 16473 7021 16507
rect 7055 16504 7067 16507
rect 7374 16504 7380 16516
rect 7055 16476 7380 16504
rect 7055 16473 7067 16476
rect 7009 16467 7067 16473
rect 7374 16464 7380 16476
rect 7432 16504 7438 16516
rect 7469 16507 7527 16513
rect 7469 16504 7481 16507
rect 7432 16476 7481 16504
rect 7432 16464 7438 16476
rect 7469 16473 7481 16476
rect 7515 16473 7527 16507
rect 7944 16504 7972 16535
rect 11238 16532 11244 16544
rect 11296 16572 11302 16584
rect 11900 16581 11928 16612
rect 12986 16600 12992 16652
rect 13044 16640 13050 16652
rect 13725 16643 13783 16649
rect 13044 16612 13676 16640
rect 13044 16600 13050 16612
rect 11885 16575 11943 16581
rect 11885 16572 11897 16575
rect 11296 16544 11897 16572
rect 11296 16532 11302 16544
rect 11885 16541 11897 16544
rect 11931 16541 11943 16575
rect 12406 16572 12756 16574
rect 11885 16535 11943 16541
rect 11992 16546 13584 16572
rect 11992 16544 12434 16546
rect 12728 16544 13584 16546
rect 8202 16504 8208 16516
rect 7944 16476 8208 16504
rect 7469 16467 7527 16473
rect 8202 16464 8208 16476
rect 8260 16464 8266 16516
rect 9309 16507 9367 16513
rect 9309 16473 9321 16507
rect 9355 16504 9367 16507
rect 10321 16507 10379 16513
rect 9355 16476 9904 16504
rect 9355 16473 9367 16476
rect 9309 16467 9367 16473
rect 7282 16445 7288 16448
rect 7269 16439 7288 16445
rect 7269 16405 7281 16439
rect 7269 16399 7288 16405
rect 7282 16396 7288 16399
rect 7340 16396 7346 16448
rect 7650 16396 7656 16448
rect 7708 16396 7714 16448
rect 8386 16396 8392 16448
rect 8444 16396 8450 16448
rect 8938 16396 8944 16448
rect 8996 16396 9002 16448
rect 9876 16445 9904 16476
rect 10321 16473 10333 16507
rect 10367 16504 10379 16507
rect 11054 16504 11060 16516
rect 10367 16476 11060 16504
rect 10367 16473 10379 16476
rect 10321 16467 10379 16473
rect 11054 16464 11060 16476
rect 11112 16504 11118 16516
rect 11793 16507 11851 16513
rect 11793 16504 11805 16507
rect 11112 16476 11805 16504
rect 11112 16464 11118 16476
rect 11793 16473 11805 16476
rect 11839 16504 11851 16507
rect 11992 16504 12020 16544
rect 11839 16476 12020 16504
rect 11839 16473 11851 16476
rect 11793 16467 11851 16473
rect 12158 16464 12164 16516
rect 12216 16504 12222 16516
rect 12437 16507 12495 16513
rect 12437 16504 12449 16507
rect 12216 16476 12449 16504
rect 12216 16464 12222 16476
rect 12437 16473 12449 16476
rect 12483 16473 12495 16507
rect 12437 16467 12495 16473
rect 12713 16507 12771 16513
rect 12713 16473 12725 16507
rect 12759 16504 12771 16507
rect 12759 16476 13216 16504
rect 12759 16473 12771 16476
rect 12713 16467 12771 16473
rect 9861 16439 9919 16445
rect 9861 16405 9873 16439
rect 9907 16405 9919 16439
rect 9861 16399 9919 16405
rect 10686 16396 10692 16448
rect 10744 16396 10750 16448
rect 11698 16396 11704 16448
rect 11756 16436 11762 16448
rect 12253 16439 12311 16445
rect 12253 16436 12265 16439
rect 11756 16408 12265 16436
rect 11756 16396 11762 16408
rect 12253 16405 12265 16408
rect 12299 16405 12311 16439
rect 12253 16399 12311 16405
rect 12526 16396 12532 16448
rect 12584 16396 12590 16448
rect 13188 16445 13216 16476
rect 13556 16445 13584 16544
rect 13648 16513 13676 16612
rect 13725 16609 13737 16643
rect 13771 16640 13783 16643
rect 13814 16640 13820 16652
rect 13771 16612 13820 16640
rect 13771 16609 13783 16612
rect 13725 16603 13783 16609
rect 13814 16600 13820 16612
rect 13872 16640 13878 16652
rect 13998 16640 14004 16652
rect 13872 16612 14004 16640
rect 13872 16600 13878 16612
rect 13998 16600 14004 16612
rect 14056 16600 14062 16652
rect 14366 16600 14372 16652
rect 14424 16600 14430 16652
rect 14476 16612 14872 16640
rect 14476 16584 14504 16612
rect 14090 16532 14096 16584
rect 14148 16572 14154 16584
rect 14458 16572 14464 16584
rect 14148 16544 14464 16572
rect 14148 16532 14154 16544
rect 14458 16532 14464 16544
rect 14516 16532 14522 16584
rect 14550 16532 14556 16584
rect 14608 16532 14614 16584
rect 14844 16581 14872 16612
rect 15010 16600 15016 16652
rect 15068 16600 15074 16652
rect 16868 16640 16896 16680
rect 17402 16668 17408 16680
rect 17460 16668 17466 16720
rect 18046 16668 18052 16720
rect 18104 16708 18110 16720
rect 21376 16708 21404 16748
rect 22281 16745 22293 16748
rect 22327 16745 22339 16779
rect 22281 16739 22339 16745
rect 22741 16779 22799 16785
rect 22741 16745 22753 16779
rect 22787 16776 22799 16779
rect 22787 16748 22876 16776
rect 22787 16745 22799 16748
rect 22741 16739 22799 16745
rect 18104 16680 21404 16708
rect 21637 16711 21695 16717
rect 18104 16668 18110 16680
rect 21637 16677 21649 16711
rect 21683 16708 21695 16711
rect 22646 16708 22652 16720
rect 21683 16680 22652 16708
rect 21683 16677 21695 16680
rect 21637 16671 21695 16677
rect 22646 16668 22652 16680
rect 22704 16668 22710 16720
rect 18064 16640 18092 16668
rect 16776 16612 16896 16640
rect 17052 16612 18092 16640
rect 16776 16581 16804 16612
rect 17052 16581 17080 16612
rect 19426 16600 19432 16652
rect 19484 16640 19490 16652
rect 19794 16640 19800 16652
rect 19484 16612 19800 16640
rect 19484 16600 19490 16612
rect 19794 16600 19800 16612
rect 19852 16640 19858 16652
rect 20438 16640 20444 16652
rect 19852 16612 20444 16640
rect 19852 16600 19858 16612
rect 20438 16600 20444 16612
rect 20496 16640 20502 16652
rect 20533 16643 20591 16649
rect 20533 16640 20545 16643
rect 20496 16612 20545 16640
rect 20496 16600 20502 16612
rect 20533 16609 20545 16612
rect 20579 16609 20591 16643
rect 20533 16603 20591 16609
rect 20622 16600 20628 16652
rect 20680 16640 20686 16652
rect 21361 16643 21419 16649
rect 21361 16640 21373 16643
rect 20680 16612 21373 16640
rect 20680 16600 20686 16612
rect 21361 16609 21373 16612
rect 21407 16609 21419 16643
rect 21361 16603 21419 16609
rect 22186 16600 22192 16652
rect 22244 16640 22250 16652
rect 22373 16643 22431 16649
rect 22373 16640 22385 16643
rect 22244 16612 22385 16640
rect 22244 16600 22250 16612
rect 22373 16609 22385 16612
rect 22419 16609 22431 16643
rect 22373 16603 22431 16609
rect 14645 16575 14703 16581
rect 14645 16541 14657 16575
rect 14691 16541 14703 16575
rect 14645 16535 14703 16541
rect 14829 16575 14887 16581
rect 14829 16541 14841 16575
rect 14875 16541 14887 16575
rect 14829 16535 14887 16541
rect 16761 16575 16819 16581
rect 16761 16541 16773 16575
rect 16807 16541 16819 16575
rect 16761 16535 16819 16541
rect 16853 16575 16911 16581
rect 16853 16541 16865 16575
rect 16899 16572 16911 16575
rect 17037 16575 17095 16581
rect 16899 16544 16988 16572
rect 16899 16541 16911 16544
rect 16853 16535 16911 16541
rect 13633 16507 13691 16513
rect 13633 16473 13645 16507
rect 13679 16504 13691 16507
rect 14568 16504 14596 16532
rect 13679 16476 14596 16504
rect 13679 16473 13691 16476
rect 13633 16467 13691 16473
rect 13173 16439 13231 16445
rect 13173 16405 13185 16439
rect 13219 16405 13231 16439
rect 13173 16399 13231 16405
rect 13541 16439 13599 16445
rect 13541 16405 13553 16439
rect 13587 16436 13599 16439
rect 13722 16436 13728 16448
rect 13587 16408 13728 16436
rect 13587 16405 13599 16408
rect 13541 16399 13599 16405
rect 13722 16396 13728 16408
rect 13780 16396 13786 16448
rect 13814 16396 13820 16448
rect 13872 16436 13878 16448
rect 14182 16436 14188 16448
rect 13872 16408 14188 16436
rect 13872 16396 13878 16408
rect 14182 16396 14188 16408
rect 14240 16436 14246 16448
rect 14660 16436 14688 16535
rect 14240 16408 14688 16436
rect 16577 16439 16635 16445
rect 14240 16396 14246 16408
rect 16577 16405 16589 16439
rect 16623 16436 16635 16439
rect 16666 16436 16672 16448
rect 16623 16408 16672 16436
rect 16623 16405 16635 16408
rect 16577 16399 16635 16405
rect 16666 16396 16672 16408
rect 16724 16396 16730 16448
rect 16960 16436 16988 16544
rect 17037 16541 17049 16575
rect 17083 16541 17095 16575
rect 17037 16535 17095 16541
rect 17129 16575 17187 16581
rect 17129 16541 17141 16575
rect 17175 16572 17187 16575
rect 17218 16572 17224 16584
rect 17175 16544 17224 16572
rect 17175 16541 17187 16544
rect 17129 16535 17187 16541
rect 17218 16532 17224 16544
rect 17276 16572 17282 16584
rect 18138 16572 18144 16584
rect 17276 16544 18144 16572
rect 17276 16532 17282 16544
rect 18138 16532 18144 16544
rect 18196 16532 18202 16584
rect 20993 16575 21051 16581
rect 20993 16541 21005 16575
rect 21039 16572 21051 16575
rect 21174 16572 21180 16584
rect 21039 16544 21180 16572
rect 21039 16541 21051 16544
rect 20993 16535 21051 16541
rect 21174 16532 21180 16544
rect 21232 16532 21238 16584
rect 21269 16575 21327 16581
rect 21269 16541 21281 16575
rect 21315 16541 21327 16575
rect 21269 16535 21327 16541
rect 20714 16513 20720 16516
rect 20691 16507 20720 16513
rect 20691 16473 20703 16507
rect 20691 16467 20720 16473
rect 20714 16464 20720 16467
rect 20772 16464 20778 16516
rect 20806 16464 20812 16516
rect 20864 16464 20870 16516
rect 20898 16464 20904 16516
rect 20956 16464 20962 16516
rect 19610 16436 19616 16448
rect 16960 16408 19616 16436
rect 19610 16396 19616 16408
rect 19668 16396 19674 16448
rect 19978 16396 19984 16448
rect 20036 16436 20042 16448
rect 21284 16436 21312 16535
rect 21818 16532 21824 16584
rect 21876 16572 21882 16584
rect 22557 16575 22615 16581
rect 21876 16544 22508 16572
rect 21876 16532 21882 16544
rect 22278 16464 22284 16516
rect 22336 16464 22342 16516
rect 22480 16504 22508 16544
rect 22557 16541 22569 16575
rect 22603 16572 22615 16575
rect 22646 16572 22652 16584
rect 22603 16544 22652 16572
rect 22603 16541 22615 16544
rect 22557 16535 22615 16541
rect 22646 16532 22652 16544
rect 22704 16532 22710 16584
rect 22848 16581 22876 16748
rect 22922 16736 22928 16788
rect 22980 16736 22986 16788
rect 26694 16736 26700 16788
rect 26752 16776 26758 16788
rect 26789 16779 26847 16785
rect 26789 16776 26801 16779
rect 26752 16748 26801 16776
rect 26752 16736 26758 16748
rect 26789 16745 26801 16748
rect 26835 16745 26847 16779
rect 26789 16739 26847 16745
rect 28074 16736 28080 16788
rect 28132 16776 28138 16788
rect 28169 16779 28227 16785
rect 28169 16776 28181 16779
rect 28132 16748 28181 16776
rect 28132 16736 28138 16748
rect 28169 16745 28181 16748
rect 28215 16745 28227 16779
rect 28169 16739 28227 16745
rect 28258 16736 28264 16788
rect 28316 16776 28322 16788
rect 28316 16748 28764 16776
rect 28316 16736 28322 16748
rect 26513 16711 26571 16717
rect 26513 16677 26525 16711
rect 26559 16708 26571 16711
rect 28626 16708 28632 16720
rect 26559 16680 28632 16708
rect 26559 16677 26571 16680
rect 26513 16671 26571 16677
rect 28626 16668 28632 16680
rect 28684 16668 28690 16720
rect 28736 16708 28764 16748
rect 29086 16736 29092 16788
rect 29144 16776 29150 16788
rect 35342 16776 35348 16788
rect 29144 16748 35348 16776
rect 29144 16736 29150 16748
rect 35342 16736 35348 16748
rect 35400 16736 35406 16788
rect 36446 16736 36452 16788
rect 36504 16776 36510 16788
rect 36814 16776 36820 16788
rect 36504 16748 36820 16776
rect 36504 16736 36510 16748
rect 36814 16736 36820 16748
rect 36872 16736 36878 16788
rect 38286 16736 38292 16788
rect 38344 16776 38350 16788
rect 38381 16779 38439 16785
rect 38381 16776 38393 16779
rect 38344 16748 38393 16776
rect 38344 16736 38350 16748
rect 38381 16745 38393 16748
rect 38427 16745 38439 16779
rect 38381 16739 38439 16745
rect 28736 16680 28948 16708
rect 22922 16600 22928 16652
rect 22980 16600 22986 16652
rect 25682 16600 25688 16652
rect 25740 16600 25746 16652
rect 25774 16600 25780 16652
rect 25832 16640 25838 16652
rect 26329 16643 26387 16649
rect 26329 16640 26341 16643
rect 25832 16612 26341 16640
rect 25832 16600 25838 16612
rect 26329 16609 26341 16612
rect 26375 16609 26387 16643
rect 26329 16603 26387 16609
rect 28166 16600 28172 16652
rect 28224 16640 28230 16652
rect 28920 16640 28948 16680
rect 32950 16668 32956 16720
rect 33008 16708 33014 16720
rect 36906 16708 36912 16720
rect 33008 16680 36912 16708
rect 33008 16668 33014 16680
rect 36906 16668 36912 16680
rect 36964 16668 36970 16720
rect 37093 16711 37151 16717
rect 37093 16677 37105 16711
rect 37139 16708 37151 16711
rect 37366 16708 37372 16720
rect 37139 16680 37372 16708
rect 37139 16677 37151 16680
rect 37093 16671 37151 16677
rect 37366 16668 37372 16680
rect 37424 16668 37430 16720
rect 36814 16640 36820 16652
rect 28224 16612 28856 16640
rect 28920 16612 28994 16640
rect 28224 16600 28230 16612
rect 22833 16575 22891 16581
rect 22833 16541 22845 16575
rect 22879 16541 22891 16575
rect 24486 16572 24492 16584
rect 22833 16535 22891 16541
rect 23768 16544 24492 16572
rect 23768 16504 23796 16544
rect 24486 16532 24492 16544
rect 24544 16572 24550 16584
rect 25317 16575 25375 16581
rect 25317 16572 25329 16575
rect 24544 16544 25329 16572
rect 24544 16532 24550 16544
rect 25317 16541 25329 16544
rect 25363 16541 25375 16575
rect 25317 16535 25375 16541
rect 22480 16476 23796 16504
rect 24762 16464 24768 16516
rect 24820 16464 24826 16516
rect 25332 16504 25360 16535
rect 25498 16532 25504 16584
rect 25556 16532 25562 16584
rect 25792 16571 25820 16600
rect 25777 16565 25835 16571
rect 25777 16531 25789 16565
rect 25823 16531 25835 16565
rect 26050 16532 26056 16584
rect 26108 16532 26114 16584
rect 26237 16575 26295 16581
rect 26237 16541 26249 16575
rect 26283 16541 26295 16575
rect 26237 16535 26295 16541
rect 25777 16525 25835 16531
rect 25590 16504 25596 16516
rect 25332 16476 25596 16504
rect 25590 16464 25596 16476
rect 25648 16464 25654 16516
rect 26252 16504 26280 16535
rect 26418 16532 26424 16584
rect 26476 16532 26482 16584
rect 28074 16532 28080 16584
rect 28132 16572 28138 16584
rect 28348 16575 28406 16581
rect 28132 16566 28212 16572
rect 28348 16566 28360 16575
rect 28132 16544 28360 16566
rect 28132 16532 28138 16544
rect 28184 16541 28360 16544
rect 28394 16541 28406 16575
rect 28184 16538 28406 16541
rect 28348 16535 28406 16538
rect 28626 16532 28632 16584
rect 28684 16581 28690 16584
rect 28828 16581 28856 16612
rect 28684 16575 28723 16581
rect 28711 16541 28723 16575
rect 28684 16535 28723 16541
rect 28813 16575 28871 16581
rect 28813 16541 28825 16575
rect 28859 16541 28871 16575
rect 28966 16572 28994 16612
rect 36740 16612 36820 16640
rect 31386 16572 31392 16584
rect 28966 16544 31392 16572
rect 28813 16535 28871 16541
rect 28684 16532 28690 16535
rect 31386 16532 31392 16544
rect 31444 16532 31450 16584
rect 31726 16544 35112 16572
rect 27982 16504 27988 16516
rect 26252 16476 27988 16504
rect 27982 16464 27988 16476
rect 28040 16464 28046 16516
rect 28442 16464 28448 16516
rect 28500 16464 28506 16516
rect 28537 16507 28595 16513
rect 28537 16473 28549 16507
rect 28583 16504 28595 16507
rect 30006 16504 30012 16516
rect 28583 16476 30012 16504
rect 28583 16473 28595 16476
rect 28537 16467 28595 16473
rect 30006 16464 30012 16476
rect 30064 16464 30070 16516
rect 31726 16504 31754 16544
rect 30116 16476 31754 16504
rect 20036 16408 21312 16436
rect 20036 16396 20042 16408
rect 22554 16396 22560 16448
rect 22612 16436 22618 16448
rect 23201 16439 23259 16445
rect 23201 16436 23213 16439
rect 22612 16408 23213 16436
rect 22612 16396 22618 16408
rect 23201 16405 23213 16408
rect 23247 16405 23259 16439
rect 23201 16399 23259 16405
rect 23382 16396 23388 16448
rect 23440 16436 23446 16448
rect 24486 16436 24492 16448
rect 23440 16408 24492 16436
rect 23440 16396 23446 16408
rect 24486 16396 24492 16408
rect 24544 16396 24550 16448
rect 27430 16396 27436 16448
rect 27488 16436 27494 16448
rect 30116 16436 30144 16476
rect 33594 16464 33600 16516
rect 33652 16504 33658 16516
rect 34054 16504 34060 16516
rect 33652 16476 34060 16504
rect 33652 16464 33658 16476
rect 34054 16464 34060 16476
rect 34112 16464 34118 16516
rect 27488 16408 30144 16436
rect 27488 16396 27494 16408
rect 30742 16396 30748 16448
rect 30800 16436 30806 16448
rect 31938 16436 31944 16448
rect 30800 16408 31944 16436
rect 30800 16396 30806 16408
rect 31938 16396 31944 16408
rect 31996 16436 32002 16448
rect 34974 16436 34980 16448
rect 31996 16408 34980 16436
rect 31996 16396 32002 16408
rect 34974 16396 34980 16408
rect 35032 16396 35038 16448
rect 35084 16436 35112 16544
rect 36354 16532 36360 16584
rect 36412 16572 36418 16584
rect 36630 16581 36636 16584
rect 36449 16575 36507 16581
rect 36449 16572 36461 16575
rect 36412 16544 36461 16572
rect 36412 16532 36418 16544
rect 36449 16541 36461 16544
rect 36495 16541 36507 16575
rect 36449 16535 36507 16541
rect 36597 16575 36636 16581
rect 36597 16541 36609 16575
rect 36597 16535 36636 16541
rect 36630 16532 36636 16535
rect 36688 16532 36694 16584
rect 36740 16581 36768 16612
rect 36814 16600 36820 16612
rect 36872 16600 36878 16652
rect 38470 16600 38476 16652
rect 38528 16600 38534 16652
rect 36725 16575 36783 16581
rect 36725 16541 36737 16575
rect 36771 16541 36783 16575
rect 36725 16535 36783 16541
rect 36955 16575 37013 16581
rect 36955 16541 36967 16575
rect 37001 16572 37013 16575
rect 37458 16572 37464 16584
rect 37001 16544 37464 16572
rect 37001 16541 37013 16544
rect 36955 16535 37013 16541
rect 37458 16532 37464 16544
rect 37516 16572 37522 16584
rect 38010 16572 38016 16584
rect 37516 16544 38016 16572
rect 37516 16532 37522 16544
rect 38010 16532 38016 16544
rect 38068 16532 38074 16584
rect 38381 16575 38439 16581
rect 38381 16541 38393 16575
rect 38427 16541 38439 16575
rect 38381 16535 38439 16541
rect 36817 16507 36875 16513
rect 36817 16473 36829 16507
rect 36863 16473 36875 16507
rect 38396 16504 38424 16535
rect 36817 16467 36875 16473
rect 37016 16476 38424 16504
rect 36832 16436 36860 16467
rect 37016 16448 37044 16476
rect 35084 16408 36860 16436
rect 36998 16396 37004 16448
rect 37056 16396 37062 16448
rect 38749 16439 38807 16445
rect 38749 16405 38761 16439
rect 38795 16436 38807 16439
rect 39482 16436 39488 16448
rect 38795 16408 39488 16436
rect 38795 16405 38807 16408
rect 38749 16399 38807 16405
rect 39482 16396 39488 16408
rect 39540 16396 39546 16448
rect 1104 16346 40572 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 40572 16346
rect 1104 16272 40572 16294
rect 4709 16235 4767 16241
rect 4709 16201 4721 16235
rect 4755 16232 4767 16235
rect 5261 16235 5319 16241
rect 5261 16232 5273 16235
rect 4755 16204 5273 16232
rect 4755 16201 4767 16204
rect 4709 16195 4767 16201
rect 5261 16201 5273 16204
rect 5307 16232 5319 16235
rect 7098 16232 7104 16244
rect 5307 16204 7104 16232
rect 5307 16201 5319 16204
rect 5261 16195 5319 16201
rect 7098 16192 7104 16204
rect 7156 16192 7162 16244
rect 7282 16192 7288 16244
rect 7340 16232 7346 16244
rect 7469 16235 7527 16241
rect 7469 16232 7481 16235
rect 7340 16204 7481 16232
rect 7340 16192 7346 16204
rect 7469 16201 7481 16204
rect 7515 16201 7527 16235
rect 7469 16195 7527 16201
rect 8202 16192 8208 16244
rect 8260 16232 8266 16244
rect 8297 16235 8355 16241
rect 8297 16232 8309 16235
rect 8260 16204 8309 16232
rect 8260 16192 8266 16204
rect 8297 16201 8309 16204
rect 8343 16201 8355 16235
rect 8297 16195 8355 16201
rect 9490 16192 9496 16244
rect 9548 16232 9554 16244
rect 10965 16235 11023 16241
rect 9548 16204 10824 16232
rect 9548 16192 9554 16204
rect 3234 16164 3240 16176
rect 2976 16136 3240 16164
rect 2976 16105 3004 16136
rect 3234 16124 3240 16136
rect 3292 16124 3298 16176
rect 3786 16124 3792 16176
rect 3844 16124 3850 16176
rect 10686 16164 10692 16176
rect 7484 16136 8432 16164
rect 2961 16099 3019 16105
rect 2961 16065 2973 16099
rect 3007 16065 3019 16099
rect 2961 16059 3019 16065
rect 5169 16099 5227 16105
rect 5169 16065 5181 16099
rect 5215 16096 5227 16099
rect 5442 16096 5448 16108
rect 5215 16068 5448 16096
rect 5215 16065 5227 16068
rect 5169 16059 5227 16065
rect 5442 16056 5448 16068
rect 5500 16056 5506 16108
rect 7484 16105 7512 16136
rect 7469 16099 7527 16105
rect 7469 16065 7481 16099
rect 7515 16065 7527 16099
rect 7469 16059 7527 16065
rect 7653 16099 7711 16105
rect 7653 16065 7665 16099
rect 7699 16065 7711 16099
rect 7653 16059 7711 16065
rect 3237 16031 3295 16037
rect 3237 15997 3249 16031
rect 3283 16028 3295 16031
rect 5353 16031 5411 16037
rect 3283 16000 4844 16028
rect 3283 15997 3295 16000
rect 3237 15991 3295 15997
rect 4816 15969 4844 16000
rect 5353 15997 5365 16031
rect 5399 16028 5411 16031
rect 5810 16028 5816 16040
rect 5399 16000 5816 16028
rect 5399 15997 5411 16000
rect 5353 15991 5411 15997
rect 5810 15988 5816 16000
rect 5868 15988 5874 16040
rect 4801 15963 4859 15969
rect 4801 15929 4813 15963
rect 4847 15929 4859 15963
rect 7668 15960 7696 16059
rect 8404 16028 8432 16136
rect 8496 16136 10692 16164
rect 8496 16105 8524 16136
rect 10686 16124 10692 16136
rect 10744 16124 10750 16176
rect 8481 16099 8539 16105
rect 8481 16065 8493 16099
rect 8527 16065 8539 16099
rect 8481 16059 8539 16065
rect 8665 16099 8723 16105
rect 8665 16065 8677 16099
rect 8711 16096 8723 16099
rect 9398 16096 9404 16108
rect 8711 16068 9404 16096
rect 8711 16065 8723 16068
rect 8665 16059 8723 16065
rect 8680 16028 8708 16059
rect 9398 16056 9404 16068
rect 9456 16056 9462 16108
rect 10796 16096 10824 16204
rect 10965 16201 10977 16235
rect 11011 16232 11023 16235
rect 11054 16232 11060 16244
rect 11011 16204 11060 16232
rect 11011 16201 11023 16204
rect 10965 16195 11023 16201
rect 11054 16192 11060 16204
rect 11112 16192 11118 16244
rect 11698 16192 11704 16244
rect 11756 16232 11762 16244
rect 11885 16235 11943 16241
rect 11885 16232 11897 16235
rect 11756 16204 11897 16232
rect 11756 16192 11762 16204
rect 11885 16201 11897 16204
rect 11931 16201 11943 16235
rect 11885 16195 11943 16201
rect 12250 16192 12256 16244
rect 12308 16232 12314 16244
rect 24762 16232 24768 16244
rect 12308 16204 24768 16232
rect 12308 16192 12314 16204
rect 24762 16192 24768 16204
rect 24820 16192 24826 16244
rect 25866 16192 25872 16244
rect 25924 16232 25930 16244
rect 26326 16232 26332 16244
rect 25924 16204 26332 16232
rect 25924 16192 25930 16204
rect 26326 16192 26332 16204
rect 26384 16192 26390 16244
rect 26418 16192 26424 16244
rect 26476 16232 26482 16244
rect 26973 16235 27031 16241
rect 26973 16232 26985 16235
rect 26476 16204 26985 16232
rect 26476 16192 26482 16204
rect 26973 16201 26985 16204
rect 27019 16201 27031 16235
rect 28074 16232 28080 16244
rect 26973 16195 27031 16201
rect 27080 16204 28080 16232
rect 10873 16167 10931 16173
rect 10873 16133 10885 16167
rect 10919 16164 10931 16167
rect 11238 16164 11244 16176
rect 10919 16136 11244 16164
rect 10919 16133 10931 16136
rect 10873 16127 10931 16133
rect 11238 16124 11244 16136
rect 11296 16124 11302 16176
rect 12529 16167 12587 16173
rect 12529 16133 12541 16167
rect 12575 16164 12587 16167
rect 12986 16164 12992 16176
rect 12575 16136 12992 16164
rect 12575 16133 12587 16136
rect 12529 16127 12587 16133
rect 12986 16124 12992 16136
rect 13044 16124 13050 16176
rect 13985 16167 14043 16173
rect 13985 16133 13997 16167
rect 14031 16164 14043 16167
rect 14090 16164 14096 16176
rect 14031 16136 14096 16164
rect 14031 16133 14043 16136
rect 13985 16127 14043 16133
rect 14090 16124 14096 16136
rect 14148 16124 14154 16176
rect 14185 16167 14243 16173
rect 14185 16133 14197 16167
rect 14231 16164 14243 16167
rect 14458 16164 14464 16176
rect 14231 16136 14464 16164
rect 14231 16133 14243 16136
rect 14185 16127 14243 16133
rect 10796 16068 11928 16096
rect 8404 16000 8708 16028
rect 11057 16031 11115 16037
rect 11057 15997 11069 16031
rect 11103 15997 11115 16031
rect 11900 16028 11928 16068
rect 11974 16056 11980 16108
rect 12032 16056 12038 16108
rect 12713 16099 12771 16105
rect 12713 16065 12725 16099
rect 12759 16096 12771 16099
rect 12802 16096 12808 16108
rect 12759 16068 12808 16096
rect 12759 16065 12771 16068
rect 12713 16059 12771 16065
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 13357 16099 13415 16105
rect 13357 16065 13369 16099
rect 13403 16065 13415 16099
rect 13357 16059 13415 16065
rect 12069 16031 12127 16037
rect 12069 16028 12081 16031
rect 11900 16000 12081 16028
rect 11057 15991 11115 15997
rect 12069 15997 12081 16000
rect 12115 16028 12127 16031
rect 13372 16028 13400 16059
rect 13630 16056 13636 16108
rect 13688 16056 13694 16108
rect 13814 16056 13820 16108
rect 13872 16096 13878 16108
rect 14200 16096 14228 16127
rect 14458 16124 14464 16136
rect 14516 16124 14522 16176
rect 14550 16124 14556 16176
rect 14608 16164 14614 16176
rect 14829 16167 14887 16173
rect 14829 16164 14841 16167
rect 14608 16136 14841 16164
rect 14608 16124 14614 16136
rect 14829 16133 14841 16136
rect 14875 16133 14887 16167
rect 16482 16164 16488 16176
rect 14829 16127 14887 16133
rect 16040 16136 16488 16164
rect 13872 16068 14228 16096
rect 15013 16099 15071 16105
rect 13872 16056 13878 16068
rect 15013 16065 15025 16099
rect 15059 16096 15071 16099
rect 15102 16096 15108 16108
rect 15059 16068 15108 16096
rect 15059 16065 15071 16068
rect 15013 16059 15071 16065
rect 15102 16056 15108 16068
rect 15160 16056 15166 16108
rect 16040 16105 16068 16136
rect 16482 16124 16488 16136
rect 16540 16124 16546 16176
rect 22278 16124 22284 16176
rect 22336 16164 22342 16176
rect 24121 16167 24179 16173
rect 24121 16164 24133 16167
rect 22336 16136 24133 16164
rect 22336 16124 22342 16136
rect 24121 16133 24133 16136
rect 24167 16133 24179 16167
rect 25682 16164 25688 16176
rect 24121 16127 24179 16133
rect 24320 16136 25688 16164
rect 15197 16099 15255 16105
rect 15197 16065 15209 16099
rect 15243 16096 15255 16099
rect 15841 16099 15899 16105
rect 15841 16096 15853 16099
rect 15243 16068 15853 16096
rect 15243 16065 15255 16068
rect 15197 16059 15255 16065
rect 15841 16065 15853 16068
rect 15887 16065 15899 16099
rect 15841 16059 15899 16065
rect 16025 16099 16083 16105
rect 16025 16065 16037 16099
rect 16071 16065 16083 16099
rect 16025 16059 16083 16065
rect 16114 16056 16120 16108
rect 16172 16056 16178 16108
rect 16301 16099 16359 16105
rect 16301 16065 16313 16099
rect 16347 16065 16359 16099
rect 16301 16059 16359 16065
rect 12115 16000 13400 16028
rect 13541 16031 13599 16037
rect 12115 15997 12127 16000
rect 12069 15991 12127 15997
rect 10505 15963 10563 15969
rect 10505 15960 10517 15963
rect 7668 15932 10517 15960
rect 4801 15923 4859 15929
rect 10505 15929 10517 15932
rect 10551 15929 10563 15963
rect 10505 15923 10563 15929
rect 10870 15920 10876 15972
rect 10928 15960 10934 15972
rect 11072 15960 11100 15991
rect 12176 15972 12204 16000
rect 13541 15997 13553 16031
rect 13587 16028 13599 16031
rect 14366 16028 14372 16040
rect 13587 16000 14372 16028
rect 13587 15997 13599 16000
rect 13541 15991 13599 15997
rect 14366 15988 14372 16000
rect 14424 15988 14430 16040
rect 16316 16028 16344 16059
rect 16390 16056 16396 16108
rect 16448 16056 16454 16108
rect 24320 16105 24348 16136
rect 25682 16124 25688 16136
rect 25740 16124 25746 16176
rect 24305 16099 24363 16105
rect 24305 16065 24317 16099
rect 24351 16065 24363 16099
rect 24305 16059 24363 16065
rect 24486 16056 24492 16108
rect 24544 16056 24550 16108
rect 24581 16099 24639 16105
rect 24581 16065 24593 16099
rect 24627 16096 24639 16099
rect 24670 16096 24676 16108
rect 24627 16068 24676 16096
rect 24627 16065 24639 16068
rect 24581 16059 24639 16065
rect 24670 16056 24676 16068
rect 24728 16096 24734 16108
rect 25222 16096 25228 16108
rect 24728 16068 25228 16096
rect 24728 16056 24734 16068
rect 25222 16056 25228 16068
rect 25280 16096 25286 16108
rect 27080 16096 27108 16204
rect 28074 16192 28080 16204
rect 28132 16232 28138 16244
rect 29546 16232 29552 16244
rect 28132 16204 29552 16232
rect 28132 16192 28138 16204
rect 29546 16192 29552 16204
rect 29604 16192 29610 16244
rect 30006 16192 30012 16244
rect 30064 16192 30070 16244
rect 30466 16232 30472 16244
rect 30208 16204 30472 16232
rect 27522 16164 27528 16176
rect 27172 16136 27528 16164
rect 27172 16105 27200 16136
rect 27522 16124 27528 16136
rect 27580 16124 27586 16176
rect 25280 16068 27108 16096
rect 27157 16099 27215 16105
rect 25280 16056 25286 16068
rect 27157 16065 27169 16099
rect 27203 16065 27215 16099
rect 27157 16059 27215 16065
rect 27430 16056 27436 16108
rect 27488 16056 27494 16108
rect 27617 16099 27675 16105
rect 27617 16065 27629 16099
rect 27663 16096 27675 16099
rect 27706 16096 27712 16108
rect 27663 16068 27712 16096
rect 27663 16065 27675 16068
rect 27617 16059 27675 16065
rect 27706 16056 27712 16068
rect 27764 16056 27770 16108
rect 27982 16056 27988 16108
rect 28040 16096 28046 16108
rect 28169 16099 28227 16105
rect 28169 16096 28181 16099
rect 28040 16068 28181 16096
rect 28040 16056 28046 16068
rect 28169 16065 28181 16068
rect 28215 16096 28227 16099
rect 28258 16096 28264 16108
rect 28215 16068 28264 16096
rect 28215 16065 28227 16068
rect 28169 16059 28227 16065
rect 28258 16056 28264 16068
rect 28316 16056 28322 16108
rect 28350 16056 28356 16108
rect 28408 16056 28414 16108
rect 30208 16105 30236 16204
rect 30466 16192 30472 16204
rect 30524 16192 30530 16244
rect 34808 16204 36952 16232
rect 30374 16124 30380 16176
rect 30432 16124 30438 16176
rect 31294 16124 31300 16176
rect 31352 16124 31358 16176
rect 33318 16124 33324 16176
rect 33376 16164 33382 16176
rect 34054 16164 34060 16176
rect 33376 16136 34060 16164
rect 33376 16124 33382 16136
rect 34054 16124 34060 16136
rect 34112 16164 34118 16176
rect 34238 16164 34244 16176
rect 34112 16136 34244 16164
rect 34112 16124 34118 16136
rect 34238 16124 34244 16136
rect 34296 16173 34302 16176
rect 34296 16167 34345 16173
rect 34296 16133 34299 16167
rect 34333 16133 34345 16167
rect 34296 16127 34345 16133
rect 34296 16124 34302 16127
rect 34422 16124 34428 16176
rect 34480 16124 34486 16176
rect 30193 16099 30251 16105
rect 30193 16065 30205 16099
rect 30239 16065 30251 16099
rect 30193 16059 30251 16065
rect 30285 16099 30343 16105
rect 30285 16065 30297 16099
rect 30331 16065 30343 16099
rect 30285 16059 30343 16065
rect 17402 16028 17408 16040
rect 16316 16000 17408 16028
rect 17402 15988 17408 16000
rect 17460 15988 17466 16040
rect 28077 16031 28135 16037
rect 28077 15997 28089 16031
rect 28123 16028 28135 16031
rect 29270 16028 29276 16040
rect 28123 16000 29276 16028
rect 28123 15997 28135 16000
rect 28077 15991 28135 15997
rect 29270 15988 29276 16000
rect 29328 15988 29334 16040
rect 10928 15932 11100 15960
rect 10928 15920 10934 15932
rect 12158 15920 12164 15972
rect 12216 15920 12222 15972
rect 13449 15963 13507 15969
rect 13449 15929 13461 15963
rect 13495 15929 13507 15963
rect 13449 15923 13507 15929
rect 11422 15852 11428 15904
rect 11480 15892 11486 15904
rect 11517 15895 11575 15901
rect 11517 15892 11529 15895
rect 11480 15864 11529 15892
rect 11480 15852 11486 15864
rect 11517 15861 11529 15864
rect 11563 15861 11575 15895
rect 11517 15855 11575 15861
rect 11790 15852 11796 15904
rect 11848 15892 11854 15904
rect 12345 15895 12403 15901
rect 12345 15892 12357 15895
rect 11848 15864 12357 15892
rect 11848 15852 11854 15864
rect 12345 15861 12357 15864
rect 12391 15861 12403 15895
rect 12345 15855 12403 15861
rect 13173 15895 13231 15901
rect 13173 15861 13185 15895
rect 13219 15892 13231 15895
rect 13262 15892 13268 15904
rect 13219 15864 13268 15892
rect 13219 15861 13231 15864
rect 13173 15855 13231 15861
rect 13262 15852 13268 15864
rect 13320 15852 13326 15904
rect 13464 15892 13492 15923
rect 15838 15920 15844 15972
rect 15896 15960 15902 15972
rect 16114 15960 16120 15972
rect 15896 15932 16120 15960
rect 15896 15920 15902 15932
rect 16114 15920 16120 15932
rect 16172 15920 16178 15972
rect 20714 15920 20720 15972
rect 20772 15960 20778 15972
rect 27246 15960 27252 15972
rect 20772 15932 27252 15960
rect 20772 15920 20778 15932
rect 27246 15920 27252 15932
rect 27304 15920 27310 15972
rect 27341 15963 27399 15969
rect 27341 15929 27353 15963
rect 27387 15960 27399 15963
rect 28442 15960 28448 15972
rect 27387 15932 28448 15960
rect 27387 15929 27399 15932
rect 27341 15923 27399 15929
rect 28442 15920 28448 15932
rect 28500 15920 28506 15972
rect 30300 15960 30328 16059
rect 30558 16056 30564 16108
rect 30616 16056 30622 16108
rect 30742 16056 30748 16108
rect 30800 16096 30806 16108
rect 31159 16099 31217 16105
rect 31159 16096 31171 16099
rect 30800 16068 31171 16096
rect 30800 16056 30806 16068
rect 31159 16065 31171 16068
rect 31205 16065 31217 16099
rect 31159 16059 31217 16065
rect 31386 16056 31392 16108
rect 31444 16056 31450 16108
rect 31478 16056 31484 16108
rect 31536 16056 31542 16108
rect 33226 16056 33232 16108
rect 33284 16096 33290 16108
rect 33870 16096 33876 16108
rect 33284 16068 33876 16096
rect 33284 16056 33290 16068
rect 33870 16056 33876 16068
rect 33928 16096 33934 16108
rect 34149 16099 34207 16105
rect 34149 16096 34161 16099
rect 33928 16068 34161 16096
rect 33928 16056 33934 16068
rect 34149 16065 34161 16068
rect 34195 16065 34207 16099
rect 34149 16059 34207 16065
rect 34514 16056 34520 16108
rect 34572 16056 34578 16108
rect 34609 16099 34667 16105
rect 34609 16065 34621 16099
rect 34655 16096 34667 16099
rect 34808 16096 34836 16204
rect 35158 16124 35164 16176
rect 35216 16124 35222 16176
rect 36814 16124 36820 16176
rect 36872 16124 36878 16176
rect 34655 16068 34836 16096
rect 34655 16065 34667 16068
rect 34609 16059 34667 16065
rect 34882 16056 34888 16108
rect 34940 16056 34946 16108
rect 36538 16056 36544 16108
rect 36596 16056 36602 16108
rect 36924 16105 36952 16204
rect 36725 16099 36783 16105
rect 36725 16065 36737 16099
rect 36771 16065 36783 16099
rect 36725 16059 36783 16065
rect 36909 16099 36967 16105
rect 36909 16065 36921 16099
rect 36955 16096 36967 16099
rect 37458 16096 37464 16108
rect 36955 16068 37464 16096
rect 36955 16065 36967 16068
rect 36909 16059 36967 16065
rect 31018 15988 31024 16040
rect 31076 16028 31082 16040
rect 31570 16028 31576 16040
rect 31076 16000 31576 16028
rect 31076 15988 31082 16000
rect 31570 15988 31576 16000
rect 31628 15988 31634 16040
rect 34238 15988 34244 16040
rect 34296 16028 34302 16040
rect 34532 16028 34560 16056
rect 34296 16000 34560 16028
rect 34296 15988 34302 16000
rect 34790 15988 34796 16040
rect 34848 15988 34854 16040
rect 34974 15988 34980 16040
rect 35032 16028 35038 16040
rect 36740 16028 36768 16059
rect 37458 16056 37464 16068
rect 37516 16056 37522 16108
rect 35032 16000 36768 16028
rect 35032 15988 35038 16000
rect 31294 15960 31300 15972
rect 30300 15932 31300 15960
rect 31294 15920 31300 15932
rect 31352 15920 31358 15972
rect 31665 15963 31723 15969
rect 31665 15929 31677 15963
rect 31711 15960 31723 15963
rect 38286 15960 38292 15972
rect 31711 15932 38292 15960
rect 31711 15929 31723 15932
rect 31665 15923 31723 15929
rect 38286 15920 38292 15932
rect 38344 15920 38350 15972
rect 13817 15895 13875 15901
rect 13817 15892 13829 15895
rect 13464 15864 13829 15892
rect 13817 15861 13829 15864
rect 13863 15861 13875 15895
rect 13817 15855 13875 15861
rect 14001 15895 14059 15901
rect 14001 15861 14013 15895
rect 14047 15892 14059 15895
rect 14182 15892 14188 15904
rect 14047 15864 14188 15892
rect 14047 15861 14059 15864
rect 14001 15855 14059 15861
rect 14182 15852 14188 15864
rect 14240 15852 14246 15904
rect 18414 15852 18420 15904
rect 18472 15892 18478 15904
rect 27522 15892 27528 15904
rect 18472 15864 27528 15892
rect 18472 15852 18478 15864
rect 27522 15852 27528 15864
rect 27580 15852 27586 15904
rect 27890 15852 27896 15904
rect 27948 15852 27954 15904
rect 27982 15852 27988 15904
rect 28040 15852 28046 15904
rect 28074 15852 28080 15904
rect 28132 15892 28138 15904
rect 28350 15892 28356 15904
rect 28132 15864 28356 15892
rect 28132 15852 28138 15864
rect 28350 15852 28356 15864
rect 28408 15852 28414 15904
rect 28902 15852 28908 15904
rect 28960 15892 28966 15904
rect 30282 15892 30288 15904
rect 28960 15864 30288 15892
rect 28960 15852 28966 15864
rect 30282 15852 30288 15864
rect 30340 15852 30346 15904
rect 30834 15852 30840 15904
rect 30892 15892 30898 15904
rect 32766 15892 32772 15904
rect 30892 15864 32772 15892
rect 30892 15852 30898 15864
rect 32766 15852 32772 15864
rect 32824 15852 32830 15904
rect 33778 15852 33784 15904
rect 33836 15892 33842 15904
rect 34882 15892 34888 15904
rect 33836 15864 34888 15892
rect 33836 15852 33842 15864
rect 34882 15852 34888 15864
rect 34940 15852 34946 15904
rect 37090 15852 37096 15904
rect 37148 15852 37154 15904
rect 1104 15802 40572 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 40572 15802
rect 1104 15728 40572 15750
rect 5442 15648 5448 15700
rect 5500 15648 5506 15700
rect 6086 15648 6092 15700
rect 6144 15688 6150 15700
rect 6181 15691 6239 15697
rect 6181 15688 6193 15691
rect 6144 15660 6193 15688
rect 6144 15648 6150 15660
rect 6181 15657 6193 15660
rect 6227 15657 6239 15691
rect 6181 15651 6239 15657
rect 9858 15648 9864 15700
rect 9916 15688 9922 15700
rect 10229 15691 10287 15697
rect 10229 15688 10241 15691
rect 9916 15660 10241 15688
rect 9916 15648 9922 15660
rect 10229 15657 10241 15660
rect 10275 15657 10287 15691
rect 10229 15651 10287 15657
rect 5994 15580 6000 15632
rect 6052 15620 6058 15632
rect 7009 15623 7067 15629
rect 7009 15620 7021 15623
rect 6052 15592 7021 15620
rect 6052 15580 6058 15592
rect 4893 15555 4951 15561
rect 4893 15521 4905 15555
rect 4939 15552 4951 15555
rect 5258 15552 5264 15564
rect 4939 15524 5264 15552
rect 4939 15521 4951 15524
rect 4893 15515 4951 15521
rect 5258 15512 5264 15524
rect 5316 15552 5322 15564
rect 5316 15524 5672 15552
rect 5316 15512 5322 15524
rect 5534 15444 5540 15496
rect 5592 15444 5598 15496
rect 5644 15493 5672 15524
rect 5810 15512 5816 15564
rect 5868 15512 5874 15564
rect 5902 15512 5908 15564
rect 5960 15552 5966 15564
rect 5960 15524 6316 15552
rect 5960 15512 5966 15524
rect 5630 15487 5688 15493
rect 5630 15453 5642 15487
rect 5676 15453 5688 15487
rect 5828 15484 5856 15512
rect 6043 15487 6101 15493
rect 6043 15484 6055 15487
rect 5828 15456 6055 15484
rect 5630 15447 5688 15453
rect 6043 15453 6055 15456
rect 6089 15484 6101 15487
rect 6178 15484 6184 15496
rect 6089 15456 6184 15484
rect 6089 15453 6101 15456
rect 6043 15447 6101 15453
rect 6178 15444 6184 15456
rect 6236 15444 6242 15496
rect 6288 15493 6316 15524
rect 6472 15493 6500 15592
rect 7009 15589 7021 15592
rect 7055 15589 7067 15623
rect 7009 15583 7067 15589
rect 6273 15487 6331 15493
rect 6273 15453 6285 15487
rect 6319 15453 6331 15487
rect 6273 15447 6331 15453
rect 6457 15487 6515 15493
rect 6457 15453 6469 15487
rect 6503 15453 6515 15487
rect 6457 15447 6515 15453
rect 6546 15444 6552 15496
rect 6604 15444 6610 15496
rect 6822 15444 6828 15496
rect 6880 15444 6886 15496
rect 7006 15444 7012 15496
rect 7064 15444 7070 15496
rect 8018 15444 8024 15496
rect 8076 15444 8082 15496
rect 10042 15444 10048 15496
rect 10100 15444 10106 15496
rect 10244 15484 10272 15651
rect 16390 15648 16396 15700
rect 16448 15648 16454 15700
rect 16758 15648 16764 15700
rect 16816 15688 16822 15700
rect 16853 15691 16911 15697
rect 16853 15688 16865 15691
rect 16816 15660 16865 15688
rect 16816 15648 16822 15660
rect 16853 15657 16865 15660
rect 16899 15657 16911 15691
rect 16853 15651 16911 15657
rect 16868 15620 16896 15651
rect 17034 15648 17040 15700
rect 17092 15648 17098 15700
rect 17402 15648 17408 15700
rect 17460 15648 17466 15700
rect 19426 15648 19432 15700
rect 19484 15688 19490 15700
rect 21542 15688 21548 15700
rect 19484 15660 21548 15688
rect 19484 15648 19490 15660
rect 21542 15648 21548 15660
rect 21600 15648 21606 15700
rect 22002 15648 22008 15700
rect 22060 15648 22066 15700
rect 22186 15648 22192 15700
rect 22244 15688 22250 15700
rect 24670 15688 24676 15700
rect 22244 15660 24676 15688
rect 22244 15648 22250 15660
rect 24670 15648 24676 15660
rect 24728 15648 24734 15700
rect 27246 15648 27252 15700
rect 27304 15688 27310 15700
rect 28718 15688 28724 15700
rect 27304 15660 28724 15688
rect 27304 15648 27310 15660
rect 28718 15648 28724 15660
rect 28776 15688 28782 15700
rect 31846 15688 31852 15700
rect 28776 15660 31852 15688
rect 28776 15648 28782 15660
rect 31846 15648 31852 15660
rect 31904 15648 31910 15700
rect 33042 15648 33048 15700
rect 33100 15648 33106 15700
rect 34330 15648 34336 15700
rect 34388 15688 34394 15700
rect 34698 15688 34704 15700
rect 34388 15660 34704 15688
rect 34388 15648 34394 15660
rect 34698 15648 34704 15660
rect 34756 15648 34762 15700
rect 34974 15648 34980 15700
rect 35032 15648 35038 15700
rect 35345 15691 35403 15697
rect 35345 15657 35357 15691
rect 35391 15688 35403 15691
rect 37918 15688 37924 15700
rect 35391 15660 37924 15688
rect 35391 15657 35403 15660
rect 35345 15651 35403 15657
rect 37918 15648 37924 15660
rect 37976 15648 37982 15700
rect 38286 15648 38292 15700
rect 38344 15648 38350 15700
rect 16868 15592 18644 15620
rect 10321 15555 10379 15561
rect 10321 15521 10333 15555
rect 10367 15552 10379 15555
rect 10505 15555 10563 15561
rect 10505 15552 10517 15555
rect 10367 15524 10517 15552
rect 10367 15521 10379 15524
rect 10321 15515 10379 15521
rect 10505 15521 10517 15524
rect 10551 15552 10563 15555
rect 11333 15555 11391 15561
rect 11333 15552 11345 15555
rect 10551 15524 11345 15552
rect 10551 15521 10563 15524
rect 10505 15515 10563 15521
rect 11333 15521 11345 15524
rect 11379 15521 11391 15555
rect 11333 15515 11391 15521
rect 17129 15555 17187 15561
rect 17129 15521 17141 15555
rect 17175 15552 17187 15555
rect 17586 15552 17592 15564
rect 17175 15524 17592 15552
rect 17175 15521 17187 15524
rect 17129 15515 17187 15521
rect 17586 15512 17592 15524
rect 17644 15512 17650 15564
rect 18506 15552 18512 15564
rect 17972 15524 18512 15552
rect 17972 15496 18000 15524
rect 18506 15512 18512 15524
rect 18564 15512 18570 15564
rect 18616 15552 18644 15592
rect 19334 15580 19340 15632
rect 19392 15620 19398 15632
rect 19392 15592 25176 15620
rect 19392 15580 19398 15592
rect 22002 15552 22008 15564
rect 18616 15524 22008 15552
rect 22002 15512 22008 15524
rect 22060 15512 22066 15564
rect 22094 15512 22100 15564
rect 22152 15552 22158 15564
rect 22281 15555 22339 15561
rect 22281 15552 22293 15555
rect 22152 15524 22293 15552
rect 22152 15512 22158 15524
rect 22281 15521 22293 15524
rect 22327 15521 22339 15555
rect 22281 15515 22339 15521
rect 22373 15555 22431 15561
rect 22373 15521 22385 15555
rect 22419 15552 22431 15555
rect 22830 15552 22836 15564
rect 22419 15524 22836 15552
rect 22419 15521 22431 15524
rect 22373 15515 22431 15521
rect 22830 15512 22836 15524
rect 22888 15512 22894 15564
rect 25148 15561 25176 15592
rect 30006 15580 30012 15632
rect 30064 15580 30070 15632
rect 31389 15623 31447 15629
rect 31389 15589 31401 15623
rect 31435 15589 31447 15623
rect 31389 15583 31447 15589
rect 31680 15592 32444 15620
rect 25133 15555 25191 15561
rect 25133 15521 25145 15555
rect 25179 15521 25191 15555
rect 29641 15555 29699 15561
rect 29641 15552 29653 15555
rect 25133 15515 25191 15521
rect 25516 15524 29653 15552
rect 10413 15487 10471 15493
rect 10413 15484 10425 15487
rect 10244 15456 10425 15484
rect 10413 15453 10425 15456
rect 10459 15453 10471 15487
rect 10413 15447 10471 15453
rect 11054 15444 11060 15496
rect 11112 15484 11118 15496
rect 11609 15487 11667 15493
rect 11609 15484 11621 15487
rect 11112 15456 11621 15484
rect 11112 15444 11118 15456
rect 11609 15453 11621 15456
rect 11655 15453 11667 15487
rect 11609 15447 11667 15453
rect 11701 15487 11759 15493
rect 11701 15453 11713 15487
rect 11747 15453 11759 15487
rect 11701 15447 11759 15453
rect 5810 15376 5816 15428
rect 5868 15376 5874 15428
rect 5905 15419 5963 15425
rect 5905 15385 5917 15419
rect 5951 15416 5963 15419
rect 6564 15416 6592 15444
rect 5951 15388 6592 15416
rect 10060 15416 10088 15444
rect 10502 15416 10508 15428
rect 10060 15388 10508 15416
rect 5951 15385 5963 15388
rect 5905 15379 5963 15385
rect 10502 15376 10508 15388
rect 10560 15416 10566 15428
rect 10689 15419 10747 15425
rect 10689 15416 10701 15419
rect 10560 15388 10701 15416
rect 10560 15376 10566 15388
rect 10689 15385 10701 15388
rect 10735 15385 10747 15419
rect 11716 15416 11744 15447
rect 11790 15444 11796 15496
rect 11848 15444 11854 15496
rect 11882 15444 11888 15496
rect 11940 15484 11946 15496
rect 11977 15487 12035 15493
rect 11977 15484 11989 15487
rect 11940 15456 11989 15484
rect 11940 15444 11946 15456
rect 11977 15453 11989 15456
rect 12023 15453 12035 15487
rect 11977 15447 12035 15453
rect 12526 15444 12532 15496
rect 12584 15484 12590 15496
rect 13170 15484 13176 15496
rect 12584 15456 13176 15484
rect 12584 15444 12590 15456
rect 13170 15444 13176 15456
rect 13228 15444 13234 15496
rect 16577 15487 16635 15493
rect 16577 15453 16589 15487
rect 16623 15453 16635 15487
rect 16577 15447 16635 15453
rect 12158 15416 12164 15428
rect 11716 15388 12164 15416
rect 10689 15379 10747 15385
rect 12158 15376 12164 15388
rect 12216 15376 12222 15428
rect 16592 15416 16620 15447
rect 16666 15444 16672 15496
rect 16724 15444 16730 15496
rect 16758 15444 16764 15496
rect 16816 15484 16822 15496
rect 16853 15487 16911 15493
rect 16853 15484 16865 15487
rect 16816 15456 16865 15484
rect 16816 15444 16822 15456
rect 16853 15453 16865 15456
rect 16899 15453 16911 15487
rect 16853 15447 16911 15453
rect 16942 15444 16948 15496
rect 17000 15444 17006 15496
rect 17221 15487 17279 15493
rect 17221 15453 17233 15487
rect 17267 15484 17279 15487
rect 17954 15484 17960 15496
rect 17267 15456 17960 15484
rect 17267 15453 17279 15456
rect 17221 15447 17279 15453
rect 17954 15444 17960 15456
rect 18012 15444 18018 15496
rect 18046 15444 18052 15496
rect 18104 15484 18110 15496
rect 18141 15487 18199 15493
rect 18141 15484 18153 15487
rect 18104 15456 18153 15484
rect 18104 15444 18110 15456
rect 18141 15453 18153 15456
rect 18187 15453 18199 15487
rect 18141 15447 18199 15453
rect 18230 15444 18236 15496
rect 18288 15484 18294 15496
rect 18325 15487 18383 15493
rect 18325 15484 18337 15487
rect 18288 15456 18337 15484
rect 18288 15444 18294 15456
rect 18325 15453 18337 15456
rect 18371 15453 18383 15487
rect 18325 15447 18383 15453
rect 18414 15444 18420 15496
rect 18472 15444 18478 15496
rect 20349 15487 20407 15493
rect 20349 15453 20361 15487
rect 20395 15484 20407 15487
rect 20530 15484 20536 15496
rect 20395 15456 20536 15484
rect 20395 15453 20407 15456
rect 20349 15447 20407 15453
rect 20530 15444 20536 15456
rect 20588 15444 20594 15496
rect 20625 15487 20683 15493
rect 20625 15453 20637 15487
rect 20671 15453 20683 15487
rect 20625 15447 20683 15453
rect 17770 15416 17776 15428
rect 16592 15388 17776 15416
rect 17770 15376 17776 15388
rect 17828 15416 17834 15428
rect 20165 15419 20223 15425
rect 20165 15416 20177 15419
rect 17828 15388 20177 15416
rect 17828 15376 17834 15388
rect 20165 15385 20177 15388
rect 20211 15385 20223 15419
rect 20640 15416 20668 15447
rect 22186 15444 22192 15496
rect 22244 15444 22250 15496
rect 22462 15444 22468 15496
rect 22520 15444 22526 15496
rect 23658 15444 23664 15496
rect 23716 15484 23722 15496
rect 24213 15487 24271 15493
rect 24213 15484 24225 15487
rect 23716 15456 24225 15484
rect 23716 15444 23722 15456
rect 24213 15453 24225 15456
rect 24259 15453 24271 15487
rect 24213 15447 24271 15453
rect 24394 15444 24400 15496
rect 24452 15444 24458 15496
rect 24670 15444 24676 15496
rect 24728 15484 24734 15496
rect 25516 15493 25544 15524
rect 29641 15521 29653 15524
rect 29687 15521 29699 15555
rect 29914 15552 29920 15564
rect 29641 15515 29699 15521
rect 29748 15524 29920 15552
rect 24765 15487 24823 15493
rect 24765 15484 24777 15487
rect 24728 15456 24777 15484
rect 24728 15444 24734 15456
rect 24765 15453 24777 15456
rect 24811 15453 24823 15487
rect 24765 15447 24823 15453
rect 25501 15487 25559 15493
rect 25501 15453 25513 15487
rect 25547 15453 25559 15487
rect 25501 15447 25559 15453
rect 25590 15444 25596 15496
rect 25648 15484 25654 15496
rect 25685 15487 25743 15493
rect 25685 15484 25697 15487
rect 25648 15456 25697 15484
rect 25648 15444 25654 15456
rect 25685 15453 25697 15456
rect 25731 15453 25743 15487
rect 25685 15447 25743 15453
rect 26234 15444 26240 15496
rect 26292 15484 26298 15496
rect 28902 15484 28908 15496
rect 26292 15456 28908 15484
rect 26292 15444 26298 15456
rect 28902 15444 28908 15456
rect 28960 15444 28966 15496
rect 28997 15487 29055 15493
rect 28997 15453 29009 15487
rect 29043 15484 29055 15487
rect 29086 15484 29092 15496
rect 29043 15456 29092 15484
rect 29043 15453 29055 15456
rect 28997 15447 29055 15453
rect 29086 15444 29092 15456
rect 29144 15444 29150 15496
rect 29181 15487 29239 15493
rect 29181 15453 29193 15487
rect 29227 15453 29239 15487
rect 29181 15447 29239 15453
rect 29273 15487 29331 15493
rect 29273 15453 29285 15487
rect 29319 15484 29331 15487
rect 29748 15484 29776 15524
rect 29914 15512 29920 15524
rect 29972 15512 29978 15564
rect 30024 15552 30052 15580
rect 30024 15524 30512 15552
rect 29319 15456 29776 15484
rect 29319 15453 29331 15456
rect 29273 15447 29331 15453
rect 23845 15419 23903 15425
rect 23845 15416 23857 15419
rect 20640 15388 23857 15416
rect 20165 15379 20223 15385
rect 23845 15385 23857 15388
rect 23891 15385 23903 15419
rect 23845 15379 23903 15385
rect 24026 15376 24032 15428
rect 24084 15376 24090 15428
rect 24118 15376 24124 15428
rect 24176 15416 24182 15428
rect 26418 15416 26424 15428
rect 24176 15388 26424 15416
rect 24176 15376 24182 15388
rect 26418 15376 26424 15388
rect 26476 15416 26482 15428
rect 29196 15416 29224 15447
rect 29822 15444 29828 15496
rect 29880 15444 29886 15496
rect 30009 15487 30067 15493
rect 30009 15453 30021 15487
rect 30055 15453 30067 15487
rect 30009 15447 30067 15453
rect 30101 15487 30159 15493
rect 30101 15453 30113 15487
rect 30147 15484 30159 15487
rect 30190 15484 30196 15496
rect 30147 15456 30196 15484
rect 30147 15453 30159 15456
rect 30101 15447 30159 15453
rect 29638 15416 29644 15428
rect 26476 15388 29644 15416
rect 26476 15376 26482 15388
rect 29638 15376 29644 15388
rect 29696 15376 29702 15428
rect 30024 15416 30052 15447
rect 30190 15444 30196 15456
rect 30248 15444 30254 15496
rect 30484 15493 30512 15524
rect 30469 15487 30527 15493
rect 30469 15453 30481 15487
rect 30515 15453 30527 15487
rect 30469 15447 30527 15453
rect 30834 15444 30840 15496
rect 30892 15444 30898 15496
rect 31018 15444 31024 15496
rect 31076 15444 31082 15496
rect 31202 15444 31208 15496
rect 31260 15444 31266 15496
rect 31404 15484 31432 15583
rect 31481 15487 31539 15493
rect 31481 15484 31493 15487
rect 31404 15456 31493 15484
rect 31481 15453 31493 15456
rect 31527 15453 31539 15487
rect 31481 15447 31539 15453
rect 30653 15419 30711 15425
rect 30653 15416 30665 15419
rect 30024 15388 30665 15416
rect 30653 15385 30665 15388
rect 30699 15416 30711 15419
rect 30742 15416 30748 15428
rect 30699 15388 30748 15416
rect 30699 15385 30711 15388
rect 30653 15379 30711 15385
rect 30742 15376 30748 15388
rect 30800 15376 30806 15428
rect 31113 15419 31171 15425
rect 31113 15385 31125 15419
rect 31159 15385 31171 15419
rect 31496 15416 31524 15447
rect 31570 15444 31576 15496
rect 31628 15444 31634 15496
rect 31680 15416 31708 15592
rect 32416 15493 32444 15592
rect 32490 15580 32496 15632
rect 32548 15580 32554 15632
rect 36538 15620 36544 15632
rect 34072 15592 36544 15620
rect 32508 15493 32536 15580
rect 32766 15512 32772 15564
rect 32824 15552 32830 15564
rect 34072 15552 34100 15592
rect 36538 15580 36544 15592
rect 36596 15580 36602 15632
rect 36630 15580 36636 15632
rect 36688 15620 36694 15632
rect 39206 15620 39212 15632
rect 36688 15592 39212 15620
rect 36688 15580 36694 15592
rect 39206 15580 39212 15592
rect 39264 15580 39270 15632
rect 32824 15524 34100 15552
rect 32824 15512 32830 15524
rect 34514 15512 34520 15564
rect 34572 15552 34578 15564
rect 35069 15555 35127 15561
rect 35069 15552 35081 15555
rect 34572 15524 35081 15552
rect 34572 15512 34578 15524
rect 35069 15521 35081 15524
rect 35115 15521 35127 15555
rect 35069 15515 35127 15521
rect 38473 15555 38531 15561
rect 38473 15521 38485 15555
rect 38519 15552 38531 15555
rect 38841 15555 38899 15561
rect 38841 15552 38853 15555
rect 38519 15524 38853 15552
rect 38519 15521 38531 15524
rect 38473 15515 38531 15521
rect 38841 15521 38853 15524
rect 38887 15521 38899 15555
rect 39301 15555 39359 15561
rect 39301 15552 39313 15555
rect 38841 15515 38899 15521
rect 38948 15524 39313 15552
rect 31946 15487 32004 15493
rect 31946 15453 31958 15487
rect 31992 15453 32004 15487
rect 31946 15447 32004 15453
rect 32401 15487 32459 15493
rect 32401 15453 32413 15487
rect 32447 15453 32459 15487
rect 32401 15447 32459 15453
rect 32494 15487 32552 15493
rect 32494 15453 32506 15487
rect 32540 15453 32552 15487
rect 32866 15487 32924 15493
rect 32866 15484 32878 15487
rect 32494 15447 32552 15453
rect 32600 15456 32878 15484
rect 31496 15388 31708 15416
rect 31113 15379 31171 15385
rect 4614 15308 4620 15360
rect 4672 15348 4678 15360
rect 4985 15351 5043 15357
rect 4985 15348 4997 15351
rect 4672 15320 4997 15348
rect 4672 15308 4678 15320
rect 4985 15317 4997 15320
rect 5031 15317 5043 15351
rect 4985 15311 5043 15317
rect 5077 15351 5135 15357
rect 5077 15317 5089 15351
rect 5123 15348 5135 15351
rect 6270 15348 6276 15360
rect 5123 15320 6276 15348
rect 5123 15317 5135 15320
rect 5077 15311 5135 15317
rect 6270 15308 6276 15320
rect 6328 15308 6334 15360
rect 6457 15351 6515 15357
rect 6457 15317 6469 15351
rect 6503 15348 6515 15351
rect 6546 15348 6552 15360
rect 6503 15320 6552 15348
rect 6503 15317 6515 15320
rect 6457 15311 6515 15317
rect 6546 15308 6552 15320
rect 6604 15308 6610 15360
rect 7926 15308 7932 15360
rect 7984 15308 7990 15360
rect 9861 15351 9919 15357
rect 9861 15317 9873 15351
rect 9907 15348 9919 15351
rect 10042 15348 10048 15360
rect 9907 15320 10048 15348
rect 9907 15317 9919 15320
rect 9861 15311 9919 15317
rect 10042 15308 10048 15320
rect 10100 15308 10106 15360
rect 10410 15308 10416 15360
rect 10468 15308 10474 15360
rect 13354 15308 13360 15360
rect 13412 15308 13418 15360
rect 17954 15308 17960 15360
rect 18012 15308 18018 15360
rect 20530 15308 20536 15360
rect 20588 15348 20594 15360
rect 21726 15348 21732 15360
rect 20588 15320 21732 15348
rect 20588 15308 20594 15320
rect 21726 15308 21732 15320
rect 21784 15348 21790 15360
rect 22646 15348 22652 15360
rect 21784 15320 22652 15348
rect 21784 15308 21790 15320
rect 22646 15308 22652 15320
rect 22704 15308 22710 15360
rect 28721 15351 28779 15357
rect 28721 15317 28733 15351
rect 28767 15348 28779 15351
rect 28902 15348 28908 15360
rect 28767 15320 28908 15348
rect 28767 15317 28779 15320
rect 28721 15311 28779 15317
rect 28902 15308 28908 15320
rect 28960 15308 28966 15360
rect 29270 15308 29276 15360
rect 29328 15348 29334 15360
rect 30190 15348 30196 15360
rect 29328 15320 30196 15348
rect 29328 15308 29334 15320
rect 30190 15308 30196 15320
rect 30248 15308 30254 15360
rect 30282 15308 30288 15360
rect 30340 15308 30346 15360
rect 30374 15308 30380 15360
rect 30432 15348 30438 15360
rect 31128 15348 31156 15379
rect 31754 15376 31760 15428
rect 31812 15376 31818 15428
rect 31846 15376 31852 15428
rect 31904 15376 31910 15428
rect 31961 15416 31989 15447
rect 32600 15416 32628 15456
rect 32866 15453 32878 15456
rect 32912 15453 32924 15487
rect 32866 15447 32924 15453
rect 34790 15444 34796 15496
rect 34848 15484 34854 15496
rect 34977 15487 35035 15493
rect 34977 15484 34989 15487
rect 34848 15456 34989 15484
rect 34848 15444 34854 15456
rect 34977 15453 34989 15456
rect 35023 15453 35035 15487
rect 34977 15447 35035 15453
rect 36906 15444 36912 15496
rect 36964 15484 36970 15496
rect 38562 15484 38568 15496
rect 36964 15456 38568 15484
rect 36964 15444 36970 15456
rect 38562 15444 38568 15456
rect 38620 15444 38626 15496
rect 38948 15484 38976 15524
rect 39301 15521 39313 15524
rect 39347 15521 39359 15555
rect 39301 15515 39359 15521
rect 38672 15456 38976 15484
rect 39025 15487 39083 15493
rect 31961 15388 32628 15416
rect 32677 15419 32735 15425
rect 30432 15320 31156 15348
rect 30432 15308 30438 15320
rect 31478 15308 31484 15360
rect 31536 15348 31542 15360
rect 31961 15348 31989 15388
rect 32677 15385 32689 15419
rect 32723 15385 32735 15419
rect 32677 15379 32735 15385
rect 32769 15419 32827 15425
rect 32769 15385 32781 15419
rect 32815 15416 32827 15419
rect 33226 15416 33232 15428
rect 32815 15388 33232 15416
rect 32815 15385 32827 15388
rect 32769 15379 32827 15385
rect 31536 15320 31989 15348
rect 31536 15308 31542 15320
rect 32122 15308 32128 15360
rect 32180 15308 32186 15360
rect 32692 15348 32720 15379
rect 33226 15376 33232 15388
rect 33284 15376 33290 15428
rect 37458 15376 37464 15428
rect 37516 15416 37522 15428
rect 38289 15419 38347 15425
rect 38289 15416 38301 15419
rect 37516 15388 38301 15416
rect 37516 15376 37522 15388
rect 38289 15385 38301 15388
rect 38335 15385 38347 15419
rect 38672 15416 38700 15456
rect 39025 15453 39037 15487
rect 39071 15484 39083 15487
rect 39114 15484 39120 15496
rect 39071 15456 39120 15484
rect 39071 15453 39083 15456
rect 39025 15447 39083 15453
rect 39114 15444 39120 15456
rect 39172 15484 39178 15496
rect 39390 15484 39396 15496
rect 39172 15456 39396 15484
rect 39172 15444 39178 15456
rect 39390 15444 39396 15456
rect 39448 15444 39454 15496
rect 38289 15379 38347 15385
rect 38580 15388 38700 15416
rect 33042 15348 33048 15360
rect 32692 15320 33048 15348
rect 33042 15308 33048 15320
rect 33100 15308 33106 15360
rect 33870 15308 33876 15360
rect 33928 15348 33934 15360
rect 36078 15348 36084 15360
rect 33928 15320 36084 15348
rect 33928 15308 33934 15320
rect 36078 15308 36084 15320
rect 36136 15348 36142 15360
rect 38580 15348 38608 15388
rect 36136 15320 38608 15348
rect 36136 15308 36142 15320
rect 38654 15308 38660 15360
rect 38712 15348 38718 15360
rect 38749 15351 38807 15357
rect 38749 15348 38761 15351
rect 38712 15320 38761 15348
rect 38712 15308 38718 15320
rect 38749 15317 38761 15320
rect 38795 15317 38807 15351
rect 38749 15311 38807 15317
rect 1104 15258 40572 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 40572 15258
rect 1104 15184 40572 15206
rect 4614 15104 4620 15156
rect 4672 15104 4678 15156
rect 5261 15147 5319 15153
rect 5261 15113 5273 15147
rect 5307 15144 5319 15147
rect 5534 15144 5540 15156
rect 5307 15116 5540 15144
rect 5307 15113 5319 15116
rect 5261 15107 5319 15113
rect 5534 15104 5540 15116
rect 5592 15104 5598 15156
rect 5718 15104 5724 15156
rect 5776 15144 5782 15156
rect 5776 15116 7328 15144
rect 5776 15104 5782 15116
rect 6733 15079 6791 15085
rect 4264 15048 6592 15076
rect 4264 15017 4292 15048
rect 4249 15011 4307 15017
rect 4249 14977 4261 15011
rect 4295 14977 4307 15011
rect 4249 14971 4307 14977
rect 5169 15011 5227 15017
rect 5169 14977 5181 15011
rect 5215 15008 5227 15011
rect 5258 15008 5264 15020
rect 5215 14980 5264 15008
rect 5215 14977 5227 14980
rect 5169 14971 5227 14977
rect 5258 14968 5264 14980
rect 5316 14968 5322 15020
rect 5353 15011 5411 15017
rect 5353 14977 5365 15011
rect 5399 14977 5411 15011
rect 5353 14971 5411 14977
rect 5813 15011 5871 15017
rect 5813 14977 5825 15011
rect 5859 15008 5871 15011
rect 5902 15008 5908 15020
rect 5859 14980 5908 15008
rect 5859 14977 5871 14980
rect 5813 14971 5871 14977
rect 4341 14943 4399 14949
rect 4341 14909 4353 14943
rect 4387 14940 4399 14943
rect 4614 14940 4620 14952
rect 4387 14912 4620 14940
rect 4387 14909 4399 14912
rect 4341 14903 4399 14909
rect 4614 14900 4620 14912
rect 4672 14900 4678 14952
rect 5368 14940 5396 14971
rect 5902 14968 5908 14980
rect 5960 14968 5966 15020
rect 5994 14968 6000 15020
rect 6052 14968 6058 15020
rect 6564 15017 6592 15048
rect 6733 15045 6745 15079
rect 6779 15076 6791 15079
rect 6822 15076 6828 15088
rect 6779 15048 6828 15076
rect 6779 15045 6791 15048
rect 6733 15039 6791 15045
rect 6822 15036 6828 15048
rect 6880 15036 6886 15088
rect 6917 15079 6975 15085
rect 6917 15045 6929 15079
rect 6963 15076 6975 15079
rect 7006 15076 7012 15088
rect 6963 15048 7012 15076
rect 6963 15045 6975 15048
rect 6917 15039 6975 15045
rect 7006 15036 7012 15048
rect 7064 15036 7070 15088
rect 6549 15011 6607 15017
rect 6549 14977 6561 15011
rect 6595 15008 6607 15011
rect 6595 14980 6960 15008
rect 6595 14977 6607 14980
rect 6549 14971 6607 14977
rect 6932 14952 6960 14980
rect 5368 14912 6684 14940
rect 6181 14807 6239 14813
rect 6181 14773 6193 14807
rect 6227 14804 6239 14807
rect 6454 14804 6460 14816
rect 6227 14776 6460 14804
rect 6227 14773 6239 14776
rect 6181 14767 6239 14773
rect 6454 14764 6460 14776
rect 6512 14764 6518 14816
rect 6656 14804 6684 14912
rect 6914 14900 6920 14952
rect 6972 14900 6978 14952
rect 7024 14940 7052 15036
rect 7193 14943 7251 14949
rect 7193 14940 7205 14943
rect 7024 14912 7205 14940
rect 7193 14909 7205 14912
rect 7239 14909 7251 14943
rect 7300 14940 7328 15116
rect 7834 15104 7840 15156
rect 7892 15144 7898 15156
rect 8478 15144 8484 15156
rect 7892 15116 8484 15144
rect 7892 15104 7898 15116
rect 8478 15104 8484 15116
rect 8536 15104 8542 15156
rect 8665 15147 8723 15153
rect 8665 15113 8677 15147
rect 8711 15144 8723 15147
rect 8938 15144 8944 15156
rect 8711 15116 8944 15144
rect 8711 15113 8723 15116
rect 8665 15107 8723 15113
rect 8680 15076 8708 15107
rect 8938 15104 8944 15116
rect 8996 15104 9002 15156
rect 10226 15144 10232 15156
rect 9140 15116 10232 15144
rect 7668 15048 8708 15076
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 15008 7435 15011
rect 7558 15008 7564 15020
rect 7423 14980 7564 15008
rect 7423 14977 7435 14980
rect 7377 14971 7435 14977
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 7668 15017 7696 15048
rect 7653 15011 7711 15017
rect 7653 14977 7665 15011
rect 7699 14977 7711 15011
rect 7653 14971 7711 14977
rect 7745 15011 7803 15017
rect 7745 14977 7757 15011
rect 7791 15008 7803 15011
rect 7926 15008 7932 15020
rect 7791 14980 7932 15008
rect 7791 14977 7803 14980
rect 7745 14971 7803 14977
rect 7926 14968 7932 14980
rect 7984 14968 7990 15020
rect 8018 14968 8024 15020
rect 8076 15008 8082 15020
rect 8297 15011 8355 15017
rect 8297 15008 8309 15011
rect 8076 14980 8309 15008
rect 8076 14968 8082 14980
rect 8297 14977 8309 14980
rect 8343 15008 8355 15011
rect 8570 15008 8576 15020
rect 8343 14980 8576 15008
rect 8343 14977 8355 14980
rect 8297 14971 8355 14977
rect 8570 14968 8576 14980
rect 8628 15008 8634 15020
rect 9140 15008 9168 15116
rect 10226 15104 10232 15116
rect 10284 15144 10290 15156
rect 10284 15116 12664 15144
rect 10284 15104 10290 15116
rect 9214 15036 9220 15088
rect 9272 15076 9278 15088
rect 12526 15076 12532 15088
rect 9272 15048 10088 15076
rect 9272 15036 9278 15048
rect 8628 14980 9168 15008
rect 8628 14968 8634 14980
rect 9398 14968 9404 15020
rect 9456 14968 9462 15020
rect 9677 15011 9735 15017
rect 9677 14977 9689 15011
rect 9723 15008 9735 15011
rect 9858 15008 9864 15020
rect 9723 14980 9864 15008
rect 9723 14977 9735 14980
rect 9677 14971 9735 14977
rect 9858 14968 9864 14980
rect 9916 14968 9922 15020
rect 10060 15017 10088 15048
rect 11992 15048 12532 15076
rect 10045 15011 10103 15017
rect 10045 14977 10057 15011
rect 10091 15008 10103 15011
rect 10091 14980 10732 15008
rect 10091 14977 10103 14980
rect 10045 14971 10103 14977
rect 7837 14943 7895 14949
rect 7837 14940 7849 14943
rect 7300 14912 7849 14940
rect 7193 14903 7251 14909
rect 7837 14909 7849 14912
rect 7883 14940 7895 14943
rect 8205 14943 8263 14949
rect 8205 14940 8217 14943
rect 7883 14912 8217 14940
rect 7883 14909 7895 14912
rect 7837 14903 7895 14909
rect 8205 14909 8217 14912
rect 8251 14940 8263 14943
rect 9309 14943 9367 14949
rect 8251 14912 9260 14940
rect 8251 14909 8263 14912
rect 8205 14903 8263 14909
rect 7006 14832 7012 14884
rect 7064 14832 7070 14884
rect 9125 14875 9183 14881
rect 9125 14872 9137 14875
rect 7116 14844 9137 14872
rect 7116 14804 7144 14844
rect 9125 14841 9137 14844
rect 9171 14841 9183 14875
rect 9125 14835 9183 14841
rect 6656 14776 7144 14804
rect 7190 14764 7196 14816
rect 7248 14764 7254 14816
rect 7282 14764 7288 14816
rect 7340 14764 7346 14816
rect 7466 14764 7472 14816
rect 7524 14764 7530 14816
rect 8021 14807 8079 14813
rect 8021 14773 8033 14807
rect 8067 14804 8079 14807
rect 8110 14804 8116 14816
rect 8067 14776 8116 14804
rect 8067 14773 8079 14776
rect 8021 14767 8079 14773
rect 8110 14764 8116 14776
rect 8168 14764 8174 14816
rect 9232 14804 9260 14912
rect 9309 14909 9321 14943
rect 9355 14909 9367 14943
rect 9309 14903 9367 14909
rect 9324 14872 9352 14903
rect 9490 14900 9496 14952
rect 9548 14940 9554 14952
rect 9769 14943 9827 14949
rect 9769 14940 9781 14943
rect 9548 14912 9781 14940
rect 9548 14900 9554 14912
rect 9769 14909 9781 14912
rect 9815 14909 9827 14943
rect 10137 14943 10195 14949
rect 10137 14940 10149 14943
rect 9769 14903 9827 14909
rect 9968 14912 10149 14940
rect 9861 14875 9919 14881
rect 9861 14872 9873 14875
rect 9324 14844 9873 14872
rect 9861 14841 9873 14844
rect 9907 14841 9919 14875
rect 9861 14835 9919 14841
rect 9968 14804 9996 14912
rect 10137 14909 10149 14912
rect 10183 14909 10195 14943
rect 10137 14903 10195 14909
rect 10226 14900 10232 14952
rect 10284 14900 10290 14952
rect 10318 14900 10324 14952
rect 10376 14900 10382 14952
rect 10704 14940 10732 14980
rect 10778 14968 10784 15020
rect 10836 14968 10842 15020
rect 11885 15011 11943 15017
rect 11885 14977 11897 15011
rect 11931 14977 11943 15011
rect 11885 14971 11943 14977
rect 11606 14940 11612 14952
rect 10704 14912 11612 14940
rect 11606 14900 11612 14912
rect 11664 14940 11670 14952
rect 11793 14943 11851 14949
rect 11793 14940 11805 14943
rect 11664 14912 11805 14940
rect 11664 14900 11670 14912
rect 11793 14909 11805 14912
rect 11839 14909 11851 14943
rect 11793 14903 11851 14909
rect 10597 14875 10655 14881
rect 10597 14872 10609 14875
rect 10152 14844 10609 14872
rect 10152 14816 10180 14844
rect 10597 14841 10609 14844
rect 10643 14841 10655 14875
rect 11900 14872 11928 14971
rect 11992 14949 12020 15048
rect 12526 15036 12532 15048
rect 12584 15036 12590 15088
rect 12636 15076 12664 15116
rect 13354 15104 13360 15156
rect 13412 15144 13418 15156
rect 13817 15147 13875 15153
rect 13817 15144 13829 15147
rect 13412 15116 13829 15144
rect 13412 15104 13418 15116
rect 13817 15113 13829 15116
rect 13863 15113 13875 15147
rect 20533 15147 20591 15153
rect 13817 15107 13875 15113
rect 13924 15116 20300 15144
rect 13372 15076 13400 15104
rect 12636 15048 13400 15076
rect 12434 14968 12440 15020
rect 12492 14968 12498 15020
rect 12636 15017 12664 15048
rect 13446 15036 13452 15088
rect 13504 15076 13510 15088
rect 13924 15076 13952 15116
rect 13504 15048 13952 15076
rect 13504 15036 13510 15048
rect 16758 15036 16764 15088
rect 16816 15076 16822 15088
rect 17313 15079 17371 15085
rect 17313 15076 17325 15079
rect 16816 15048 17325 15076
rect 16816 15036 16822 15048
rect 17313 15045 17325 15048
rect 17359 15076 17371 15079
rect 17494 15076 17500 15088
rect 17359 15048 17500 15076
rect 17359 15045 17371 15048
rect 17313 15039 17371 15045
rect 17494 15036 17500 15048
rect 17552 15036 17558 15088
rect 17862 15036 17868 15088
rect 17920 15036 17926 15088
rect 18138 15036 18144 15088
rect 18196 15076 18202 15088
rect 18196 15048 20116 15076
rect 18196 15036 18202 15048
rect 12621 15011 12679 15017
rect 12621 14977 12633 15011
rect 12667 14977 12679 15011
rect 12621 14971 12679 14977
rect 12710 14968 12716 15020
rect 12768 14968 12774 15020
rect 12894 14968 12900 15020
rect 12952 15008 12958 15020
rect 13081 15011 13139 15017
rect 13081 15008 13093 15011
rect 12952 14980 13093 15008
rect 12952 14968 12958 14980
rect 13081 14977 13093 14980
rect 13127 14977 13139 15011
rect 13081 14971 13139 14977
rect 13170 14968 13176 15020
rect 13228 14968 13234 15020
rect 13262 14968 13268 15020
rect 13320 15008 13326 15020
rect 13541 15011 13599 15017
rect 13541 15008 13553 15011
rect 13320 14980 13553 15008
rect 13320 14968 13326 14980
rect 13541 14977 13553 14980
rect 13587 15008 13599 15011
rect 14185 15011 14243 15017
rect 14185 15008 14197 15011
rect 13587 14980 14197 15008
rect 13587 14977 13599 14980
rect 13541 14971 13599 14977
rect 14185 14977 14197 14980
rect 14231 14977 14243 15011
rect 14185 14971 14243 14977
rect 14921 15011 14979 15017
rect 14921 14977 14933 15011
rect 14967 14977 14979 15011
rect 14921 14971 14979 14977
rect 11977 14943 12035 14949
rect 11977 14909 11989 14943
rect 12023 14909 12035 14943
rect 11977 14903 12035 14909
rect 12066 14900 12072 14952
rect 12124 14900 12130 14952
rect 12912 14940 12940 14968
rect 12406 14912 12940 14940
rect 14936 14940 14964 14971
rect 15102 14968 15108 15020
rect 15160 15008 15166 15020
rect 15381 15011 15439 15017
rect 15381 15008 15393 15011
rect 15160 14980 15393 15008
rect 15160 14968 15166 14980
rect 15381 14977 15393 14980
rect 15427 14977 15439 15011
rect 15381 14971 15439 14977
rect 15838 14968 15844 15020
rect 15896 14968 15902 15020
rect 16301 15011 16359 15017
rect 16301 14977 16313 15011
rect 16347 15008 16359 15011
rect 16482 15008 16488 15020
rect 16347 14980 16488 15008
rect 16347 14977 16359 14980
rect 16301 14971 16359 14977
rect 16482 14968 16488 14980
rect 16540 14968 16546 15020
rect 16850 14968 16856 15020
rect 16908 14968 16914 15020
rect 17589 15011 17647 15017
rect 17589 14977 17601 15011
rect 17635 15008 17647 15011
rect 19334 15008 19340 15020
rect 17635 14980 19340 15008
rect 17635 14977 17647 14980
rect 17589 14971 17647 14977
rect 19334 14968 19340 14980
rect 19392 14968 19398 15020
rect 19610 14968 19616 15020
rect 19668 15008 19674 15020
rect 19705 15011 19763 15017
rect 19705 15008 19717 15011
rect 19668 14980 19717 15008
rect 19668 14968 19674 14980
rect 19705 14977 19717 14980
rect 19751 14977 19763 15011
rect 19705 14971 19763 14977
rect 19794 14968 19800 15020
rect 19852 14968 19858 15020
rect 19978 14968 19984 15020
rect 20036 14968 20042 15020
rect 20088 15017 20116 15048
rect 20162 15036 20168 15088
rect 20220 15036 20226 15088
rect 20073 15011 20131 15017
rect 20073 14977 20085 15011
rect 20119 14977 20131 15011
rect 20272 15008 20300 15116
rect 20533 15113 20545 15147
rect 20579 15144 20591 15147
rect 20622 15144 20628 15156
rect 20579 15116 20628 15144
rect 20579 15113 20591 15116
rect 20533 15107 20591 15113
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 22646 15104 22652 15156
rect 22704 15144 22710 15156
rect 22741 15147 22799 15153
rect 22741 15144 22753 15147
rect 22704 15116 22753 15144
rect 22704 15104 22710 15116
rect 22741 15113 22753 15116
rect 22787 15144 22799 15147
rect 23106 15144 23112 15156
rect 22787 15116 23112 15144
rect 22787 15113 22799 15116
rect 22741 15107 22799 15113
rect 23106 15104 23112 15116
rect 23164 15104 23170 15156
rect 24581 15147 24639 15153
rect 24581 15113 24593 15147
rect 24627 15144 24639 15147
rect 24670 15144 24676 15156
rect 24627 15116 24676 15144
rect 24627 15113 24639 15116
rect 24581 15107 24639 15113
rect 24670 15104 24676 15116
rect 24728 15104 24734 15156
rect 24780 15116 28994 15144
rect 20381 15079 20439 15085
rect 20381 15045 20393 15079
rect 20427 15076 20439 15079
rect 21266 15076 21272 15088
rect 20427 15048 21272 15076
rect 20427 15045 20439 15048
rect 20381 15039 20439 15045
rect 21266 15036 21272 15048
rect 21324 15076 21330 15088
rect 21542 15076 21548 15088
rect 21324 15048 21548 15076
rect 21324 15036 21330 15048
rect 21542 15036 21548 15048
rect 21600 15036 21606 15088
rect 24780 15076 24808 15116
rect 25130 15076 25136 15088
rect 24136 15048 24808 15076
rect 24872 15048 25136 15076
rect 20272 14980 22232 15008
rect 20073 14971 20131 14977
rect 14936 14912 16712 14940
rect 12406 14872 12434 14912
rect 11900 14844 12434 14872
rect 12912 14872 12940 14912
rect 12912 14844 13860 14872
rect 10597 14835 10655 14841
rect 9232 14776 9996 14804
rect 10134 14764 10140 14816
rect 10192 14764 10198 14816
rect 11609 14807 11667 14813
rect 11609 14773 11621 14807
rect 11655 14804 11667 14807
rect 11698 14804 11704 14816
rect 11655 14776 11704 14804
rect 11655 14773 11667 14776
rect 11609 14767 11667 14773
rect 11698 14764 11704 14776
rect 11756 14764 11762 14816
rect 12894 14764 12900 14816
rect 12952 14764 12958 14816
rect 13630 14764 13636 14816
rect 13688 14764 13694 14816
rect 13832 14813 13860 14844
rect 14826 14832 14832 14884
rect 14884 14872 14890 14884
rect 16684 14881 16712 14912
rect 15381 14875 15439 14881
rect 15381 14872 15393 14875
rect 14884 14844 15393 14872
rect 14884 14832 14890 14844
rect 15381 14841 15393 14844
rect 15427 14841 15439 14875
rect 15381 14835 15439 14841
rect 16669 14875 16727 14881
rect 16669 14841 16681 14875
rect 16715 14841 16727 14875
rect 16868 14872 16896 14968
rect 17034 14900 17040 14952
rect 17092 14900 17098 14952
rect 17773 14943 17831 14949
rect 17773 14909 17785 14943
rect 17819 14940 17831 14943
rect 17954 14940 17960 14952
rect 17819 14912 17960 14940
rect 17819 14909 17831 14912
rect 17773 14903 17831 14909
rect 17954 14900 17960 14912
rect 18012 14900 18018 14952
rect 19812 14940 19840 14968
rect 20438 14940 20444 14952
rect 19812 14912 20444 14940
rect 20438 14900 20444 14912
rect 20496 14940 20502 14952
rect 21266 14940 21272 14952
rect 20496 14912 21272 14940
rect 20496 14900 20502 14912
rect 21266 14900 21272 14912
rect 21324 14900 21330 14952
rect 17405 14875 17463 14881
rect 17405 14872 17417 14875
rect 16868 14844 17417 14872
rect 16669 14835 16727 14841
rect 17405 14841 17417 14844
rect 17451 14841 17463 14875
rect 17405 14835 17463 14841
rect 18690 14832 18696 14884
rect 18748 14872 18754 14884
rect 21174 14872 21180 14884
rect 18748 14844 21180 14872
rect 18748 14832 18754 14844
rect 21174 14832 21180 14844
rect 21232 14832 21238 14884
rect 22204 14872 22232 14980
rect 22278 14968 22284 15020
rect 22336 15008 22342 15020
rect 22465 15011 22523 15017
rect 22465 15008 22477 15011
rect 22336 14980 22477 15008
rect 22336 14968 22342 14980
rect 22465 14977 22477 14980
rect 22511 14977 22523 15011
rect 22465 14971 22523 14977
rect 22830 14968 22836 15020
rect 22888 15008 22894 15020
rect 24136 15008 24164 15048
rect 22888 14980 24164 15008
rect 22888 14968 22894 14980
rect 24210 14968 24216 15020
rect 24268 15008 24274 15020
rect 24268 14980 24532 15008
rect 24268 14968 24274 14980
rect 24504 14952 24532 14980
rect 24670 14968 24676 15020
rect 24728 15014 24734 15020
rect 24872 15017 24900 15048
rect 25130 15036 25136 15048
rect 25188 15036 25194 15088
rect 28966 15076 28994 15116
rect 31018 15104 31024 15156
rect 31076 15144 31082 15156
rect 31754 15144 31760 15156
rect 31076 15116 31760 15144
rect 31076 15104 31082 15116
rect 31754 15104 31760 15116
rect 31812 15144 31818 15156
rect 33962 15144 33968 15156
rect 31812 15116 33968 15144
rect 31812 15104 31818 15116
rect 33962 15104 33968 15116
rect 34020 15104 34026 15156
rect 34425 15147 34483 15153
rect 34425 15113 34437 15147
rect 34471 15144 34483 15147
rect 34974 15144 34980 15156
rect 34471 15116 34980 15144
rect 34471 15113 34483 15116
rect 34425 15107 34483 15113
rect 34974 15104 34980 15116
rect 35032 15144 35038 15156
rect 35032 15116 35940 15144
rect 35032 15104 35038 15116
rect 30282 15076 30288 15088
rect 28966 15048 30288 15076
rect 30282 15036 30288 15048
rect 30340 15036 30346 15088
rect 33134 15036 33140 15088
rect 33192 15076 33198 15088
rect 34149 15079 34207 15085
rect 34149 15076 34161 15079
rect 33192 15048 34161 15076
rect 33192 15036 33198 15048
rect 34149 15045 34161 15048
rect 34195 15045 34207 15079
rect 34149 15039 34207 15045
rect 35434 15036 35440 15088
rect 35492 15076 35498 15088
rect 35912 15085 35940 15116
rect 38470 15104 38476 15156
rect 38528 15144 38534 15156
rect 39022 15144 39028 15156
rect 38528 15116 39028 15144
rect 38528 15104 38534 15116
rect 39022 15104 39028 15116
rect 39080 15104 39086 15156
rect 35713 15079 35771 15085
rect 35713 15076 35725 15079
rect 35492 15048 35725 15076
rect 35492 15036 35498 15048
rect 35713 15045 35725 15048
rect 35759 15045 35771 15079
rect 35713 15039 35771 15045
rect 35897 15079 35955 15085
rect 35897 15045 35909 15079
rect 35943 15045 35955 15079
rect 35897 15039 35955 15045
rect 24765 15014 24823 15017
rect 24728 15011 24823 15014
rect 24728 14986 24777 15011
rect 24728 14968 24734 14986
rect 24765 14977 24777 14986
rect 24811 14977 24823 15011
rect 24765 14971 24823 14977
rect 24857 15011 24915 15017
rect 24857 14977 24869 15011
rect 24903 14977 24915 15011
rect 24857 14971 24915 14977
rect 25041 15011 25099 15017
rect 25041 14977 25053 15011
rect 25087 15008 25099 15011
rect 28994 15008 29000 15020
rect 25087 14980 29000 15008
rect 25087 14977 25099 14980
rect 25041 14971 25099 14977
rect 22373 14943 22431 14949
rect 22373 14909 22385 14943
rect 22419 14940 22431 14943
rect 22646 14940 22652 14952
rect 22419 14912 22652 14940
rect 22419 14909 22431 14912
rect 22373 14903 22431 14909
rect 22646 14900 22652 14912
rect 22704 14940 22710 14952
rect 24394 14940 24400 14952
rect 22704 14912 24400 14940
rect 22704 14900 22710 14912
rect 24394 14900 24400 14912
rect 24452 14900 24458 14952
rect 24486 14900 24492 14952
rect 24544 14940 24550 14952
rect 25056 14940 25084 14971
rect 28994 14968 29000 14980
rect 29052 14968 29058 15020
rect 33873 15011 33931 15017
rect 33873 14977 33885 15011
rect 33919 14977 33931 15011
rect 33873 14971 33931 14977
rect 24544 14912 25084 14940
rect 24544 14900 24550 14912
rect 31478 14900 31484 14952
rect 31536 14940 31542 14952
rect 33888 14940 33916 14971
rect 33962 14968 33968 15020
rect 34020 15008 34026 15020
rect 34057 15011 34115 15017
rect 34057 15008 34069 15011
rect 34020 14980 34069 15008
rect 34020 14968 34026 14980
rect 34057 14977 34069 14980
rect 34103 14977 34115 15011
rect 34057 14971 34115 14977
rect 34241 15011 34299 15017
rect 34241 14977 34253 15011
rect 34287 15008 34299 15011
rect 35342 15008 35348 15020
rect 34287 14980 35348 15008
rect 34287 14977 34299 14980
rect 34241 14971 34299 14977
rect 35342 14968 35348 14980
rect 35400 14968 35406 15020
rect 38654 14968 38660 15020
rect 38712 14968 38718 15020
rect 38838 14968 38844 15020
rect 38896 14968 38902 15020
rect 34606 14940 34612 14952
rect 31536 14912 34612 14940
rect 31536 14900 31542 14912
rect 34606 14900 34612 14912
rect 34664 14900 34670 14952
rect 24670 14872 24676 14884
rect 22204 14844 24676 14872
rect 24670 14832 24676 14844
rect 24728 14832 24734 14884
rect 24949 14875 25007 14881
rect 24949 14841 24961 14875
rect 24995 14872 25007 14875
rect 27706 14872 27712 14884
rect 24995 14844 27712 14872
rect 24995 14841 25007 14844
rect 24949 14835 25007 14841
rect 27706 14832 27712 14844
rect 27764 14832 27770 14884
rect 33318 14832 33324 14884
rect 33376 14872 33382 14884
rect 37550 14872 37556 14884
rect 33376 14844 37556 14872
rect 33376 14832 33382 14844
rect 37550 14832 37556 14844
rect 37608 14832 37614 14884
rect 13817 14807 13875 14813
rect 13817 14773 13829 14807
rect 13863 14773 13875 14807
rect 13817 14767 13875 14773
rect 14734 14764 14740 14816
rect 14792 14764 14798 14816
rect 16482 14764 16488 14816
rect 16540 14804 16546 14816
rect 16853 14807 16911 14813
rect 16853 14804 16865 14807
rect 16540 14776 16865 14804
rect 16540 14764 16546 14776
rect 16853 14773 16865 14776
rect 16899 14773 16911 14807
rect 16853 14767 16911 14773
rect 17770 14764 17776 14816
rect 17828 14764 17834 14816
rect 19518 14764 19524 14816
rect 19576 14764 19582 14816
rect 20349 14807 20407 14813
rect 20349 14773 20361 14807
rect 20395 14804 20407 14807
rect 20714 14804 20720 14816
rect 20395 14776 20720 14804
rect 20395 14773 20407 14776
rect 20349 14767 20407 14773
rect 20714 14764 20720 14776
rect 20772 14764 20778 14816
rect 20806 14764 20812 14816
rect 20864 14804 20870 14816
rect 22097 14807 22155 14813
rect 22097 14804 22109 14807
rect 20864 14776 22109 14804
rect 20864 14764 20870 14776
rect 22097 14773 22109 14776
rect 22143 14773 22155 14807
rect 22097 14767 22155 14773
rect 22557 14807 22615 14813
rect 22557 14773 22569 14807
rect 22603 14804 22615 14807
rect 22922 14804 22928 14816
rect 22603 14776 22928 14804
rect 22603 14773 22615 14776
rect 22557 14767 22615 14773
rect 22922 14764 22928 14776
rect 22980 14804 22986 14816
rect 24394 14804 24400 14816
rect 22980 14776 24400 14804
rect 22980 14764 22986 14776
rect 24394 14764 24400 14776
rect 24452 14764 24458 14816
rect 34054 14764 34060 14816
rect 34112 14804 34118 14816
rect 34422 14804 34428 14816
rect 34112 14776 34428 14804
rect 34112 14764 34118 14776
rect 34422 14764 34428 14776
rect 34480 14764 34486 14816
rect 36081 14807 36139 14813
rect 36081 14773 36093 14807
rect 36127 14804 36139 14807
rect 38654 14804 38660 14816
rect 36127 14776 38660 14804
rect 36127 14773 36139 14776
rect 36081 14767 36139 14773
rect 38654 14764 38660 14776
rect 38712 14764 38718 14816
rect 39022 14764 39028 14816
rect 39080 14764 39086 14816
rect 1104 14714 40572 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 40572 14714
rect 1104 14640 40572 14662
rect 4525 14603 4583 14609
rect 4525 14569 4537 14603
rect 4571 14600 4583 14603
rect 5810 14600 5816 14612
rect 4571 14572 5816 14600
rect 4571 14569 4583 14572
rect 4525 14563 4583 14569
rect 5810 14560 5816 14572
rect 5868 14560 5874 14612
rect 6270 14560 6276 14612
rect 6328 14560 6334 14612
rect 7006 14560 7012 14612
rect 7064 14600 7070 14612
rect 9309 14603 9367 14609
rect 7064 14572 9260 14600
rect 7064 14560 7070 14572
rect 4614 14492 4620 14544
rect 4672 14492 4678 14544
rect 6181 14535 6239 14541
rect 6181 14501 6193 14535
rect 6227 14501 6239 14535
rect 7837 14535 7895 14541
rect 7837 14532 7849 14535
rect 6181 14495 6239 14501
rect 6748 14504 7849 14532
rect 4246 14424 4252 14476
rect 4304 14424 4310 14476
rect 6196 14464 6224 14495
rect 6104 14436 6224 14464
rect 4157 14399 4215 14405
rect 4157 14365 4169 14399
rect 4203 14396 4215 14399
rect 4338 14396 4344 14408
rect 4203 14368 4344 14396
rect 4203 14365 4215 14368
rect 4157 14359 4215 14365
rect 4338 14356 4344 14368
rect 4396 14356 4402 14408
rect 4706 14356 4712 14408
rect 4764 14396 4770 14408
rect 4831 14399 4889 14405
rect 4831 14396 4843 14399
rect 4764 14368 4843 14396
rect 4764 14356 4770 14368
rect 4831 14365 4843 14368
rect 4877 14365 4889 14399
rect 4831 14359 4889 14365
rect 4985 14399 5043 14405
rect 4985 14365 4997 14399
rect 5031 14396 5043 14399
rect 5902 14396 5908 14408
rect 5031 14368 5908 14396
rect 5031 14365 5043 14368
rect 4985 14359 5043 14365
rect 5902 14356 5908 14368
rect 5960 14356 5966 14408
rect 5994 14220 6000 14272
rect 6052 14220 6058 14272
rect 6104 14260 6132 14436
rect 6454 14424 6460 14476
rect 6512 14424 6518 14476
rect 6546 14424 6552 14476
rect 6604 14424 6610 14476
rect 6748 14473 6776 14504
rect 7837 14501 7849 14504
rect 7883 14501 7895 14535
rect 9122 14532 9128 14544
rect 7837 14495 7895 14501
rect 8358 14504 9128 14532
rect 6733 14467 6791 14473
rect 6733 14433 6745 14467
rect 6779 14433 6791 14467
rect 6733 14427 6791 14433
rect 6822 14424 6828 14476
rect 6880 14464 6886 14476
rect 7558 14464 7564 14476
rect 6880 14436 7328 14464
rect 6880 14424 6886 14436
rect 6641 14399 6699 14405
rect 6641 14365 6653 14399
rect 6687 14396 6699 14399
rect 7098 14396 7104 14408
rect 6687 14368 7104 14396
rect 6687 14365 6699 14368
rect 6641 14359 6699 14365
rect 7098 14356 7104 14368
rect 7156 14356 7162 14408
rect 7190 14356 7196 14408
rect 7248 14356 7254 14408
rect 7300 14405 7328 14436
rect 7484 14436 7564 14464
rect 7484 14405 7512 14436
rect 7558 14424 7564 14436
rect 7616 14424 7622 14476
rect 8358 14430 8386 14504
rect 9122 14492 9128 14504
rect 9180 14492 9186 14544
rect 9232 14532 9260 14572
rect 9309 14569 9321 14603
rect 9355 14600 9367 14603
rect 9398 14600 9404 14612
rect 9355 14572 9404 14600
rect 9355 14569 9367 14572
rect 9309 14563 9367 14569
rect 9398 14560 9404 14572
rect 9456 14560 9462 14612
rect 9490 14560 9496 14612
rect 9548 14600 9554 14612
rect 9950 14600 9956 14612
rect 9548 14572 9956 14600
rect 9548 14560 9554 14572
rect 9950 14560 9956 14572
rect 10008 14600 10014 14612
rect 10134 14600 10140 14612
rect 10008 14572 10140 14600
rect 10008 14560 10014 14572
rect 10134 14560 10140 14572
rect 10192 14560 10198 14612
rect 10229 14603 10287 14609
rect 10229 14569 10241 14603
rect 10275 14600 10287 14603
rect 10318 14600 10324 14612
rect 10275 14572 10324 14600
rect 10275 14569 10287 14572
rect 10229 14563 10287 14569
rect 10318 14560 10324 14572
rect 10376 14560 10382 14612
rect 10778 14560 10784 14612
rect 10836 14600 10842 14612
rect 14734 14600 14740 14612
rect 10836 14572 14740 14600
rect 10836 14560 10842 14572
rect 14734 14560 14740 14572
rect 14792 14560 14798 14612
rect 15654 14560 15660 14612
rect 15712 14560 15718 14612
rect 15838 14560 15844 14612
rect 15896 14560 15902 14612
rect 16022 14560 16028 14612
rect 16080 14560 16086 14612
rect 17405 14603 17463 14609
rect 17405 14569 17417 14603
rect 17451 14600 17463 14603
rect 17954 14600 17960 14612
rect 17451 14572 17960 14600
rect 17451 14569 17463 14572
rect 17405 14563 17463 14569
rect 17954 14560 17960 14572
rect 18012 14560 18018 14612
rect 18230 14560 18236 14612
rect 18288 14600 18294 14612
rect 18874 14600 18880 14612
rect 18288 14572 18880 14600
rect 18288 14560 18294 14572
rect 18874 14560 18880 14572
rect 18932 14560 18938 14612
rect 19518 14560 19524 14612
rect 19576 14560 19582 14612
rect 19794 14560 19800 14612
rect 19852 14560 19858 14612
rect 20349 14603 20407 14609
rect 20349 14569 20361 14603
rect 20395 14600 20407 14603
rect 20622 14600 20628 14612
rect 20395 14572 20628 14600
rect 20395 14569 20407 14572
rect 20349 14563 20407 14569
rect 20622 14560 20628 14572
rect 20680 14560 20686 14612
rect 20993 14603 21051 14609
rect 20993 14569 21005 14603
rect 21039 14600 21051 14603
rect 21039 14572 22140 14600
rect 21039 14569 21051 14572
rect 20993 14563 21051 14569
rect 14921 14535 14979 14541
rect 14921 14532 14933 14535
rect 9232 14504 14933 14532
rect 8358 14405 8412 14430
rect 8754 14424 8760 14476
rect 8812 14464 8818 14476
rect 10134 14464 10140 14476
rect 8812 14436 9720 14464
rect 8812 14424 8818 14436
rect 9692 14408 9720 14436
rect 9876 14436 10140 14464
rect 7286 14399 7344 14405
rect 7286 14365 7298 14399
rect 7332 14365 7344 14399
rect 7286 14359 7344 14365
rect 7469 14399 7527 14405
rect 7469 14365 7481 14399
rect 7515 14365 7527 14399
rect 7469 14359 7527 14365
rect 7699 14399 7757 14405
rect 8358 14402 8447 14405
rect 7699 14365 7711 14399
rect 7745 14365 7757 14399
rect 8384 14399 8447 14402
rect 8384 14368 8401 14399
rect 7699 14359 7757 14365
rect 8389 14365 8401 14368
rect 8435 14365 8447 14399
rect 8389 14359 8447 14365
rect 6181 14331 6239 14337
rect 6181 14297 6193 14331
rect 6227 14328 6239 14331
rect 6822 14328 6828 14340
rect 6227 14300 6828 14328
rect 6227 14297 6239 14300
rect 6181 14291 6239 14297
rect 6822 14288 6828 14300
rect 6880 14288 6886 14340
rect 7558 14288 7564 14340
rect 7616 14288 7622 14340
rect 7714 14328 7742 14359
rect 8478 14356 8484 14408
rect 8536 14356 8542 14408
rect 8570 14356 8576 14408
rect 8628 14356 8634 14408
rect 8662 14356 8668 14408
rect 8720 14356 8726 14408
rect 9490 14405 9496 14408
rect 9488 14396 9496 14405
rect 9451 14368 9496 14396
rect 9488 14359 9496 14368
rect 9490 14356 9496 14359
rect 9548 14356 9554 14408
rect 9674 14356 9680 14408
rect 9732 14356 9738 14408
rect 9876 14405 9904 14436
rect 10134 14424 10140 14436
rect 10192 14424 10198 14476
rect 9860 14399 9918 14405
rect 9860 14365 9872 14399
rect 9906 14365 9918 14399
rect 9860 14359 9918 14365
rect 9950 14356 9956 14408
rect 10008 14356 10014 14408
rect 10042 14356 10048 14408
rect 10100 14356 10106 14408
rect 10244 14405 10272 14504
rect 14921 14501 14933 14504
rect 14967 14501 14979 14535
rect 14921 14495 14979 14501
rect 15289 14535 15347 14541
rect 15289 14501 15301 14535
rect 15335 14532 15347 14535
rect 15746 14532 15752 14544
rect 15335 14504 15752 14532
rect 15335 14501 15347 14504
rect 15289 14495 15347 14501
rect 15746 14492 15752 14504
rect 15804 14492 15810 14544
rect 15930 14492 15936 14544
rect 15988 14532 15994 14544
rect 20162 14532 20168 14544
rect 15988 14504 20168 14532
rect 15988 14492 15994 14504
rect 16117 14467 16175 14473
rect 15028 14436 15608 14464
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14365 10287 14399
rect 10229 14359 10287 14365
rect 10321 14399 10379 14405
rect 10321 14365 10333 14399
rect 10367 14365 10379 14399
rect 10321 14359 10379 14365
rect 9503 14328 9531 14356
rect 7714 14300 9531 14328
rect 9585 14331 9643 14337
rect 9585 14297 9597 14331
rect 9631 14328 9643 14331
rect 10060 14328 10088 14356
rect 10336 14328 10364 14359
rect 10410 14356 10416 14408
rect 10468 14396 10474 14408
rect 10505 14399 10563 14405
rect 10505 14396 10517 14399
rect 10468 14368 10517 14396
rect 10468 14356 10474 14368
rect 10505 14365 10517 14368
rect 10551 14365 10563 14399
rect 10505 14359 10563 14365
rect 11606 14356 11612 14408
rect 11664 14396 11670 14408
rect 15028 14405 15056 14436
rect 15580 14408 15608 14436
rect 16117 14433 16129 14467
rect 16163 14464 16175 14467
rect 16850 14464 16856 14476
rect 16163 14436 16856 14464
rect 16163 14433 16175 14436
rect 16117 14427 16175 14433
rect 16850 14424 16856 14436
rect 16908 14424 16914 14476
rect 17221 14467 17279 14473
rect 17221 14433 17233 14467
rect 17267 14464 17279 14467
rect 17586 14464 17592 14476
rect 17267 14436 17592 14464
rect 17267 14433 17279 14436
rect 17221 14427 17279 14433
rect 17586 14424 17592 14436
rect 17644 14424 17650 14476
rect 18690 14424 18696 14476
rect 18748 14424 18754 14476
rect 18874 14424 18880 14476
rect 18932 14424 18938 14476
rect 18984 14473 19012 14504
rect 20162 14492 20168 14504
rect 20220 14492 20226 14544
rect 20809 14535 20867 14541
rect 20809 14501 20821 14535
rect 20855 14532 20867 14535
rect 20855 14504 21312 14532
rect 20855 14501 20867 14504
rect 20809 14495 20867 14501
rect 18969 14467 19027 14473
rect 18969 14433 18981 14467
rect 19015 14433 19027 14467
rect 18969 14427 19027 14433
rect 19521 14467 19579 14473
rect 19521 14433 19533 14467
rect 19567 14464 19579 14467
rect 19794 14464 19800 14476
rect 19567 14436 19800 14464
rect 19567 14433 19579 14436
rect 19521 14427 19579 14433
rect 19794 14424 19800 14436
rect 19852 14424 19858 14476
rect 20441 14467 20499 14473
rect 20441 14433 20453 14467
rect 20487 14464 20499 14467
rect 20824 14464 20852 14495
rect 20487 14436 20852 14464
rect 20487 14433 20499 14436
rect 20441 14427 20499 14433
rect 21174 14424 21180 14476
rect 21232 14424 21238 14476
rect 12529 14399 12587 14405
rect 12529 14396 12541 14399
rect 11664 14368 12541 14396
rect 11664 14356 11670 14368
rect 12529 14365 12541 14368
rect 12575 14365 12587 14399
rect 12529 14359 12587 14365
rect 14829 14399 14887 14405
rect 14829 14365 14841 14399
rect 14875 14365 14887 14399
rect 14829 14359 14887 14365
rect 15013 14399 15071 14405
rect 15013 14365 15025 14399
rect 15059 14365 15071 14399
rect 15013 14359 15071 14365
rect 15473 14399 15531 14405
rect 15473 14365 15485 14399
rect 15519 14365 15531 14399
rect 15473 14359 15531 14365
rect 9631 14300 9812 14328
rect 10060 14300 10364 14328
rect 9631 14297 9643 14300
rect 9585 14291 9643 14297
rect 7374 14260 7380 14272
rect 6104 14232 7380 14260
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 8202 14220 8208 14272
rect 8260 14220 8266 14272
rect 8662 14220 8668 14272
rect 8720 14260 8726 14272
rect 9398 14260 9404 14272
rect 8720 14232 9404 14260
rect 8720 14220 8726 14232
rect 9398 14220 9404 14232
rect 9456 14220 9462 14272
rect 9784 14260 9812 14300
rect 12986 14288 12992 14340
rect 13044 14328 13050 14340
rect 14844 14328 14872 14359
rect 15286 14328 15292 14340
rect 13044 14300 13308 14328
rect 14844 14300 15292 14328
rect 13044 14288 13050 14300
rect 10410 14260 10416 14272
rect 9784 14232 10416 14260
rect 10410 14220 10416 14232
rect 10468 14220 10474 14272
rect 11882 14220 11888 14272
rect 11940 14260 11946 14272
rect 12066 14260 12072 14272
rect 11940 14232 12072 14260
rect 11940 14220 11946 14232
rect 12066 14220 12072 14232
rect 12124 14220 12130 14272
rect 12621 14263 12679 14269
rect 12621 14229 12633 14263
rect 12667 14260 12679 14263
rect 13170 14260 13176 14272
rect 12667 14232 13176 14260
rect 12667 14229 12679 14232
rect 12621 14223 12679 14229
rect 13170 14220 13176 14232
rect 13228 14220 13234 14272
rect 13280 14260 13308 14300
rect 15286 14288 15292 14300
rect 15344 14288 15350 14340
rect 15488 14328 15516 14359
rect 15562 14356 15568 14408
rect 15620 14356 15626 14408
rect 15930 14396 15936 14408
rect 15672 14368 15936 14396
rect 15672 14328 15700 14368
rect 15930 14356 15936 14368
rect 15988 14356 15994 14408
rect 16393 14399 16451 14405
rect 16393 14365 16405 14399
rect 16439 14396 16451 14399
rect 16758 14396 16764 14408
rect 16439 14368 16764 14396
rect 16439 14365 16451 14368
rect 16393 14359 16451 14365
rect 16758 14356 16764 14368
rect 16816 14356 16822 14408
rect 17129 14399 17187 14405
rect 17129 14365 17141 14399
rect 17175 14365 17187 14399
rect 17129 14359 17187 14365
rect 15488 14300 15700 14328
rect 15749 14331 15807 14337
rect 15749 14297 15761 14331
rect 15795 14328 15807 14331
rect 17144 14328 17172 14359
rect 17310 14356 17316 14408
rect 17368 14396 17374 14408
rect 17405 14399 17463 14405
rect 17405 14396 17417 14399
rect 17368 14368 17417 14396
rect 17368 14356 17374 14368
rect 17405 14365 17417 14368
rect 17451 14365 17463 14399
rect 17405 14359 17463 14365
rect 18785 14399 18843 14405
rect 18785 14365 18797 14399
rect 18831 14365 18843 14399
rect 18785 14359 18843 14365
rect 18800 14328 18828 14359
rect 19610 14356 19616 14408
rect 19668 14356 19674 14408
rect 20162 14356 20168 14408
rect 20220 14396 20226 14408
rect 20257 14399 20315 14405
rect 20257 14396 20269 14399
rect 20220 14368 20269 14396
rect 20220 14356 20226 14368
rect 20257 14365 20269 14368
rect 20303 14365 20315 14399
rect 20257 14359 20315 14365
rect 20530 14356 20536 14408
rect 20588 14356 20594 14408
rect 20717 14399 20775 14405
rect 20717 14365 20729 14399
rect 20763 14365 20775 14399
rect 21192 14396 21220 14424
rect 20717 14359 20775 14365
rect 21100 14368 21220 14396
rect 21284 14396 21312 14504
rect 21726 14492 21732 14544
rect 21784 14492 21790 14544
rect 22112 14532 22140 14572
rect 22186 14560 22192 14612
rect 22244 14560 22250 14612
rect 22646 14560 22652 14612
rect 22704 14560 22710 14612
rect 23293 14603 23351 14609
rect 23293 14569 23305 14603
rect 23339 14600 23351 14603
rect 24946 14600 24952 14612
rect 23339 14572 24952 14600
rect 23339 14569 23351 14572
rect 23293 14563 23351 14569
rect 24946 14560 24952 14572
rect 25004 14560 25010 14612
rect 25498 14560 25504 14612
rect 25556 14600 25562 14612
rect 25593 14603 25651 14609
rect 25593 14600 25605 14603
rect 25556 14572 25605 14600
rect 25556 14560 25562 14572
rect 25593 14569 25605 14572
rect 25639 14569 25651 14603
rect 25593 14563 25651 14569
rect 27798 14560 27804 14612
rect 27856 14600 27862 14612
rect 27893 14603 27951 14609
rect 27893 14600 27905 14603
rect 27856 14572 27905 14600
rect 27856 14560 27862 14572
rect 27893 14569 27905 14572
rect 27939 14569 27951 14603
rect 27893 14563 27951 14569
rect 28534 14560 28540 14612
rect 28592 14560 28598 14612
rect 28994 14600 29000 14612
rect 28644 14572 29000 14600
rect 22830 14532 22836 14544
rect 22112 14504 22836 14532
rect 22830 14492 22836 14504
rect 22888 14492 22894 14544
rect 24026 14492 24032 14544
rect 24084 14532 24090 14544
rect 25225 14535 25283 14541
rect 25225 14532 25237 14535
rect 24084 14504 25237 14532
rect 24084 14492 24090 14504
rect 25225 14501 25237 14504
rect 25271 14532 25283 14535
rect 27246 14532 27252 14544
rect 25271 14504 27252 14532
rect 25271 14501 25283 14504
rect 25225 14495 25283 14501
rect 27246 14492 27252 14504
rect 27304 14492 27310 14544
rect 21744 14464 21772 14492
rect 23566 14464 23572 14476
rect 21744 14436 21956 14464
rect 21637 14399 21695 14405
rect 21637 14396 21649 14399
rect 21284 14368 21649 14396
rect 18966 14328 18972 14340
rect 15795 14300 16988 14328
rect 17144 14300 17448 14328
rect 18800 14300 18972 14328
rect 15795 14297 15807 14300
rect 15749 14291 15807 14297
rect 13446 14260 13452 14272
rect 13280 14232 13452 14260
rect 13446 14220 13452 14232
rect 13504 14260 13510 14272
rect 16758 14260 16764 14272
rect 13504 14232 16764 14260
rect 13504 14220 13510 14232
rect 16758 14220 16764 14232
rect 16816 14220 16822 14272
rect 16960 14269 16988 14300
rect 17420 14272 17448 14300
rect 18966 14288 18972 14300
rect 19024 14288 19030 14340
rect 19337 14331 19395 14337
rect 19337 14297 19349 14331
rect 19383 14328 19395 14331
rect 19981 14331 20039 14337
rect 19981 14328 19993 14331
rect 19383 14300 19993 14328
rect 19383 14297 19395 14300
rect 19337 14291 19395 14297
rect 19981 14297 19993 14300
rect 20027 14297 20039 14331
rect 19981 14291 20039 14297
rect 20346 14288 20352 14340
rect 20404 14328 20410 14340
rect 20732 14328 20760 14359
rect 20404 14300 20760 14328
rect 20977 14331 21035 14337
rect 20404 14288 20410 14300
rect 20548 14272 20576 14300
rect 20977 14297 20989 14331
rect 21023 14328 21035 14331
rect 21100 14328 21128 14368
rect 21637 14365 21649 14368
rect 21683 14365 21695 14399
rect 21637 14359 21695 14365
rect 21023 14300 21128 14328
rect 21177 14331 21235 14337
rect 21023 14297 21035 14300
rect 20977 14291 21035 14297
rect 21177 14297 21189 14331
rect 21223 14328 21235 14331
rect 21266 14328 21272 14340
rect 21223 14300 21272 14328
rect 21223 14297 21235 14300
rect 21177 14291 21235 14297
rect 21266 14288 21272 14300
rect 21324 14288 21330 14340
rect 21652 14328 21680 14359
rect 21726 14356 21732 14408
rect 21784 14356 21790 14408
rect 21928 14405 21956 14436
rect 23032 14436 23572 14464
rect 21913 14399 21971 14405
rect 21913 14365 21925 14399
rect 21959 14365 21971 14399
rect 21913 14359 21971 14365
rect 22005 14399 22063 14405
rect 22005 14365 22017 14399
rect 22051 14396 22063 14399
rect 22094 14396 22100 14408
rect 22051 14368 22100 14396
rect 22051 14365 22063 14368
rect 22005 14359 22063 14365
rect 22094 14356 22100 14368
rect 22152 14356 22158 14408
rect 22738 14356 22744 14408
rect 22796 14356 22802 14408
rect 23032 14405 23060 14436
rect 23566 14424 23572 14436
rect 23624 14464 23630 14476
rect 24302 14464 24308 14476
rect 23624 14436 24308 14464
rect 23624 14424 23630 14436
rect 24302 14424 24308 14436
rect 24360 14424 24366 14476
rect 24946 14424 24952 14476
rect 25004 14464 25010 14476
rect 25314 14464 25320 14476
rect 25004 14436 25320 14464
rect 25004 14424 25010 14436
rect 25314 14424 25320 14436
rect 25372 14424 25378 14476
rect 26053 14467 26111 14473
rect 26053 14433 26065 14467
rect 26099 14464 26111 14467
rect 26099 14436 27660 14464
rect 26099 14433 26111 14436
rect 26053 14427 26111 14433
rect 22833 14399 22891 14405
rect 22833 14365 22845 14399
rect 22879 14365 22891 14399
rect 22833 14359 22891 14365
rect 23017 14399 23075 14405
rect 23017 14365 23029 14399
rect 23063 14365 23075 14399
rect 23017 14359 23075 14365
rect 22281 14331 22339 14337
rect 22281 14328 22293 14331
rect 21652 14300 22293 14328
rect 22281 14297 22293 14300
rect 22327 14297 22339 14331
rect 22281 14291 22339 14297
rect 22462 14288 22468 14340
rect 22520 14328 22526 14340
rect 22848 14328 22876 14359
rect 23106 14356 23112 14408
rect 23164 14396 23170 14408
rect 24578 14396 24584 14408
rect 23164 14368 24584 14396
rect 23164 14356 23170 14368
rect 24578 14356 24584 14368
rect 24636 14356 24642 14408
rect 24670 14356 24676 14408
rect 24728 14396 24734 14408
rect 25038 14396 25044 14408
rect 24728 14368 25044 14396
rect 24728 14356 24734 14368
rect 25038 14356 25044 14368
rect 25096 14356 25102 14408
rect 25225 14399 25283 14405
rect 25225 14365 25237 14399
rect 25271 14365 25283 14399
rect 25225 14359 25283 14365
rect 25777 14399 25835 14405
rect 25777 14365 25789 14399
rect 25823 14396 25835 14399
rect 25866 14396 25872 14408
rect 25823 14368 25872 14396
rect 25823 14365 25835 14368
rect 25777 14359 25835 14365
rect 22520 14300 22876 14328
rect 25240 14328 25268 14359
rect 25866 14356 25872 14368
rect 25924 14356 25930 14408
rect 25958 14356 25964 14408
rect 26016 14356 26022 14408
rect 26421 14399 26479 14405
rect 26421 14365 26433 14399
rect 26467 14365 26479 14399
rect 26421 14359 26479 14365
rect 26605 14399 26663 14405
rect 26605 14365 26617 14399
rect 26651 14396 26663 14399
rect 27430 14396 27436 14408
rect 26651 14368 27436 14396
rect 26651 14365 26663 14368
rect 26605 14359 26663 14365
rect 26436 14328 26464 14359
rect 27430 14356 27436 14368
rect 27488 14356 27494 14408
rect 25240 14300 26648 14328
rect 22520 14288 22526 14300
rect 26620 14272 26648 14300
rect 16945 14263 17003 14269
rect 16945 14229 16957 14263
rect 16991 14229 17003 14263
rect 16945 14223 17003 14229
rect 17402 14220 17408 14272
rect 17460 14220 17466 14272
rect 17862 14220 17868 14272
rect 17920 14260 17926 14272
rect 18509 14263 18567 14269
rect 18509 14260 18521 14263
rect 17920 14232 18521 14260
rect 17920 14220 17926 14232
rect 18509 14229 18521 14232
rect 18555 14229 18567 14263
rect 18509 14223 18567 14229
rect 20530 14220 20536 14272
rect 20588 14220 20594 14272
rect 23750 14220 23756 14272
rect 23808 14260 23814 14272
rect 23934 14260 23940 14272
rect 23808 14232 23940 14260
rect 23808 14220 23814 14232
rect 23934 14220 23940 14232
rect 23992 14220 23998 14272
rect 26418 14220 26424 14272
rect 26476 14220 26482 14272
rect 26602 14220 26608 14272
rect 26660 14220 26666 14272
rect 27632 14260 27660 14436
rect 28074 14356 28080 14408
rect 28132 14356 28138 14408
rect 28169 14399 28227 14405
rect 28169 14365 28181 14399
rect 28215 14365 28227 14399
rect 28169 14359 28227 14365
rect 27706 14288 27712 14340
rect 27764 14328 27770 14340
rect 28184 14328 28212 14359
rect 28258 14356 28264 14408
rect 28316 14356 28322 14408
rect 28353 14399 28411 14405
rect 28353 14365 28365 14399
rect 28399 14396 28411 14399
rect 28644 14396 28672 14572
rect 28994 14560 29000 14572
rect 29052 14560 29058 14612
rect 35894 14560 35900 14612
rect 35952 14600 35958 14612
rect 36078 14600 36084 14612
rect 35952 14572 36084 14600
rect 35952 14560 35958 14572
rect 36078 14560 36084 14572
rect 36136 14600 36142 14612
rect 36446 14600 36452 14612
rect 36136 14572 36452 14600
rect 36136 14560 36142 14572
rect 36446 14560 36452 14572
rect 36504 14560 36510 14612
rect 36633 14603 36691 14609
rect 36633 14569 36645 14603
rect 36679 14600 36691 14603
rect 37458 14600 37464 14612
rect 36679 14572 37464 14600
rect 36679 14569 36691 14572
rect 36633 14563 36691 14569
rect 37458 14560 37464 14572
rect 37516 14560 37522 14612
rect 28902 14492 28908 14544
rect 28960 14492 28966 14544
rect 29638 14492 29644 14544
rect 29696 14532 29702 14544
rect 29696 14504 37044 14532
rect 29696 14492 29702 14504
rect 28813 14467 28871 14473
rect 28813 14433 28825 14467
rect 28859 14464 28871 14467
rect 30101 14467 30159 14473
rect 30101 14464 30113 14467
rect 28859 14436 30113 14464
rect 28859 14433 28871 14436
rect 28813 14427 28871 14433
rect 28920 14408 28948 14436
rect 30101 14433 30113 14436
rect 30147 14433 30159 14467
rect 31018 14464 31024 14476
rect 30101 14427 30159 14433
rect 30300 14436 31024 14464
rect 28399 14368 28672 14396
rect 28721 14399 28779 14405
rect 28399 14365 28411 14368
rect 28353 14359 28411 14365
rect 28721 14365 28733 14399
rect 28767 14365 28779 14399
rect 28721 14359 28779 14365
rect 27764 14300 28212 14328
rect 27764 14288 27770 14300
rect 28534 14288 28540 14340
rect 28592 14328 28598 14340
rect 28736 14328 28764 14359
rect 28902 14356 28908 14408
rect 28960 14356 28966 14408
rect 28994 14356 29000 14408
rect 29052 14356 29058 14408
rect 30300 14405 30328 14436
rect 31018 14424 31024 14436
rect 31076 14464 31082 14476
rect 33594 14464 33600 14476
rect 31076 14436 33600 14464
rect 31076 14424 31082 14436
rect 33594 14424 33600 14436
rect 33652 14424 33658 14476
rect 36280 14436 36860 14464
rect 30285 14399 30343 14405
rect 30285 14365 30297 14399
rect 30331 14365 30343 14399
rect 30285 14359 30343 14365
rect 30466 14356 30472 14408
rect 30524 14396 30530 14408
rect 30561 14399 30619 14405
rect 30561 14396 30573 14399
rect 30524 14368 30573 14396
rect 30524 14356 30530 14368
rect 30561 14365 30573 14368
rect 30607 14365 30619 14399
rect 30561 14359 30619 14365
rect 35894 14356 35900 14408
rect 35952 14396 35958 14408
rect 36280 14405 36308 14436
rect 36832 14408 36860 14436
rect 36081 14399 36139 14405
rect 36081 14396 36093 14399
rect 35952 14368 36093 14396
rect 35952 14356 35958 14368
rect 36081 14365 36093 14368
rect 36127 14365 36139 14399
rect 36081 14359 36139 14365
rect 36265 14399 36323 14405
rect 36265 14365 36277 14399
rect 36311 14365 36323 14399
rect 36265 14359 36323 14365
rect 36449 14399 36507 14405
rect 36449 14365 36461 14399
rect 36495 14365 36507 14399
rect 36449 14359 36507 14365
rect 28592 14300 28764 14328
rect 28592 14288 28598 14300
rect 32950 14288 32956 14340
rect 33008 14328 33014 14340
rect 36357 14331 36415 14337
rect 36357 14328 36369 14331
rect 33008 14300 36369 14328
rect 33008 14288 33014 14300
rect 36357 14297 36369 14300
rect 36403 14297 36415 14331
rect 36357 14291 36415 14297
rect 36464 14328 36492 14359
rect 36630 14356 36636 14408
rect 36688 14396 36694 14408
rect 36725 14399 36783 14405
rect 36725 14396 36737 14399
rect 36688 14368 36737 14396
rect 36688 14356 36694 14368
rect 36725 14365 36737 14368
rect 36771 14365 36783 14399
rect 36725 14359 36783 14365
rect 36814 14356 36820 14408
rect 36872 14396 36878 14408
rect 37016 14405 37044 14504
rect 36909 14399 36967 14405
rect 36909 14396 36921 14399
rect 36872 14368 36921 14396
rect 36872 14356 36878 14368
rect 36909 14365 36921 14368
rect 36955 14365 36967 14399
rect 36909 14359 36967 14365
rect 37001 14399 37059 14405
rect 37001 14365 37013 14399
rect 37047 14365 37059 14399
rect 37001 14359 37059 14365
rect 37093 14399 37151 14405
rect 37093 14365 37105 14399
rect 37139 14365 37151 14399
rect 37093 14359 37151 14365
rect 37108 14328 37136 14359
rect 36464 14300 37136 14328
rect 30374 14260 30380 14272
rect 27632 14232 30380 14260
rect 30374 14220 30380 14232
rect 30432 14220 30438 14272
rect 30469 14263 30527 14269
rect 30469 14229 30481 14263
rect 30515 14260 30527 14263
rect 30558 14260 30564 14272
rect 30515 14232 30564 14260
rect 30515 14229 30527 14232
rect 30469 14223 30527 14229
rect 30558 14220 30564 14232
rect 30616 14220 30622 14272
rect 35342 14220 35348 14272
rect 35400 14260 35406 14272
rect 36464 14260 36492 14300
rect 35400 14232 36492 14260
rect 35400 14220 35406 14232
rect 37274 14220 37280 14272
rect 37332 14220 37338 14272
rect 1104 14170 40572 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 40572 14170
rect 1104 14096 40572 14118
rect 4157 14059 4215 14065
rect 4157 14025 4169 14059
rect 4203 14056 4215 14059
rect 4246 14056 4252 14068
rect 4203 14028 4252 14056
rect 4203 14025 4215 14028
rect 4157 14019 4215 14025
rect 4246 14016 4252 14028
rect 4304 14016 4310 14068
rect 5994 14016 6000 14068
rect 6052 14056 6058 14068
rect 7558 14056 7564 14068
rect 6052 14028 7564 14056
rect 6052 14016 6058 14028
rect 7558 14016 7564 14028
rect 7616 14016 7622 14068
rect 10134 14056 10140 14068
rect 9508 14028 10140 14056
rect 5902 13988 5908 14000
rect 4632 13960 5908 13988
rect 4154 13880 4160 13932
rect 4212 13920 4218 13932
rect 4341 13923 4399 13929
rect 4341 13920 4353 13923
rect 4212 13892 4353 13920
rect 4212 13880 4218 13892
rect 4341 13889 4353 13892
rect 4387 13889 4399 13923
rect 4341 13883 4399 13889
rect 4433 13923 4491 13929
rect 4433 13889 4445 13923
rect 4479 13920 4491 13923
rect 4522 13920 4528 13932
rect 4479 13892 4528 13920
rect 4479 13889 4491 13892
rect 4433 13883 4491 13889
rect 4522 13880 4528 13892
rect 4580 13880 4586 13932
rect 4632 13929 4660 13960
rect 5902 13948 5908 13960
rect 5960 13948 5966 14000
rect 7098 13948 7104 14000
rect 7156 13988 7162 14000
rect 8662 13988 8668 14000
rect 7156 13960 8668 13988
rect 7156 13948 7162 13960
rect 8662 13948 8668 13960
rect 8720 13948 8726 14000
rect 4617 13923 4675 13929
rect 4617 13889 4629 13923
rect 4663 13889 4675 13923
rect 4617 13883 4675 13889
rect 4706 13880 4712 13932
rect 4764 13880 4770 13932
rect 9401 13923 9459 13929
rect 9401 13889 9413 13923
rect 9447 13920 9459 13923
rect 9508 13920 9536 14028
rect 10134 14016 10140 14028
rect 10192 14016 10198 14068
rect 13170 14056 13176 14068
rect 10612 14028 13176 14056
rect 9585 13991 9643 13997
rect 9585 13957 9597 13991
rect 9631 13988 9643 13991
rect 9950 13988 9956 14000
rect 9631 13960 9956 13988
rect 9631 13957 9643 13960
rect 9585 13951 9643 13957
rect 9950 13948 9956 13960
rect 10008 13948 10014 14000
rect 9447 13892 9536 13920
rect 9677 13923 9735 13929
rect 9447 13889 9459 13892
rect 9401 13883 9459 13889
rect 9677 13889 9689 13923
rect 9723 13920 9735 13923
rect 9766 13920 9772 13932
rect 9723 13892 9772 13920
rect 9723 13889 9735 13892
rect 9677 13883 9735 13889
rect 9766 13880 9772 13892
rect 9824 13920 9830 13932
rect 10410 13920 10416 13932
rect 9824 13892 10416 13920
rect 9824 13880 9830 13892
rect 10410 13880 10416 13892
rect 10468 13880 10474 13932
rect 10502 13880 10508 13932
rect 10560 13880 10566 13932
rect 10612 13929 10640 14028
rect 13170 14016 13176 14028
rect 13228 14016 13234 14068
rect 16025 14059 16083 14065
rect 16025 14025 16037 14059
rect 16071 14056 16083 14059
rect 16666 14056 16672 14068
rect 16071 14028 16672 14056
rect 16071 14025 16083 14028
rect 16025 14019 16083 14025
rect 16666 14016 16672 14028
rect 16724 14016 16730 14068
rect 16758 14016 16764 14068
rect 16816 14056 16822 14068
rect 19705 14059 19763 14065
rect 19705 14056 19717 14059
rect 16816 14028 19717 14056
rect 16816 14016 16822 14028
rect 19705 14025 19717 14028
rect 19751 14025 19763 14059
rect 19705 14019 19763 14025
rect 20070 14016 20076 14068
rect 20128 14056 20134 14068
rect 21726 14056 21732 14068
rect 20128 14028 21732 14056
rect 20128 14016 20134 14028
rect 21726 14016 21732 14028
rect 21784 14016 21790 14068
rect 22278 14056 22284 14068
rect 21836 14028 22284 14056
rect 12526 13988 12532 14000
rect 10888 13960 12532 13988
rect 10888 13929 10916 13960
rect 12526 13948 12532 13960
rect 12584 13948 12590 14000
rect 13633 13991 13691 13997
rect 13633 13988 13645 13991
rect 12820 13960 13645 13988
rect 12820 13932 12848 13960
rect 13633 13957 13645 13960
rect 13679 13957 13691 13991
rect 13633 13951 13691 13957
rect 16206 13948 16212 14000
rect 16264 13988 16270 14000
rect 17218 13988 17224 14000
rect 16264 13960 17224 13988
rect 16264 13948 16270 13960
rect 17218 13948 17224 13960
rect 17276 13988 17282 14000
rect 17862 13988 17868 14000
rect 17276 13960 17868 13988
rect 17276 13948 17282 13960
rect 17862 13948 17868 13960
rect 17920 13948 17926 14000
rect 18966 13948 18972 14000
rect 19024 13988 19030 14000
rect 19024 13960 20024 13988
rect 19024 13948 19030 13960
rect 10597 13923 10655 13929
rect 10597 13889 10609 13923
rect 10643 13889 10655 13923
rect 10597 13883 10655 13889
rect 10689 13923 10747 13929
rect 10689 13889 10701 13923
rect 10735 13889 10747 13923
rect 10689 13883 10747 13889
rect 10867 13923 10925 13929
rect 10867 13889 10879 13923
rect 10913 13889 10925 13923
rect 10867 13883 10925 13889
rect 7282 13812 7288 13864
rect 7340 13852 7346 13864
rect 10612 13852 10640 13883
rect 7340 13824 10640 13852
rect 10704 13852 10732 13883
rect 11054 13880 11060 13932
rect 11112 13880 11118 13932
rect 11241 13923 11299 13929
rect 11241 13889 11253 13923
rect 11287 13920 11299 13923
rect 11514 13920 11520 13932
rect 11287 13892 11520 13920
rect 11287 13889 11299 13892
rect 11241 13883 11299 13889
rect 11514 13880 11520 13892
rect 11572 13880 11578 13932
rect 11793 13923 11851 13929
rect 11793 13889 11805 13923
rect 11839 13889 11851 13923
rect 11793 13883 11851 13889
rect 11977 13923 12035 13929
rect 11977 13889 11989 13923
rect 12023 13920 12035 13923
rect 12342 13920 12348 13932
rect 12023 13892 12348 13920
rect 12023 13889 12035 13892
rect 11977 13883 12035 13889
rect 10704 13824 10916 13852
rect 7340 13812 7346 13824
rect 4338 13744 4344 13796
rect 4396 13784 4402 13796
rect 5166 13784 5172 13796
rect 4396 13756 5172 13784
rect 4396 13744 4402 13756
rect 5166 13744 5172 13756
rect 5224 13784 5230 13796
rect 5718 13784 5724 13796
rect 5224 13756 5724 13784
rect 5224 13744 5230 13756
rect 5718 13744 5724 13756
rect 5776 13784 5782 13796
rect 9858 13784 9864 13796
rect 5776 13756 9864 13784
rect 5776 13744 5782 13756
rect 9858 13744 9864 13756
rect 9916 13744 9922 13796
rect 10888 13784 10916 13824
rect 10962 13812 10968 13864
rect 11020 13852 11026 13864
rect 11149 13855 11207 13861
rect 11149 13852 11161 13855
rect 11020 13824 11161 13852
rect 11020 13812 11026 13824
rect 11149 13821 11161 13824
rect 11195 13821 11207 13855
rect 11808 13852 11836 13883
rect 12342 13880 12348 13892
rect 12400 13880 12406 13932
rect 12618 13880 12624 13932
rect 12676 13880 12682 13932
rect 12802 13880 12808 13932
rect 12860 13880 12866 13932
rect 12897 13923 12955 13929
rect 12897 13889 12909 13923
rect 12943 13920 12955 13923
rect 12986 13920 12992 13932
rect 12943 13892 12992 13920
rect 12943 13889 12955 13892
rect 12897 13883 12955 13889
rect 12986 13880 12992 13892
rect 13044 13880 13050 13932
rect 13173 13923 13231 13929
rect 13173 13889 13185 13923
rect 13219 13920 13231 13923
rect 13262 13920 13268 13932
rect 13219 13892 13268 13920
rect 13219 13889 13231 13892
rect 13173 13883 13231 13889
rect 13262 13880 13268 13892
rect 13320 13880 13326 13932
rect 13354 13880 13360 13932
rect 13412 13920 13418 13932
rect 13909 13923 13967 13929
rect 13412 13892 13860 13920
rect 13412 13880 13418 13892
rect 12434 13852 12440 13864
rect 11808 13824 12440 13852
rect 11149 13815 11207 13821
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 12636 13852 12664 13880
rect 13630 13852 13636 13864
rect 12636 13824 13216 13852
rect 11054 13784 11060 13796
rect 10888 13756 11060 13784
rect 11054 13744 11060 13756
rect 11112 13744 11118 13796
rect 12452 13784 12480 13812
rect 12710 13784 12716 13796
rect 12452 13756 12716 13784
rect 12710 13744 12716 13756
rect 12768 13744 12774 13796
rect 13188 13784 13216 13824
rect 13372 13824 13636 13852
rect 13372 13784 13400 13824
rect 13630 13812 13636 13824
rect 13688 13852 13694 13864
rect 13725 13855 13783 13861
rect 13725 13852 13737 13855
rect 13688 13824 13737 13852
rect 13688 13812 13694 13824
rect 13725 13821 13737 13824
rect 13771 13821 13783 13855
rect 13725 13815 13783 13821
rect 13188 13756 13400 13784
rect 13832 13784 13860 13892
rect 13909 13889 13921 13923
rect 13955 13920 13967 13923
rect 14458 13920 14464 13932
rect 13955 13892 14464 13920
rect 13955 13889 13967 13892
rect 13909 13883 13967 13889
rect 14458 13880 14464 13892
rect 14516 13880 14522 13932
rect 16393 13923 16451 13929
rect 16393 13889 16405 13923
rect 16439 13889 16451 13923
rect 16393 13883 16451 13889
rect 13832 13756 14228 13784
rect 9214 13676 9220 13728
rect 9272 13676 9278 13728
rect 10226 13676 10232 13728
rect 10284 13676 10290 13728
rect 11790 13676 11796 13728
rect 11848 13716 11854 13728
rect 11977 13719 12035 13725
rect 11977 13716 11989 13719
rect 11848 13688 11989 13716
rect 11848 13676 11854 13688
rect 11977 13685 11989 13688
rect 12023 13685 12035 13719
rect 11977 13679 12035 13685
rect 12434 13676 12440 13728
rect 12492 13676 12498 13728
rect 12802 13676 12808 13728
rect 12860 13716 12866 13728
rect 12989 13719 13047 13725
rect 12989 13716 13001 13719
rect 12860 13688 13001 13716
rect 12860 13676 12866 13688
rect 12989 13685 13001 13688
rect 13035 13685 13047 13719
rect 12989 13679 13047 13685
rect 13078 13676 13084 13728
rect 13136 13716 13142 13728
rect 13173 13719 13231 13725
rect 13173 13716 13185 13719
rect 13136 13688 13185 13716
rect 13136 13676 13142 13688
rect 13173 13685 13185 13688
rect 13219 13685 13231 13719
rect 13173 13679 13231 13685
rect 14090 13676 14096 13728
rect 14148 13676 14154 13728
rect 14200 13716 14228 13756
rect 15194 13744 15200 13796
rect 15252 13784 15258 13796
rect 15562 13784 15568 13796
rect 15252 13756 15568 13784
rect 15252 13744 15258 13756
rect 15562 13744 15568 13756
rect 15620 13784 15626 13796
rect 16408 13784 16436 13883
rect 19242 13880 19248 13932
rect 19300 13920 19306 13932
rect 19613 13923 19671 13929
rect 19613 13920 19625 13923
rect 19300 13892 19625 13920
rect 19300 13880 19306 13892
rect 19613 13889 19625 13892
rect 19659 13889 19671 13923
rect 19613 13883 19671 13889
rect 19797 13923 19855 13929
rect 19797 13889 19809 13923
rect 19843 13920 19855 13923
rect 19886 13920 19892 13932
rect 19843 13892 19892 13920
rect 19843 13889 19855 13892
rect 19797 13883 19855 13889
rect 19886 13880 19892 13892
rect 19944 13880 19950 13932
rect 19996 13920 20024 13960
rect 20346 13948 20352 14000
rect 20404 13988 20410 14000
rect 21836 13988 21864 14028
rect 22278 14016 22284 14028
rect 22336 14016 22342 14068
rect 23661 14059 23719 14065
rect 23661 14025 23673 14059
rect 23707 14056 23719 14059
rect 23750 14056 23756 14068
rect 23707 14028 23756 14056
rect 23707 14025 23719 14028
rect 23661 14019 23719 14025
rect 23750 14016 23756 14028
rect 23808 14016 23814 14068
rect 23845 14059 23903 14065
rect 23845 14025 23857 14059
rect 23891 14056 23903 14059
rect 23934 14056 23940 14068
rect 23891 14028 23940 14056
rect 23891 14025 23903 14028
rect 23845 14019 23903 14025
rect 23934 14016 23940 14028
rect 23992 14016 23998 14068
rect 24029 14059 24087 14065
rect 24029 14025 24041 14059
rect 24075 14056 24087 14059
rect 24210 14056 24216 14068
rect 24075 14028 24216 14056
rect 24075 14025 24087 14028
rect 24029 14019 24087 14025
rect 24210 14016 24216 14028
rect 24268 14016 24274 14068
rect 24302 14016 24308 14068
rect 24360 14016 24366 14068
rect 24486 14065 24492 14068
rect 24473 14059 24492 14065
rect 24473 14025 24485 14059
rect 24473 14019 24492 14025
rect 24486 14016 24492 14019
rect 24544 14016 24550 14068
rect 25777 14059 25835 14065
rect 25777 14025 25789 14059
rect 25823 14056 25835 14059
rect 25958 14056 25964 14068
rect 25823 14028 25964 14056
rect 25823 14025 25835 14028
rect 25777 14019 25835 14025
rect 25958 14016 25964 14028
rect 26016 14016 26022 14068
rect 26160 14028 26464 14056
rect 20404 13960 21864 13988
rect 20404 13948 20410 13960
rect 22002 13948 22008 14000
rect 22060 13988 22066 14000
rect 24118 13988 24124 14000
rect 22060 13960 24124 13988
rect 22060 13948 22066 13960
rect 24118 13948 24124 13960
rect 24176 13948 24182 14000
rect 24670 13948 24676 14000
rect 24728 13948 24734 14000
rect 20714 13920 20720 13932
rect 19996 13892 20720 13920
rect 20714 13880 20720 13892
rect 20772 13920 20778 13932
rect 23014 13920 23020 13932
rect 20772 13918 21864 13920
rect 22020 13918 23020 13920
rect 20772 13892 23020 13918
rect 20772 13880 20778 13892
rect 21836 13890 22048 13892
rect 23014 13880 23020 13892
rect 23072 13880 23078 13932
rect 23937 13923 23995 13929
rect 23937 13889 23949 13923
rect 23983 13889 23995 13923
rect 23937 13883 23995 13889
rect 24213 13923 24271 13929
rect 24213 13889 24225 13923
rect 24259 13920 24271 13923
rect 24688 13920 24716 13948
rect 24259 13892 24716 13920
rect 24259 13889 24271 13892
rect 24213 13883 24271 13889
rect 20162 13812 20168 13864
rect 20220 13852 20226 13864
rect 20220 13824 20852 13852
rect 20220 13812 20226 13824
rect 18598 13784 18604 13796
rect 15620 13756 18604 13784
rect 15620 13744 15626 13756
rect 18598 13744 18604 13756
rect 18656 13744 18662 13796
rect 19886 13744 19892 13796
rect 19944 13784 19950 13796
rect 20254 13784 20260 13796
rect 19944 13756 20260 13784
rect 19944 13744 19950 13756
rect 20254 13744 20260 13756
rect 20312 13744 20318 13796
rect 20824 13784 20852 13824
rect 22094 13812 22100 13864
rect 22152 13852 22158 13864
rect 23106 13852 23112 13864
rect 22152 13824 23112 13852
rect 22152 13812 22158 13824
rect 23106 13812 23112 13824
rect 23164 13812 23170 13864
rect 23952 13852 23980 13883
rect 25038 13880 25044 13932
rect 25096 13920 25102 13932
rect 25685 13923 25743 13929
rect 25685 13920 25697 13923
rect 25096 13892 25697 13920
rect 25096 13880 25102 13892
rect 25685 13889 25697 13892
rect 25731 13889 25743 13923
rect 25685 13883 25743 13889
rect 25869 13923 25927 13929
rect 25869 13889 25881 13923
rect 25915 13920 25927 13923
rect 26160 13920 26188 14028
rect 26234 13948 26240 14000
rect 26292 13948 26298 14000
rect 26436 13988 26464 14028
rect 26694 14016 26700 14068
rect 26752 14056 26758 14068
rect 27062 14056 27068 14068
rect 26752 14028 27068 14056
rect 26752 14016 26758 14028
rect 27062 14016 27068 14028
rect 27120 14016 27126 14068
rect 27985 14059 28043 14065
rect 27985 14025 27997 14059
rect 28031 14056 28043 14059
rect 28258 14056 28264 14068
rect 28031 14028 28264 14056
rect 28031 14025 28043 14028
rect 27985 14019 28043 14025
rect 28258 14016 28264 14028
rect 28316 14016 28322 14068
rect 32950 14056 32956 14068
rect 28363 14028 32956 14056
rect 26436 13960 27016 13988
rect 25915 13892 26188 13920
rect 26252 13918 26280 13948
rect 26988 13929 27016 13960
rect 27246 13948 27252 14000
rect 27304 13988 27310 14000
rect 28363 13988 28391 14028
rect 32950 14016 32956 14028
rect 33008 14016 33014 14068
rect 33045 14059 33103 14065
rect 33045 14025 33057 14059
rect 33091 14025 33103 14059
rect 33045 14019 33103 14025
rect 27304 13960 28391 13988
rect 27304 13948 27310 13960
rect 28442 13948 28448 14000
rect 28500 13948 28506 14000
rect 28534 13948 28540 14000
rect 28592 13988 28598 14000
rect 28718 13988 28724 14000
rect 28592 13960 28724 13988
rect 28592 13948 28598 13960
rect 28718 13948 28724 13960
rect 28776 13948 28782 14000
rect 32030 13948 32036 14000
rect 32088 13988 32094 14000
rect 32214 13988 32220 14000
rect 32088 13960 32220 13988
rect 32088 13948 32094 13960
rect 32214 13948 32220 13960
rect 32272 13988 32278 14000
rect 33060 13988 33088 14019
rect 36998 14016 37004 14068
rect 37056 14056 37062 14068
rect 37093 14059 37151 14065
rect 37093 14056 37105 14059
rect 37056 14028 37105 14056
rect 37056 14016 37062 14028
rect 37093 14025 37105 14028
rect 37139 14025 37151 14059
rect 37093 14019 37151 14025
rect 38841 14059 38899 14065
rect 38841 14025 38853 14059
rect 38887 14056 38899 14059
rect 39206 14056 39212 14068
rect 38887 14028 39212 14056
rect 38887 14025 38899 14028
rect 38841 14019 38899 14025
rect 39206 14016 39212 14028
rect 39264 14016 39270 14068
rect 34698 13988 34704 14000
rect 32272 13960 32904 13988
rect 33060 13960 34704 13988
rect 32272 13948 32278 13960
rect 26421 13923 26479 13929
rect 26421 13918 26433 13923
rect 25915 13889 25927 13892
rect 26252 13890 26433 13918
rect 25869 13883 25927 13889
rect 26421 13889 26433 13890
rect 26467 13889 26479 13923
rect 26421 13883 26479 13889
rect 26973 13923 27031 13929
rect 26973 13889 26985 13923
rect 27019 13889 27031 13923
rect 26973 13883 27031 13889
rect 27157 13923 27215 13929
rect 27157 13889 27169 13923
rect 27203 13920 27215 13923
rect 27430 13920 27436 13932
rect 27203 13892 27436 13920
rect 27203 13889 27215 13892
rect 27157 13883 27215 13889
rect 24118 13852 24124 13864
rect 23952 13824 24124 13852
rect 21266 13784 21272 13796
rect 20824 13756 21272 13784
rect 21266 13744 21272 13756
rect 21324 13744 21330 13796
rect 22830 13744 22836 13796
rect 22888 13784 22894 13796
rect 23952 13784 23980 13824
rect 24118 13812 24124 13824
rect 24176 13852 24182 13864
rect 24486 13852 24492 13864
rect 24176 13824 24492 13852
rect 24176 13812 24182 13824
rect 24486 13812 24492 13824
rect 24544 13812 24550 13864
rect 25700 13852 25728 13883
rect 26050 13852 26056 13864
rect 25700 13824 26056 13852
rect 26050 13812 26056 13824
rect 26108 13812 26114 13864
rect 26237 13855 26295 13861
rect 26237 13821 26249 13855
rect 26283 13821 26295 13855
rect 26237 13815 26295 13821
rect 26252 13784 26280 13815
rect 26510 13812 26516 13864
rect 26568 13812 26574 13864
rect 26605 13855 26663 13861
rect 26605 13821 26617 13855
rect 26651 13821 26663 13855
rect 26605 13815 26663 13821
rect 22888 13756 23980 13784
rect 24412 13756 26280 13784
rect 26620 13784 26648 13815
rect 26694 13812 26700 13864
rect 26752 13812 26758 13864
rect 26988 13852 27016 13883
rect 27430 13880 27436 13892
rect 27488 13880 27494 13932
rect 28074 13880 28080 13932
rect 28132 13920 28138 13932
rect 28169 13923 28227 13929
rect 28169 13920 28181 13923
rect 28132 13892 28181 13920
rect 28132 13880 28138 13892
rect 28169 13889 28181 13892
rect 28215 13889 28227 13923
rect 28810 13920 28816 13932
rect 28169 13883 28227 13889
rect 28276 13892 28816 13920
rect 27246 13852 27252 13864
rect 26988 13824 27252 13852
rect 27246 13812 27252 13824
rect 27304 13812 27310 13864
rect 27614 13812 27620 13864
rect 27672 13852 27678 13864
rect 28276 13852 28304 13892
rect 28810 13880 28816 13892
rect 28868 13920 28874 13932
rect 28905 13923 28963 13929
rect 28905 13920 28917 13923
rect 28868 13892 28917 13920
rect 28868 13880 28874 13892
rect 28905 13889 28917 13892
rect 28951 13920 28963 13923
rect 29546 13920 29552 13932
rect 28951 13892 29552 13920
rect 28951 13889 28963 13892
rect 28905 13883 28963 13889
rect 29546 13880 29552 13892
rect 29604 13880 29610 13932
rect 30558 13880 30564 13932
rect 30616 13880 30622 13932
rect 30653 13923 30711 13929
rect 30653 13889 30665 13923
rect 30699 13920 30711 13923
rect 31386 13920 31392 13932
rect 30699 13892 31392 13920
rect 30699 13889 30711 13892
rect 30653 13883 30711 13889
rect 31386 13880 31392 13892
rect 31444 13920 31450 13932
rect 31570 13920 31576 13932
rect 31444 13892 31576 13920
rect 31444 13880 31450 13892
rect 31570 13880 31576 13892
rect 31628 13880 31634 13932
rect 32585 13923 32643 13929
rect 32585 13889 32597 13923
rect 32631 13889 32643 13923
rect 32585 13883 32643 13889
rect 27672 13824 28304 13852
rect 28353 13855 28411 13861
rect 27672 13812 27678 13824
rect 28353 13821 28365 13855
rect 28399 13852 28411 13855
rect 30282 13852 30288 13864
rect 28399 13824 30288 13852
rect 28399 13821 28411 13824
rect 28353 13815 28411 13821
rect 30282 13812 30288 13824
rect 30340 13812 30346 13864
rect 30742 13812 30748 13864
rect 30800 13852 30806 13864
rect 30837 13855 30895 13861
rect 30837 13852 30849 13855
rect 30800 13824 30849 13852
rect 30800 13812 30806 13824
rect 30837 13821 30849 13824
rect 30883 13821 30895 13855
rect 32600 13852 32628 13883
rect 32766 13880 32772 13932
rect 32824 13880 32830 13932
rect 32876 13929 32904 13960
rect 34698 13948 34704 13960
rect 34756 13948 34762 14000
rect 36078 13948 36084 14000
rect 36136 13988 36142 14000
rect 36814 13988 36820 14000
rect 36136 13960 36820 13988
rect 36136 13948 36142 13960
rect 36814 13948 36820 13960
rect 36872 13948 36878 14000
rect 37182 13948 37188 14000
rect 37240 13988 37246 14000
rect 37277 13991 37335 13997
rect 37277 13988 37289 13991
rect 37240 13960 37289 13988
rect 37240 13948 37246 13960
rect 37277 13957 37289 13960
rect 37323 13957 37335 13991
rect 39390 13988 39396 14000
rect 37277 13951 37335 13957
rect 37384 13960 39396 13988
rect 32861 13923 32919 13929
rect 32861 13889 32873 13923
rect 32907 13889 32919 13923
rect 32861 13883 32919 13889
rect 36722 13880 36728 13932
rect 36780 13880 36786 13932
rect 36906 13880 36912 13932
rect 36964 13880 36970 13932
rect 32950 13852 32956 13864
rect 32600 13824 32956 13852
rect 30837 13815 30895 13821
rect 27154 13784 27160 13796
rect 26620 13756 27160 13784
rect 22888 13744 22894 13756
rect 18230 13716 18236 13728
rect 14200 13688 18236 13716
rect 18230 13676 18236 13688
rect 18288 13676 18294 13728
rect 19518 13676 19524 13728
rect 19576 13716 19582 13728
rect 22848 13716 22876 13744
rect 19576 13688 22876 13716
rect 19576 13676 19582 13688
rect 23934 13676 23940 13728
rect 23992 13716 23998 13728
rect 24412 13716 24440 13756
rect 23992 13688 24440 13716
rect 23992 13676 23998 13688
rect 24486 13676 24492 13728
rect 24544 13676 24550 13728
rect 26252 13716 26280 13756
rect 27154 13744 27160 13756
rect 27212 13744 27218 13796
rect 27798 13744 27804 13796
rect 27856 13784 27862 13796
rect 28721 13787 28779 13793
rect 27856 13756 28212 13784
rect 27856 13744 27862 13756
rect 28074 13716 28080 13728
rect 26252 13688 28080 13716
rect 28074 13676 28080 13688
rect 28132 13676 28138 13728
rect 28184 13725 28212 13756
rect 28721 13753 28733 13787
rect 28767 13784 28779 13787
rect 28994 13784 29000 13796
rect 28767 13756 29000 13784
rect 28767 13753 28779 13756
rect 28721 13747 28779 13753
rect 28994 13744 29000 13756
rect 29052 13744 29058 13796
rect 30852 13784 30880 13815
rect 32950 13812 32956 13824
rect 33008 13852 33014 13864
rect 33008 13824 33364 13852
rect 33008 13812 33014 13824
rect 33226 13784 33232 13796
rect 30852 13756 33232 13784
rect 33226 13744 33232 13756
rect 33284 13744 33290 13796
rect 33336 13784 33364 13824
rect 33594 13812 33600 13864
rect 33652 13852 33658 13864
rect 37384 13852 37412 13960
rect 39390 13948 39396 13960
rect 39448 13948 39454 14000
rect 37458 13880 37464 13932
rect 37516 13880 37522 13932
rect 37550 13880 37556 13932
rect 37608 13880 37614 13932
rect 38378 13880 38384 13932
rect 38436 13880 38442 13932
rect 38657 13923 38715 13929
rect 38657 13889 38669 13923
rect 38703 13920 38715 13923
rect 39758 13920 39764 13932
rect 38703 13892 39764 13920
rect 38703 13889 38715 13892
rect 38657 13883 38715 13889
rect 33652 13824 37412 13852
rect 33652 13812 33658 13824
rect 37642 13812 37648 13864
rect 37700 13852 37706 13864
rect 38473 13855 38531 13861
rect 38473 13852 38485 13855
rect 37700 13824 38485 13852
rect 37700 13812 37706 13824
rect 38473 13821 38485 13824
rect 38519 13821 38531 13855
rect 38473 13815 38531 13821
rect 36814 13784 36820 13796
rect 33336 13756 36820 13784
rect 36814 13744 36820 13756
rect 36872 13744 36878 13796
rect 37737 13787 37795 13793
rect 37737 13784 37749 13787
rect 36924 13756 37749 13784
rect 28169 13719 28227 13725
rect 28169 13685 28181 13719
rect 28215 13685 28227 13719
rect 28169 13679 28227 13685
rect 29178 13676 29184 13728
rect 29236 13716 29242 13728
rect 30742 13716 30748 13728
rect 29236 13688 30748 13716
rect 29236 13676 29242 13688
rect 30742 13676 30748 13688
rect 30800 13676 30806 13728
rect 32122 13676 32128 13728
rect 32180 13716 32186 13728
rect 32582 13716 32588 13728
rect 32180 13688 32588 13716
rect 32180 13676 32186 13688
rect 32582 13676 32588 13688
rect 32640 13676 32646 13728
rect 36924 13725 36952 13756
rect 37737 13753 37749 13756
rect 37783 13753 37795 13787
rect 37737 13747 37795 13753
rect 38102 13744 38108 13796
rect 38160 13784 38166 13796
rect 38672 13784 38700 13883
rect 39758 13880 39764 13892
rect 39816 13880 39822 13932
rect 38160 13756 38700 13784
rect 38160 13744 38166 13756
rect 38838 13744 38844 13796
rect 38896 13784 38902 13796
rect 39482 13784 39488 13796
rect 38896 13756 39488 13784
rect 38896 13744 38902 13756
rect 39482 13744 39488 13756
rect 39540 13744 39546 13796
rect 36909 13719 36967 13725
rect 36909 13685 36921 13719
rect 36955 13685 36967 13719
rect 36909 13679 36967 13685
rect 37274 13676 37280 13728
rect 37332 13676 37338 13728
rect 38562 13676 38568 13728
rect 38620 13676 38626 13728
rect 1104 13626 40572 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 40572 13626
rect 1104 13552 40572 13574
rect 3513 13515 3571 13521
rect 3513 13481 3525 13515
rect 3559 13512 3571 13515
rect 4062 13512 4068 13524
rect 3559 13484 4068 13512
rect 3559 13481 3571 13484
rect 3513 13475 3571 13481
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 4341 13515 4399 13521
rect 4341 13481 4353 13515
rect 4387 13512 4399 13515
rect 4614 13512 4620 13524
rect 4387 13484 4620 13512
rect 4387 13481 4399 13484
rect 4341 13475 4399 13481
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 5350 13512 5356 13524
rect 4724 13484 5356 13512
rect 4154 13404 4160 13456
rect 4212 13444 4218 13456
rect 4724 13444 4752 13484
rect 5350 13472 5356 13484
rect 5408 13472 5414 13524
rect 5902 13472 5908 13524
rect 5960 13512 5966 13524
rect 6733 13515 6791 13521
rect 6733 13512 6745 13515
rect 5960 13484 6745 13512
rect 5960 13472 5966 13484
rect 6733 13481 6745 13484
rect 6779 13481 6791 13515
rect 9214 13512 9220 13524
rect 6733 13475 6791 13481
rect 7208 13484 9220 13512
rect 4212 13416 4752 13444
rect 4212 13404 4218 13416
rect 5920 13376 5948 13472
rect 7208 13376 7236 13484
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 15933 13515 15991 13521
rect 15933 13481 15945 13515
rect 15979 13512 15991 13515
rect 16022 13512 16028 13524
rect 15979 13484 16028 13512
rect 15979 13481 15991 13484
rect 15933 13475 15991 13481
rect 16022 13472 16028 13484
rect 16080 13472 16086 13524
rect 16301 13515 16359 13521
rect 16301 13481 16313 13515
rect 16347 13512 16359 13515
rect 16666 13512 16672 13524
rect 16347 13484 16672 13512
rect 16347 13481 16359 13484
rect 16301 13475 16359 13481
rect 16666 13472 16672 13484
rect 16724 13472 16730 13524
rect 16850 13472 16856 13524
rect 16908 13472 16914 13524
rect 17034 13472 17040 13524
rect 17092 13472 17098 13524
rect 17218 13472 17224 13524
rect 17276 13472 17282 13524
rect 17954 13472 17960 13524
rect 18012 13472 18018 13524
rect 19889 13515 19947 13521
rect 19889 13512 19901 13515
rect 18064 13484 19901 13512
rect 7653 13447 7711 13453
rect 7653 13413 7665 13447
rect 7699 13444 7711 13447
rect 8110 13444 8116 13456
rect 7699 13416 8116 13444
rect 7699 13413 7711 13416
rect 7653 13407 7711 13413
rect 8110 13404 8116 13416
rect 8168 13404 8174 13456
rect 9858 13444 9864 13456
rect 9232 13416 9864 13444
rect 3436 13348 4660 13376
rect 3436 13317 3464 13348
rect 4632 13320 4660 13348
rect 5000 13348 5948 13376
rect 7116 13348 7236 13376
rect 7285 13379 7343 13385
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13277 3479 13311
rect 3421 13271 3479 13277
rect 3605 13311 3663 13317
rect 3605 13277 3617 13311
rect 3651 13308 3663 13311
rect 3970 13308 3976 13320
rect 3651 13280 3976 13308
rect 3651 13277 3663 13280
rect 3605 13271 3663 13277
rect 3970 13268 3976 13280
rect 4028 13308 4034 13320
rect 4525 13311 4583 13317
rect 4525 13308 4537 13311
rect 4028 13280 4537 13308
rect 4028 13268 4034 13280
rect 4525 13277 4537 13280
rect 4571 13277 4583 13311
rect 4525 13271 4583 13277
rect 3786 13200 3792 13252
rect 3844 13200 3850 13252
rect 4154 13200 4160 13252
rect 4212 13200 4218 13252
rect 4540 13240 4568 13271
rect 4614 13268 4620 13320
rect 4672 13308 4678 13320
rect 4709 13311 4767 13317
rect 4709 13308 4721 13311
rect 4672 13280 4721 13308
rect 4672 13268 4678 13280
rect 4709 13277 4721 13280
rect 4755 13277 4767 13311
rect 4709 13271 4767 13277
rect 4798 13268 4804 13320
rect 4856 13268 4862 13320
rect 5000 13317 5028 13348
rect 7116 13320 7144 13348
rect 7285 13345 7297 13379
rect 7331 13376 7343 13379
rect 7466 13376 7472 13388
rect 7331 13348 7472 13376
rect 7331 13345 7343 13348
rect 7285 13339 7343 13345
rect 7466 13336 7472 13348
rect 7524 13336 7530 13388
rect 8202 13376 8208 13388
rect 7852 13348 8208 13376
rect 4985 13311 5043 13317
rect 4985 13277 4997 13311
rect 5031 13277 5043 13311
rect 4985 13271 5043 13277
rect 5166 13268 5172 13320
rect 5224 13268 5230 13320
rect 5261 13311 5319 13317
rect 5261 13277 5273 13311
rect 5307 13308 5319 13311
rect 5810 13308 5816 13320
rect 5307 13280 5816 13308
rect 5307 13277 5319 13280
rect 5261 13271 5319 13277
rect 5276 13240 5304 13271
rect 5810 13268 5816 13280
rect 5868 13268 5874 13320
rect 6638 13268 6644 13320
rect 6696 13308 6702 13320
rect 6917 13311 6975 13317
rect 6917 13308 6929 13311
rect 6696 13280 6929 13308
rect 6696 13268 6702 13280
rect 6917 13277 6929 13280
rect 6963 13308 6975 13311
rect 6963 13280 7052 13308
rect 6963 13277 6975 13280
rect 6917 13271 6975 13277
rect 4540 13212 5304 13240
rect 7024 13240 7052 13280
rect 7098 13268 7104 13320
rect 7156 13268 7162 13320
rect 7193 13311 7251 13317
rect 7193 13277 7205 13311
rect 7239 13308 7251 13311
rect 7742 13308 7748 13320
rect 7239 13280 7748 13308
rect 7239 13277 7251 13280
rect 7193 13271 7251 13277
rect 7742 13268 7748 13280
rect 7800 13268 7806 13320
rect 7852 13317 7880 13348
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 9232 13385 9260 13416
rect 9858 13404 9864 13416
rect 9916 13404 9922 13456
rect 11054 13404 11060 13456
rect 11112 13444 11118 13456
rect 16868 13444 16896 13472
rect 11112 13416 12296 13444
rect 11112 13404 11118 13416
rect 12268 13388 12296 13416
rect 16224 13416 16896 13444
rect 17589 13447 17647 13453
rect 9217 13379 9275 13385
rect 9217 13345 9229 13379
rect 9263 13345 9275 13379
rect 9217 13339 9275 13345
rect 9766 13336 9772 13388
rect 9824 13336 9830 13388
rect 11241 13379 11299 13385
rect 11241 13345 11253 13379
rect 11287 13376 11299 13379
rect 11514 13376 11520 13388
rect 11287 13348 11520 13376
rect 11287 13345 11299 13348
rect 11241 13339 11299 13345
rect 11514 13336 11520 13348
rect 11572 13336 11578 13388
rect 12250 13336 12256 13388
rect 12308 13376 12314 13388
rect 12308 13348 13032 13376
rect 12308 13336 12314 13348
rect 7837 13311 7895 13317
rect 7837 13277 7849 13311
rect 7883 13277 7895 13311
rect 7837 13271 7895 13277
rect 7930 13311 7988 13317
rect 7930 13277 7942 13311
rect 7976 13277 7988 13311
rect 7930 13271 7988 13277
rect 7466 13240 7472 13252
rect 7024 13212 7472 13240
rect 7466 13200 7472 13212
rect 7524 13240 7530 13252
rect 7945 13240 7973 13271
rect 8018 13268 8024 13320
rect 8076 13308 8082 13320
rect 8113 13311 8171 13317
rect 8113 13308 8125 13311
rect 8076 13280 8125 13308
rect 8076 13268 8082 13280
rect 8113 13277 8125 13280
rect 8159 13277 8171 13311
rect 8113 13271 8171 13277
rect 8343 13311 8401 13317
rect 8343 13277 8355 13311
rect 8389 13308 8401 13311
rect 8754 13308 8760 13320
rect 8389 13280 8760 13308
rect 8389 13277 8401 13280
rect 8343 13271 8401 13277
rect 8754 13268 8760 13280
rect 8812 13268 8818 13320
rect 9950 13268 9956 13320
rect 10008 13268 10014 13320
rect 11149 13311 11207 13317
rect 11149 13277 11161 13311
rect 11195 13308 11207 13311
rect 11195 13280 11744 13308
rect 11195 13277 11207 13280
rect 11149 13271 11207 13277
rect 7524 13212 7973 13240
rect 7524 13200 7530 13212
rect 8202 13200 8208 13252
rect 8260 13200 8266 13252
rect 9968 13240 9996 13268
rect 11330 13240 11336 13252
rect 9968 13212 11336 13240
rect 11330 13200 11336 13212
rect 11388 13200 11394 13252
rect 11514 13200 11520 13252
rect 11572 13200 11578 13252
rect 4798 13132 4804 13184
rect 4856 13172 4862 13184
rect 4893 13175 4951 13181
rect 4893 13172 4905 13175
rect 4856 13144 4905 13172
rect 4856 13132 4862 13144
rect 4893 13141 4905 13144
rect 4939 13141 4951 13175
rect 4893 13135 4951 13141
rect 5445 13175 5503 13181
rect 5445 13141 5457 13175
rect 5491 13172 5503 13175
rect 5534 13172 5540 13184
rect 5491 13144 5540 13172
rect 5491 13141 5503 13144
rect 5445 13135 5503 13141
rect 5534 13132 5540 13144
rect 5592 13172 5598 13184
rect 6454 13172 6460 13184
rect 5592 13144 6460 13172
rect 5592 13132 5598 13144
rect 6454 13132 6460 13144
rect 6512 13132 6518 13184
rect 7742 13132 7748 13184
rect 7800 13132 7806 13184
rect 8294 13132 8300 13184
rect 8352 13172 8358 13184
rect 8481 13175 8539 13181
rect 8481 13172 8493 13175
rect 8352 13144 8493 13172
rect 8352 13132 8358 13144
rect 8481 13141 8493 13144
rect 8527 13141 8539 13175
rect 8481 13135 8539 13141
rect 8662 13132 8668 13184
rect 8720 13172 8726 13184
rect 10321 13175 10379 13181
rect 10321 13172 10333 13175
rect 8720 13144 10333 13172
rect 8720 13132 8726 13144
rect 10321 13141 10333 13144
rect 10367 13141 10379 13175
rect 11716 13172 11744 13280
rect 12342 13268 12348 13320
rect 12400 13268 12406 13320
rect 12529 13311 12587 13317
rect 12529 13277 12541 13311
rect 12575 13308 12587 13311
rect 12710 13308 12716 13320
rect 12575 13280 12716 13308
rect 12575 13277 12587 13280
rect 12529 13271 12587 13277
rect 12710 13268 12716 13280
rect 12768 13268 12774 13320
rect 12802 13268 12808 13320
rect 12860 13268 12866 13320
rect 13004 13317 13032 13348
rect 13170 13336 13176 13388
rect 13228 13336 13234 13388
rect 14093 13379 14151 13385
rect 14093 13345 14105 13379
rect 14139 13376 14151 13379
rect 14734 13376 14740 13388
rect 14139 13348 14740 13376
rect 14139 13345 14151 13348
rect 14093 13339 14151 13345
rect 14734 13336 14740 13348
rect 14792 13336 14798 13388
rect 16224 13385 16252 13416
rect 17589 13413 17601 13447
rect 17635 13413 17647 13447
rect 17589 13407 17647 13413
rect 16209 13379 16267 13385
rect 16209 13345 16221 13379
rect 16255 13345 16267 13379
rect 17604 13376 17632 13407
rect 18064 13376 18092 13484
rect 19889 13481 19901 13484
rect 19935 13481 19947 13515
rect 19889 13475 19947 13481
rect 21726 13472 21732 13524
rect 21784 13512 21790 13524
rect 22097 13515 22155 13521
rect 22097 13512 22109 13515
rect 21784 13484 22109 13512
rect 21784 13472 21790 13484
rect 22097 13481 22109 13484
rect 22143 13481 22155 13515
rect 22097 13475 22155 13481
rect 22204 13484 22692 13512
rect 20714 13376 20720 13388
rect 16209 13339 16267 13345
rect 16316 13348 17632 13376
rect 17696 13348 18092 13376
rect 19444 13348 20720 13376
rect 12989 13311 13047 13317
rect 12989 13277 13001 13311
rect 13035 13277 13047 13311
rect 12989 13271 13047 13277
rect 13078 13268 13084 13320
rect 13136 13268 13142 13320
rect 13357 13311 13415 13317
rect 13357 13277 13369 13311
rect 13403 13277 13415 13311
rect 13357 13271 13415 13277
rect 12728 13240 12756 13268
rect 13170 13240 13176 13252
rect 12728 13212 13176 13240
rect 13170 13200 13176 13212
rect 13228 13240 13234 13252
rect 13372 13240 13400 13271
rect 14366 13268 14372 13320
rect 14424 13268 14430 13320
rect 15194 13268 15200 13320
rect 15252 13268 15258 13320
rect 15286 13268 15292 13320
rect 15344 13268 15350 13320
rect 16316 13317 16344 13348
rect 16301 13311 16359 13317
rect 16301 13277 16313 13311
rect 16347 13277 16359 13311
rect 16301 13271 16359 13277
rect 16666 13268 16672 13320
rect 16724 13268 16730 13320
rect 16758 13268 16764 13320
rect 16816 13308 16822 13320
rect 16945 13311 17003 13317
rect 16945 13308 16957 13311
rect 16816 13280 16957 13308
rect 16816 13268 16822 13280
rect 16945 13277 16957 13280
rect 16991 13277 17003 13311
rect 16945 13271 17003 13277
rect 17218 13268 17224 13320
rect 17276 13268 17282 13320
rect 17313 13311 17371 13317
rect 17313 13277 17325 13311
rect 17359 13277 17371 13311
rect 17313 13271 17371 13277
rect 13228 13212 13400 13240
rect 13464 13212 16528 13240
rect 13228 13200 13234 13212
rect 12434 13172 12440 13184
rect 11716 13144 12440 13172
rect 10321 13135 10379 13141
rect 12434 13132 12440 13144
rect 12492 13132 12498 13184
rect 12986 13132 12992 13184
rect 13044 13172 13050 13184
rect 13464 13172 13492 13212
rect 13044 13144 13492 13172
rect 13541 13175 13599 13181
rect 13044 13132 13050 13144
rect 13541 13141 13553 13175
rect 13587 13172 13599 13175
rect 13722 13172 13728 13184
rect 13587 13144 13728 13172
rect 13587 13141 13599 13144
rect 13541 13135 13599 13141
rect 13722 13132 13728 13144
rect 13780 13132 13786 13184
rect 13814 13132 13820 13184
rect 13872 13172 13878 13184
rect 15013 13175 15071 13181
rect 15013 13172 15025 13175
rect 13872 13144 15025 13172
rect 13872 13132 13878 13144
rect 15013 13141 15025 13144
rect 15059 13141 15071 13175
rect 15013 13135 15071 13141
rect 15654 13132 15660 13184
rect 15712 13172 15718 13184
rect 16393 13175 16451 13181
rect 16393 13172 16405 13175
rect 15712 13144 16405 13172
rect 15712 13132 15718 13144
rect 16393 13141 16405 13144
rect 16439 13141 16451 13175
rect 16500 13172 16528 13212
rect 17126 13200 17132 13252
rect 17184 13240 17190 13252
rect 17328 13240 17356 13271
rect 17402 13268 17408 13320
rect 17460 13308 17466 13320
rect 17696 13308 17724 13348
rect 17460 13280 17724 13308
rect 17773 13311 17831 13317
rect 17460 13268 17466 13280
rect 17773 13277 17785 13311
rect 17819 13277 17831 13311
rect 17773 13271 17831 13277
rect 17184 13212 17356 13240
rect 17184 13200 17190 13212
rect 17494 13200 17500 13252
rect 17552 13200 17558 13252
rect 17586 13172 17592 13184
rect 16500 13144 17592 13172
rect 16393 13135 16451 13141
rect 17586 13132 17592 13144
rect 17644 13132 17650 13184
rect 17788 13172 17816 13271
rect 17862 13268 17868 13320
rect 17920 13268 17926 13320
rect 17954 13268 17960 13320
rect 18012 13308 18018 13320
rect 18506 13308 18512 13320
rect 18012 13280 18512 13308
rect 18012 13268 18018 13280
rect 18506 13268 18512 13280
rect 18564 13268 18570 13320
rect 18598 13268 18604 13320
rect 18656 13308 18662 13320
rect 19245 13311 19303 13317
rect 19245 13308 19257 13311
rect 18656 13280 19257 13308
rect 18656 13268 18662 13280
rect 19245 13277 19257 13280
rect 19291 13277 19303 13311
rect 19245 13271 19303 13277
rect 18049 13243 18107 13249
rect 18049 13209 18061 13243
rect 18095 13240 18107 13243
rect 18966 13240 18972 13252
rect 18095 13212 18972 13240
rect 18095 13209 18107 13212
rect 18049 13203 18107 13209
rect 18966 13200 18972 13212
rect 19024 13200 19030 13252
rect 19260 13240 19288 13271
rect 19334 13268 19340 13320
rect 19392 13268 19398 13320
rect 19444 13240 19472 13348
rect 20714 13336 20720 13348
rect 20772 13336 20778 13388
rect 21726 13376 21732 13388
rect 20916 13348 21732 13376
rect 20916 13320 20944 13348
rect 21726 13336 21732 13348
rect 21784 13376 21790 13388
rect 22094 13376 22100 13388
rect 21784 13348 22100 13376
rect 21784 13336 21790 13348
rect 22094 13336 22100 13348
rect 22152 13336 22158 13388
rect 19521 13311 19579 13317
rect 19521 13277 19533 13311
rect 19567 13277 19579 13311
rect 19521 13271 19579 13277
rect 19613 13311 19671 13317
rect 19613 13277 19625 13311
rect 19659 13308 19671 13311
rect 19978 13308 19984 13320
rect 19659 13280 19984 13308
rect 19659 13277 19671 13280
rect 19613 13271 19671 13277
rect 19260 13212 19472 13240
rect 18506 13172 18512 13184
rect 17788 13144 18512 13172
rect 18506 13132 18512 13144
rect 18564 13132 18570 13184
rect 18874 13132 18880 13184
rect 18932 13172 18938 13184
rect 19536 13172 19564 13271
rect 19978 13268 19984 13280
rect 20036 13268 20042 13320
rect 20070 13268 20076 13320
rect 20128 13268 20134 13320
rect 20346 13268 20352 13320
rect 20404 13268 20410 13320
rect 20898 13268 20904 13320
rect 20956 13268 20962 13320
rect 21085 13311 21143 13317
rect 21085 13277 21097 13311
rect 21131 13277 21143 13311
rect 21085 13271 21143 13277
rect 19794 13200 19800 13252
rect 19852 13200 19858 13252
rect 20257 13243 20315 13249
rect 20257 13209 20269 13243
rect 20303 13209 20315 13243
rect 20257 13203 20315 13209
rect 20272 13172 20300 13203
rect 20622 13200 20628 13252
rect 20680 13240 20686 13252
rect 21100 13240 21128 13271
rect 21174 13268 21180 13320
rect 21232 13268 21238 13320
rect 21269 13311 21327 13317
rect 21269 13277 21281 13311
rect 21315 13308 21327 13311
rect 21542 13308 21548 13320
rect 21315 13280 21548 13308
rect 21315 13277 21327 13280
rect 21269 13271 21327 13277
rect 21542 13268 21548 13280
rect 21600 13268 21606 13320
rect 22204 13308 22232 13484
rect 22370 13404 22376 13456
rect 22428 13444 22434 13456
rect 22428 13416 22508 13444
rect 22428 13404 22434 13416
rect 22112 13280 22232 13308
rect 22112 13240 22140 13280
rect 22370 13268 22376 13320
rect 22428 13268 22434 13320
rect 22480 13317 22508 13416
rect 22465 13311 22523 13317
rect 22465 13277 22477 13311
rect 22511 13277 22523 13311
rect 22465 13271 22523 13277
rect 22557 13311 22615 13317
rect 22557 13277 22569 13311
rect 22603 13308 22615 13311
rect 22664 13308 22692 13484
rect 23014 13472 23020 13524
rect 23072 13512 23078 13524
rect 23750 13512 23756 13524
rect 23072 13484 23756 13512
rect 23072 13472 23078 13484
rect 23750 13472 23756 13484
rect 23808 13472 23814 13524
rect 26326 13472 26332 13524
rect 26384 13512 26390 13524
rect 27065 13515 27123 13521
rect 27065 13512 27077 13515
rect 26384 13484 27077 13512
rect 26384 13472 26390 13484
rect 27065 13481 27077 13484
rect 27111 13481 27123 13515
rect 30466 13512 30472 13524
rect 27065 13475 27123 13481
rect 28276 13484 30472 13512
rect 28276 13456 28304 13484
rect 30466 13472 30472 13484
rect 30524 13472 30530 13524
rect 31754 13512 31760 13524
rect 31589 13484 31760 13512
rect 22738 13404 22744 13456
rect 22796 13444 22802 13456
rect 22833 13447 22891 13453
rect 22833 13444 22845 13447
rect 22796 13416 22845 13444
rect 22796 13404 22802 13416
rect 22833 13413 22845 13416
rect 22879 13413 22891 13447
rect 22833 13407 22891 13413
rect 27522 13404 27528 13456
rect 27580 13444 27586 13456
rect 28258 13444 28264 13456
rect 27580 13416 28264 13444
rect 27580 13404 27586 13416
rect 28258 13404 28264 13416
rect 28316 13404 28322 13456
rect 30009 13447 30067 13453
rect 30009 13413 30021 13447
rect 30055 13444 30067 13447
rect 31589 13444 31617 13484
rect 31754 13472 31760 13484
rect 31812 13472 31818 13524
rect 32122 13472 32128 13524
rect 32180 13512 32186 13524
rect 32398 13512 32404 13524
rect 32180 13484 32404 13512
rect 32180 13472 32186 13484
rect 32398 13472 32404 13484
rect 32456 13472 32462 13524
rect 34146 13472 34152 13524
rect 34204 13512 34210 13524
rect 34701 13515 34759 13521
rect 34701 13512 34713 13515
rect 34204 13484 34713 13512
rect 34204 13472 34210 13484
rect 34701 13481 34713 13484
rect 34747 13481 34759 13515
rect 34701 13475 34759 13481
rect 35161 13515 35219 13521
rect 35161 13481 35173 13515
rect 35207 13512 35219 13515
rect 36722 13512 36728 13524
rect 35207 13484 36728 13512
rect 35207 13481 35219 13484
rect 35161 13475 35219 13481
rect 36722 13472 36728 13484
rect 36780 13472 36786 13524
rect 36814 13472 36820 13524
rect 36872 13512 36878 13524
rect 36872 13484 38792 13512
rect 36872 13472 36878 13484
rect 31846 13444 31852 13456
rect 30055 13416 31617 13444
rect 31726 13416 31852 13444
rect 30055 13413 30067 13416
rect 30009 13407 30067 13413
rect 22922 13336 22928 13388
rect 22980 13376 22986 13388
rect 31726 13376 31754 13416
rect 31846 13404 31852 13416
rect 31904 13404 31910 13456
rect 32309 13447 32367 13453
rect 32309 13413 32321 13447
rect 32355 13444 32367 13447
rect 32766 13444 32772 13456
rect 32355 13416 32772 13444
rect 32355 13413 32367 13416
rect 32309 13407 32367 13413
rect 32766 13404 32772 13416
rect 32824 13404 32830 13456
rect 32858 13404 32864 13456
rect 32916 13404 32922 13456
rect 33226 13404 33232 13456
rect 33284 13404 33290 13456
rect 33413 13447 33471 13453
rect 33413 13413 33425 13447
rect 33459 13444 33471 13447
rect 38764 13444 38792 13484
rect 38930 13472 38936 13524
rect 38988 13472 38994 13524
rect 39117 13515 39175 13521
rect 39117 13481 39129 13515
rect 39163 13481 39175 13515
rect 39117 13475 39175 13481
rect 39132 13444 39160 13475
rect 33459 13416 37274 13444
rect 38764 13416 39160 13444
rect 33459 13413 33471 13416
rect 33413 13407 33471 13413
rect 32876 13376 32904 13404
rect 33244 13376 33272 13404
rect 22980 13348 31754 13376
rect 32692 13348 32904 13376
rect 33152 13348 33272 13376
rect 34885 13379 34943 13385
rect 22980 13336 22986 13348
rect 22603 13280 22692 13308
rect 22603 13277 22615 13280
rect 22557 13271 22615 13277
rect 20680 13212 22140 13240
rect 20680 13200 20686 13212
rect 18932 13144 20300 13172
rect 18932 13132 18938 13144
rect 21542 13132 21548 13184
rect 21600 13132 21606 13184
rect 22480 13172 22508 13271
rect 22664 13240 22692 13280
rect 22741 13311 22799 13317
rect 22741 13277 22753 13311
rect 22787 13308 22799 13311
rect 22830 13308 22836 13320
rect 22787 13280 22836 13308
rect 22787 13277 22799 13280
rect 22741 13271 22799 13277
rect 22830 13268 22836 13280
rect 22888 13268 22894 13320
rect 26142 13268 26148 13320
rect 26200 13268 26206 13320
rect 26234 13268 26240 13320
rect 26292 13268 26298 13320
rect 26602 13268 26608 13320
rect 26660 13268 26666 13320
rect 27154 13268 27160 13320
rect 27212 13268 27218 13320
rect 27982 13308 27988 13320
rect 27264 13280 27988 13308
rect 23201 13243 23259 13249
rect 23201 13240 23213 13243
rect 22664 13212 23213 13240
rect 23201 13209 23213 13212
rect 23247 13209 23259 13243
rect 23201 13203 23259 13209
rect 23382 13200 23388 13252
rect 23440 13240 23446 13252
rect 24854 13240 24860 13252
rect 23440 13212 24860 13240
rect 23440 13200 23446 13212
rect 24854 13200 24860 13212
rect 24912 13240 24918 13252
rect 25590 13240 25596 13252
rect 24912 13212 25596 13240
rect 24912 13200 24918 13212
rect 25590 13200 25596 13212
rect 25648 13240 25654 13252
rect 27264 13240 27292 13280
rect 27982 13268 27988 13280
rect 28040 13308 28046 13320
rect 30101 13311 30159 13317
rect 28040 13280 29408 13308
rect 28040 13268 28046 13280
rect 27798 13240 27804 13252
rect 25648 13212 27292 13240
rect 27356 13212 27804 13240
rect 25648 13200 25654 13212
rect 22830 13172 22836 13184
rect 22480 13144 22836 13172
rect 22830 13132 22836 13144
rect 22888 13132 22894 13184
rect 23014 13181 23020 13184
rect 23001 13175 23020 13181
rect 23001 13141 23013 13175
rect 23001 13135 23020 13141
rect 23014 13132 23020 13135
rect 23072 13132 23078 13184
rect 23106 13132 23112 13184
rect 23164 13172 23170 13184
rect 23400 13172 23428 13200
rect 23164 13144 23428 13172
rect 23164 13132 23170 13144
rect 24210 13132 24216 13184
rect 24268 13172 24274 13184
rect 25866 13172 25872 13184
rect 24268 13144 25872 13172
rect 24268 13132 24274 13144
rect 25866 13132 25872 13144
rect 25924 13172 25930 13184
rect 27356 13172 27384 13212
rect 27798 13200 27804 13212
rect 27856 13240 27862 13252
rect 29270 13240 29276 13252
rect 27856 13212 29276 13240
rect 27856 13200 27862 13212
rect 29270 13200 29276 13212
rect 29328 13200 29334 13252
rect 29380 13240 29408 13280
rect 30101 13277 30113 13311
rect 30147 13308 30159 13311
rect 30190 13308 30196 13320
rect 30147 13280 30196 13308
rect 30147 13277 30159 13280
rect 30101 13271 30159 13277
rect 30190 13268 30196 13280
rect 30248 13268 30254 13320
rect 30282 13268 30288 13320
rect 30340 13268 30346 13320
rect 31478 13268 31484 13320
rect 31536 13308 31542 13320
rect 31757 13311 31815 13317
rect 31757 13308 31769 13311
rect 31536 13280 31769 13308
rect 31536 13268 31542 13280
rect 31757 13277 31769 13280
rect 31803 13308 31815 13311
rect 31846 13308 31852 13320
rect 31803 13280 31852 13308
rect 31803 13277 31815 13280
rect 31757 13271 31815 13277
rect 31846 13268 31852 13280
rect 31904 13268 31910 13320
rect 32125 13311 32183 13317
rect 32125 13277 32137 13311
rect 32171 13277 32183 13311
rect 32125 13271 32183 13277
rect 31386 13240 31392 13252
rect 29380 13212 31392 13240
rect 31386 13200 31392 13212
rect 31444 13200 31450 13252
rect 31938 13200 31944 13252
rect 31996 13200 32002 13252
rect 32033 13243 32091 13249
rect 32033 13209 32045 13243
rect 32079 13209 32091 13243
rect 32033 13203 32091 13209
rect 25924 13144 27384 13172
rect 25924 13132 25930 13144
rect 27706 13132 27712 13184
rect 27764 13172 27770 13184
rect 28350 13172 28356 13184
rect 27764 13144 28356 13172
rect 27764 13132 27770 13144
rect 28350 13132 28356 13144
rect 28408 13132 28414 13184
rect 29178 13132 29184 13184
rect 29236 13172 29242 13184
rect 30926 13172 30932 13184
rect 29236 13144 30932 13172
rect 29236 13132 29242 13144
rect 30926 13132 30932 13144
rect 30984 13132 30990 13184
rect 31478 13132 31484 13184
rect 31536 13172 31542 13184
rect 32048 13172 32076 13203
rect 31536 13144 32076 13172
rect 32140 13172 32168 13271
rect 32490 13268 32496 13320
rect 32548 13268 32554 13320
rect 32692 13317 32720 13348
rect 32677 13311 32735 13317
rect 32677 13277 32689 13311
rect 32723 13277 32735 13311
rect 32677 13271 32735 13277
rect 32766 13268 32772 13320
rect 32824 13268 32830 13320
rect 33152 13317 33180 13348
rect 34885 13345 34897 13379
rect 34931 13376 34943 13379
rect 35434 13376 35440 13388
rect 34931 13348 35440 13376
rect 34931 13345 34943 13348
rect 34885 13339 34943 13345
rect 35434 13336 35440 13348
rect 35492 13336 35498 13388
rect 37246 13376 37274 13416
rect 38562 13376 38568 13388
rect 37246 13348 38568 13376
rect 38562 13336 38568 13348
rect 38620 13376 38626 13388
rect 39209 13379 39267 13385
rect 39209 13376 39221 13379
rect 38620 13348 39221 13376
rect 38620 13336 38626 13348
rect 39209 13345 39221 13348
rect 39255 13345 39267 13379
rect 39209 13339 39267 13345
rect 32862 13311 32920 13317
rect 32862 13277 32874 13311
rect 32908 13277 32920 13311
rect 32862 13271 32920 13277
rect 33137 13311 33195 13317
rect 33137 13277 33149 13311
rect 33183 13277 33195 13311
rect 33137 13271 33195 13277
rect 32508 13240 32536 13268
rect 32876 13240 32904 13271
rect 33226 13268 33232 13320
rect 33284 13317 33290 13320
rect 33284 13311 33333 13317
rect 33284 13277 33287 13311
rect 33321 13308 33333 13311
rect 33321 13280 34192 13308
rect 33321 13277 33333 13280
rect 33284 13271 33333 13277
rect 33284 13268 33290 13271
rect 32508 13212 32904 13240
rect 33042 13200 33048 13252
rect 33100 13240 33106 13252
rect 33962 13240 33968 13252
rect 33100 13212 33968 13240
rect 33100 13200 33106 13212
rect 33962 13200 33968 13212
rect 34020 13200 34026 13252
rect 32490 13172 32496 13184
rect 32140 13144 32496 13172
rect 31536 13132 31542 13144
rect 32490 13132 32496 13144
rect 32548 13132 32554 13184
rect 34164 13172 34192 13280
rect 34698 13268 34704 13320
rect 34756 13268 34762 13320
rect 34977 13311 35035 13317
rect 34977 13308 34989 13311
rect 34808 13280 34989 13308
rect 34808 13252 34836 13280
rect 34977 13277 34989 13280
rect 35023 13277 35035 13311
rect 34977 13271 35035 13277
rect 38102 13268 38108 13320
rect 38160 13308 38166 13320
rect 38749 13311 38807 13317
rect 38749 13308 38761 13311
rect 38160 13280 38761 13308
rect 38160 13268 38166 13280
rect 38749 13277 38761 13280
rect 38795 13277 38807 13311
rect 38749 13271 38807 13277
rect 38841 13311 38899 13317
rect 38841 13277 38853 13311
rect 38887 13277 38899 13311
rect 38841 13271 38899 13277
rect 39117 13311 39175 13317
rect 39117 13277 39129 13311
rect 39163 13302 39175 13311
rect 39850 13308 39856 13320
rect 39408 13302 39856 13308
rect 39163 13280 39856 13302
rect 39163 13277 39436 13280
rect 39117 13274 39436 13277
rect 39117 13271 39175 13274
rect 34790 13200 34796 13252
rect 34848 13200 34854 13252
rect 35342 13172 35348 13184
rect 34164 13144 35348 13172
rect 35342 13132 35348 13144
rect 35400 13132 35406 13184
rect 38102 13132 38108 13184
rect 38160 13172 38166 13184
rect 38565 13175 38623 13181
rect 38565 13172 38577 13175
rect 38160 13144 38577 13172
rect 38160 13132 38166 13144
rect 38565 13141 38577 13144
rect 38611 13141 38623 13175
rect 38565 13135 38623 13141
rect 38746 13132 38752 13184
rect 38804 13172 38810 13184
rect 38856 13172 38884 13271
rect 39850 13268 39856 13280
rect 39908 13268 39914 13320
rect 39025 13243 39083 13249
rect 39025 13209 39037 13243
rect 39071 13240 39083 13243
rect 39071 13212 39344 13240
rect 39071 13209 39083 13212
rect 39025 13203 39083 13209
rect 39316 13184 39344 13212
rect 38804 13144 38884 13172
rect 38804 13132 38810 13144
rect 39298 13132 39304 13184
rect 39356 13172 39362 13184
rect 39485 13175 39543 13181
rect 39485 13172 39497 13175
rect 39356 13144 39497 13172
rect 39356 13132 39362 13144
rect 39485 13141 39497 13144
rect 39531 13141 39543 13175
rect 39485 13135 39543 13141
rect 1104 13082 40572 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 40572 13082
rect 1104 13008 40572 13030
rect 3234 12968 3240 12980
rect 2148 12940 3240 12968
rect 2148 12841 2176 12940
rect 3234 12928 3240 12940
rect 3292 12928 3298 12980
rect 4614 12928 4620 12980
rect 4672 12928 4678 12980
rect 4706 12928 4712 12980
rect 4764 12968 4770 12980
rect 5169 12971 5227 12977
rect 5169 12968 5181 12971
rect 4764 12940 5181 12968
rect 4764 12928 4770 12940
rect 5169 12937 5181 12940
rect 5215 12937 5227 12971
rect 5169 12931 5227 12937
rect 6914 12928 6920 12980
rect 6972 12968 6978 12980
rect 7742 12968 7748 12980
rect 6972 12940 7748 12968
rect 6972 12928 6978 12940
rect 7742 12928 7748 12940
rect 7800 12968 7806 12980
rect 8481 12971 8539 12977
rect 8481 12968 8493 12971
rect 7800 12940 8493 12968
rect 7800 12928 7806 12940
rect 8481 12937 8493 12940
rect 8527 12937 8539 12971
rect 8481 12931 8539 12937
rect 10597 12971 10655 12977
rect 10597 12937 10609 12971
rect 10643 12937 10655 12971
rect 10597 12931 10655 12937
rect 11885 12971 11943 12977
rect 11885 12937 11897 12971
rect 11931 12968 11943 12971
rect 12434 12968 12440 12980
rect 11931 12940 12440 12968
rect 11931 12937 11943 12940
rect 11885 12931 11943 12937
rect 3786 12900 3792 12912
rect 3634 12872 3792 12900
rect 3786 12860 3792 12872
rect 3844 12860 3850 12912
rect 4632 12900 4660 12928
rect 7377 12903 7435 12909
rect 4632 12872 5672 12900
rect 2133 12835 2191 12841
rect 2133 12801 2145 12835
rect 2179 12801 2191 12835
rect 2133 12795 2191 12801
rect 4338 12792 4344 12844
rect 4396 12792 4402 12844
rect 4430 12792 4436 12844
rect 4488 12792 4494 12844
rect 4614 12792 4620 12844
rect 4672 12792 4678 12844
rect 4709 12835 4767 12841
rect 4709 12801 4721 12835
rect 4755 12832 4767 12835
rect 4890 12832 4896 12844
rect 4755 12804 4896 12832
rect 4755 12801 4767 12804
rect 4709 12795 4767 12801
rect 4890 12792 4896 12804
rect 4948 12792 4954 12844
rect 5444 12835 5502 12841
rect 5444 12801 5456 12835
rect 5490 12801 5502 12835
rect 5444 12795 5502 12801
rect 2409 12767 2467 12773
rect 2409 12733 2421 12767
rect 2455 12764 2467 12767
rect 4157 12767 4215 12773
rect 4157 12764 4169 12767
rect 2455 12736 4169 12764
rect 2455 12733 2467 12736
rect 2409 12727 2467 12733
rect 4157 12733 4169 12736
rect 4203 12733 4215 12767
rect 5460 12764 5488 12795
rect 5534 12792 5540 12844
rect 5592 12792 5598 12844
rect 5644 12841 5672 12872
rect 7377 12869 7389 12903
rect 7423 12900 7435 12903
rect 7466 12900 7472 12912
rect 7423 12872 7472 12900
rect 7423 12869 7435 12872
rect 7377 12863 7435 12869
rect 7466 12860 7472 12872
rect 7524 12860 7530 12912
rect 10612 12900 10640 12931
rect 12434 12928 12440 12940
rect 12492 12928 12498 12980
rect 12526 12928 12532 12980
rect 12584 12928 12590 12980
rect 13170 12928 13176 12980
rect 13228 12928 13234 12980
rect 15378 12968 15384 12980
rect 14768 12940 15384 12968
rect 7760 12872 10640 12900
rect 5629 12835 5687 12841
rect 5629 12801 5641 12835
rect 5675 12832 5687 12835
rect 5902 12832 5908 12844
rect 5675 12804 5908 12832
rect 5675 12801 5687 12804
rect 5629 12795 5687 12801
rect 5902 12792 5908 12804
rect 5960 12792 5966 12844
rect 6914 12792 6920 12844
rect 6972 12832 6978 12844
rect 6972 12804 7052 12832
rect 6972 12792 6978 12804
rect 5460 12736 5672 12764
rect 4157 12727 4215 12733
rect 4430 12656 4436 12708
rect 4488 12696 4494 12708
rect 5258 12696 5264 12708
rect 4488 12668 5264 12696
rect 4488 12656 4494 12668
rect 5258 12656 5264 12668
rect 5316 12656 5322 12708
rect 5644 12696 5672 12736
rect 5718 12724 5724 12776
rect 5776 12724 5782 12776
rect 6730 12764 6736 12776
rect 5828 12736 6736 12764
rect 5828 12696 5856 12736
rect 6730 12724 6736 12736
rect 6788 12724 6794 12776
rect 7024 12773 7052 12804
rect 7098 12792 7104 12844
rect 7156 12792 7162 12844
rect 7282 12792 7288 12844
rect 7340 12832 7346 12844
rect 7760 12841 7788 12872
rect 11514 12860 11520 12912
rect 11572 12900 11578 12912
rect 11572 12872 12020 12900
rect 11572 12860 11578 12872
rect 7653 12835 7711 12841
rect 7653 12832 7665 12835
rect 7340 12804 7665 12832
rect 7340 12792 7346 12804
rect 7653 12801 7665 12804
rect 7699 12801 7711 12835
rect 7653 12795 7711 12801
rect 7745 12835 7803 12841
rect 7745 12801 7757 12835
rect 7791 12801 7803 12835
rect 7745 12795 7803 12801
rect 7834 12792 7840 12844
rect 7892 12792 7898 12844
rect 8018 12792 8024 12844
rect 8076 12792 8082 12844
rect 8294 12792 8300 12844
rect 8352 12792 8358 12844
rect 8570 12792 8576 12844
rect 8628 12792 8634 12844
rect 10226 12792 10232 12844
rect 10284 12832 10290 12844
rect 10781 12835 10839 12841
rect 10781 12832 10793 12835
rect 10284 12804 10793 12832
rect 10284 12792 10290 12804
rect 10781 12801 10793 12804
rect 10827 12801 10839 12835
rect 10781 12795 10839 12801
rect 10873 12835 10931 12841
rect 10873 12801 10885 12835
rect 10919 12832 10931 12835
rect 10962 12832 10968 12844
rect 10919 12804 10968 12832
rect 10919 12801 10931 12804
rect 10873 12795 10931 12801
rect 10962 12792 10968 12804
rect 11020 12792 11026 12844
rect 11241 12835 11299 12841
rect 11241 12801 11253 12835
rect 11287 12832 11299 12835
rect 11701 12835 11759 12841
rect 11701 12832 11713 12835
rect 11287 12804 11713 12832
rect 11287 12801 11299 12804
rect 11241 12795 11299 12801
rect 11701 12801 11713 12804
rect 11747 12832 11759 12835
rect 11790 12832 11796 12844
rect 11747 12804 11796 12832
rect 11747 12801 11759 12804
rect 11701 12795 11759 12801
rect 11790 12792 11796 12804
rect 11848 12792 11854 12844
rect 11992 12841 12020 12872
rect 12406 12872 13492 12900
rect 11977 12835 12035 12841
rect 11977 12801 11989 12835
rect 12023 12801 12035 12835
rect 12406 12832 12434 12872
rect 11977 12795 12035 12801
rect 12084 12804 12434 12832
rect 12897 12835 12955 12841
rect 7009 12767 7067 12773
rect 7009 12733 7021 12767
rect 7055 12733 7067 12767
rect 7009 12727 7067 12733
rect 9674 12724 9680 12776
rect 9732 12764 9738 12776
rect 11054 12764 11060 12776
rect 9732 12736 11060 12764
rect 9732 12724 9738 12736
rect 11054 12724 11060 12736
rect 11112 12764 11118 12776
rect 11149 12767 11207 12773
rect 11149 12764 11161 12767
rect 11112 12736 11161 12764
rect 11112 12724 11118 12736
rect 11149 12733 11161 12736
rect 11195 12733 11207 12767
rect 12084 12764 12112 12804
rect 12897 12801 12909 12835
rect 12943 12832 12955 12835
rect 12986 12832 12992 12844
rect 12943 12804 12992 12832
rect 12943 12801 12955 12804
rect 12897 12795 12955 12801
rect 12986 12792 12992 12804
rect 13044 12792 13050 12844
rect 13265 12835 13323 12841
rect 13265 12801 13277 12835
rect 13311 12801 13323 12835
rect 13265 12795 13323 12801
rect 11149 12727 11207 12733
rect 11256 12736 12112 12764
rect 7558 12696 7564 12708
rect 5644 12668 5856 12696
rect 5920 12668 7564 12696
rect 3881 12631 3939 12637
rect 3881 12597 3893 12631
rect 3927 12628 3939 12631
rect 5442 12628 5448 12640
rect 3927 12600 5448 12628
rect 3927 12597 3939 12600
rect 3881 12591 3939 12597
rect 5442 12588 5448 12600
rect 5500 12588 5506 12640
rect 5810 12588 5816 12640
rect 5868 12628 5874 12640
rect 5920 12628 5948 12668
rect 7558 12656 7564 12668
rect 7616 12696 7622 12708
rect 8662 12696 8668 12708
rect 7616 12668 8668 12696
rect 7616 12656 7622 12668
rect 8662 12656 8668 12668
rect 8720 12656 8726 12708
rect 8938 12656 8944 12708
rect 8996 12696 9002 12708
rect 11256 12696 11284 12736
rect 12342 12724 12348 12776
rect 12400 12764 12406 12776
rect 13280 12764 13308 12795
rect 12400 12736 13308 12764
rect 12400 12724 12406 12736
rect 8996 12668 11284 12696
rect 8996 12656 9002 12668
rect 11330 12656 11336 12708
rect 11388 12696 11394 12708
rect 11517 12699 11575 12705
rect 11517 12696 11529 12699
rect 11388 12668 11529 12696
rect 11388 12656 11394 12668
rect 11517 12665 11529 12668
rect 11563 12665 11575 12699
rect 11517 12659 11575 12665
rect 12805 12699 12863 12705
rect 12805 12665 12817 12699
rect 12851 12696 12863 12699
rect 13354 12696 13360 12708
rect 12851 12668 13360 12696
rect 12851 12665 12863 12668
rect 12805 12659 12863 12665
rect 13354 12656 13360 12668
rect 13412 12656 13418 12708
rect 13464 12696 13492 12872
rect 13722 12792 13728 12844
rect 13780 12792 13786 12844
rect 14093 12835 14151 12841
rect 14093 12801 14105 12835
rect 14139 12832 14151 12835
rect 14366 12832 14372 12844
rect 14139 12804 14372 12832
rect 14139 12801 14151 12804
rect 14093 12795 14151 12801
rect 14366 12792 14372 12804
rect 14424 12792 14430 12844
rect 14550 12792 14556 12844
rect 14608 12792 14614 12844
rect 14768 12841 14796 12940
rect 15378 12928 15384 12940
rect 15436 12968 15442 12980
rect 15436 12940 17448 12968
rect 15436 12928 15442 12940
rect 16666 12860 16672 12912
rect 16724 12900 16730 12912
rect 17420 12900 17448 12940
rect 17494 12928 17500 12980
rect 17552 12928 17558 12980
rect 17586 12928 17592 12980
rect 17644 12968 17650 12980
rect 18598 12968 18604 12980
rect 17644 12940 18604 12968
rect 17644 12928 17650 12940
rect 18598 12928 18604 12940
rect 18656 12928 18662 12980
rect 18966 12928 18972 12980
rect 19024 12968 19030 12980
rect 19702 12968 19708 12980
rect 19024 12940 19708 12968
rect 19024 12928 19030 12940
rect 19702 12928 19708 12940
rect 19760 12928 19766 12980
rect 20162 12928 20168 12980
rect 20220 12968 20226 12980
rect 20806 12968 20812 12980
rect 20220 12940 20812 12968
rect 20220 12928 20226 12940
rect 20806 12928 20812 12940
rect 20864 12928 20870 12980
rect 20990 12928 20996 12980
rect 21048 12928 21054 12980
rect 21082 12928 21088 12980
rect 21140 12968 21146 12980
rect 21634 12968 21640 12980
rect 21140 12940 21640 12968
rect 21140 12928 21146 12940
rect 21634 12928 21640 12940
rect 21692 12968 21698 12980
rect 21692 12940 22232 12968
rect 21692 12928 21698 12940
rect 16724 12872 17356 12900
rect 17420 12872 18828 12900
rect 16724 12860 16730 12872
rect 14737 12835 14796 12841
rect 14737 12801 14749 12835
rect 14783 12804 14796 12835
rect 14783 12801 14795 12804
rect 14737 12795 14795 12801
rect 15286 12792 15292 12844
rect 15344 12832 15350 12844
rect 16945 12835 17003 12841
rect 16945 12832 16957 12835
rect 15344 12804 16957 12832
rect 15344 12792 15350 12804
rect 16945 12801 16957 12804
rect 16991 12832 17003 12835
rect 17328 12832 17356 12872
rect 17405 12835 17463 12841
rect 17405 12832 17417 12835
rect 16991 12804 17264 12832
rect 17328 12804 17417 12832
rect 16991 12801 17003 12804
rect 16945 12795 17003 12801
rect 17034 12724 17040 12776
rect 17092 12764 17098 12776
rect 17129 12767 17187 12773
rect 17129 12764 17141 12767
rect 17092 12736 17141 12764
rect 17092 12724 17098 12736
rect 17129 12733 17141 12736
rect 17175 12733 17187 12767
rect 17236 12764 17264 12804
rect 17405 12801 17417 12804
rect 17451 12801 17463 12835
rect 17405 12795 17463 12801
rect 17310 12764 17316 12776
rect 17236 12736 17316 12764
rect 17129 12727 17187 12733
rect 17310 12724 17316 12736
rect 17368 12724 17374 12776
rect 17420 12764 17448 12795
rect 17678 12792 17684 12844
rect 17736 12792 17742 12844
rect 17770 12792 17776 12844
rect 17828 12792 17834 12844
rect 17954 12792 17960 12844
rect 18012 12792 18018 12844
rect 18046 12792 18052 12844
rect 18104 12792 18110 12844
rect 18506 12792 18512 12844
rect 18564 12792 18570 12844
rect 17420 12736 18000 12764
rect 17972 12708 18000 12736
rect 18690 12724 18696 12776
rect 18748 12724 18754 12776
rect 18800 12764 18828 12872
rect 18874 12860 18880 12912
rect 18932 12900 18938 12912
rect 21821 12903 21879 12909
rect 21821 12900 21833 12903
rect 18932 12872 21833 12900
rect 18932 12860 18938 12872
rect 21821 12869 21833 12872
rect 21867 12869 21879 12903
rect 21821 12863 21879 12869
rect 18966 12792 18972 12844
rect 19024 12792 19030 12844
rect 20070 12792 20076 12844
rect 20128 12832 20134 12844
rect 21177 12835 21235 12841
rect 21177 12832 21189 12835
rect 20128 12804 21189 12832
rect 20128 12792 20134 12804
rect 21177 12801 21189 12804
rect 21223 12801 21235 12835
rect 21177 12795 21235 12801
rect 21358 12792 21364 12844
rect 21416 12832 21422 12844
rect 21545 12835 21603 12841
rect 21545 12832 21557 12835
rect 21416 12804 21557 12832
rect 21416 12792 21422 12804
rect 21545 12801 21557 12804
rect 21591 12801 21603 12835
rect 21545 12795 21603 12801
rect 21376 12764 21404 12792
rect 18800 12736 21404 12764
rect 21836 12764 21864 12863
rect 22094 12792 22100 12844
rect 22152 12792 22158 12844
rect 22204 12832 22232 12940
rect 22922 12928 22928 12980
rect 22980 12928 22986 12980
rect 23198 12928 23204 12980
rect 23256 12968 23262 12980
rect 26973 12971 27031 12977
rect 26973 12968 26985 12971
rect 23256 12940 23428 12968
rect 23256 12928 23262 12940
rect 22940 12900 22968 12928
rect 23400 12909 23428 12940
rect 24136 12940 26985 12968
rect 22480 12872 22968 12900
rect 23385 12903 23443 12909
rect 22281 12835 22339 12841
rect 22281 12832 22293 12835
rect 22204 12804 22293 12832
rect 22281 12801 22293 12804
rect 22327 12801 22339 12835
rect 22281 12795 22339 12801
rect 22370 12792 22376 12844
rect 22428 12832 22434 12844
rect 22480 12832 22508 12872
rect 23385 12869 23397 12903
rect 23431 12869 23443 12903
rect 23385 12863 23443 12869
rect 22428 12804 22508 12832
rect 22557 12835 22615 12841
rect 22428 12792 22434 12804
rect 22557 12801 22569 12835
rect 22603 12832 22615 12835
rect 22738 12832 22744 12844
rect 22603 12804 22744 12832
rect 22603 12801 22615 12804
rect 22557 12795 22615 12801
rect 22738 12792 22744 12804
rect 22796 12792 22802 12844
rect 22833 12835 22891 12841
rect 22833 12801 22845 12835
rect 22879 12832 22891 12835
rect 22922 12832 22928 12844
rect 22879 12804 22928 12832
rect 22879 12801 22891 12804
rect 22833 12795 22891 12801
rect 22922 12792 22928 12804
rect 22980 12832 22986 12844
rect 23201 12835 23259 12841
rect 23201 12832 23213 12835
rect 22980 12804 23213 12832
rect 22980 12792 22986 12804
rect 23201 12801 23213 12804
rect 23247 12801 23259 12835
rect 23201 12795 23259 12801
rect 23474 12792 23480 12844
rect 23532 12792 23538 12844
rect 23842 12792 23848 12844
rect 23900 12792 23906 12844
rect 23934 12792 23940 12844
rect 23992 12792 23998 12844
rect 24136 12841 24164 12940
rect 26973 12937 26985 12940
rect 27019 12937 27031 12971
rect 26973 12931 27031 12937
rect 28902 12928 28908 12980
rect 28960 12928 28966 12980
rect 29086 12928 29092 12980
rect 29144 12928 29150 12980
rect 29730 12928 29736 12980
rect 29788 12968 29794 12980
rect 30098 12968 30104 12980
rect 29788 12940 30104 12968
rect 29788 12928 29794 12940
rect 30098 12928 30104 12940
rect 30156 12968 30162 12980
rect 31205 12971 31263 12977
rect 31205 12968 31217 12971
rect 30156 12940 31217 12968
rect 30156 12928 30162 12940
rect 31205 12937 31217 12940
rect 31251 12937 31263 12971
rect 31205 12931 31263 12937
rect 32677 12971 32735 12977
rect 32677 12937 32689 12971
rect 32723 12968 32735 12971
rect 32950 12968 32956 12980
rect 32723 12940 32956 12968
rect 32723 12937 32735 12940
rect 32677 12931 32735 12937
rect 32950 12928 32956 12940
rect 33008 12928 33014 12980
rect 35437 12971 35495 12977
rect 35437 12937 35449 12971
rect 35483 12968 35495 12971
rect 38378 12968 38384 12980
rect 35483 12940 38384 12968
rect 35483 12937 35495 12940
rect 35437 12931 35495 12937
rect 38378 12928 38384 12940
rect 38436 12928 38442 12980
rect 38654 12928 38660 12980
rect 38712 12928 38718 12980
rect 25958 12900 25964 12912
rect 25332 12872 25964 12900
rect 24121 12835 24179 12841
rect 24121 12801 24133 12835
rect 24167 12801 24179 12835
rect 24121 12795 24179 12801
rect 24578 12792 24584 12844
rect 24636 12792 24642 12844
rect 24673 12835 24731 12841
rect 24673 12801 24685 12835
rect 24719 12832 24731 12835
rect 24854 12832 24860 12844
rect 24719 12804 24860 12832
rect 24719 12801 24731 12804
rect 24673 12795 24731 12801
rect 24854 12792 24860 12804
rect 24912 12792 24918 12844
rect 25332 12841 25360 12872
rect 25958 12860 25964 12872
rect 26016 12900 26022 12912
rect 26510 12900 26516 12912
rect 26016 12872 26516 12900
rect 26016 12860 26022 12872
rect 26510 12860 26516 12872
rect 26568 12860 26574 12912
rect 26786 12860 26792 12912
rect 26844 12900 26850 12912
rect 27341 12903 27399 12909
rect 27341 12900 27353 12903
rect 26844 12872 27353 12900
rect 26844 12860 26850 12872
rect 27341 12869 27353 12872
rect 27387 12869 27399 12903
rect 27341 12863 27399 12869
rect 28000 12872 29224 12900
rect 25041 12835 25099 12841
rect 25041 12801 25053 12835
rect 25087 12832 25099 12835
rect 25317 12835 25375 12841
rect 25317 12832 25329 12835
rect 25087 12804 25329 12832
rect 25087 12801 25099 12804
rect 25041 12795 25099 12801
rect 25317 12801 25329 12804
rect 25363 12801 25375 12835
rect 25317 12795 25375 12801
rect 25590 12792 25596 12844
rect 25648 12792 25654 12844
rect 27157 12835 27215 12841
rect 27157 12801 27169 12835
rect 27203 12801 27215 12835
rect 27157 12795 27215 12801
rect 22186 12764 22192 12776
rect 21836 12736 22192 12764
rect 22186 12724 22192 12736
rect 22244 12724 22250 12776
rect 23109 12767 23167 12773
rect 23109 12733 23121 12767
rect 23155 12764 23167 12767
rect 23492 12764 23520 12792
rect 23155 12736 23520 12764
rect 24765 12767 24823 12773
rect 23155 12733 23167 12736
rect 23109 12727 23167 12733
rect 24765 12733 24777 12767
rect 24811 12764 24823 12767
rect 25222 12764 25228 12776
rect 24811 12736 25228 12764
rect 24811 12733 24823 12736
rect 24765 12727 24823 12733
rect 25222 12724 25228 12736
rect 25280 12764 25286 12776
rect 25409 12767 25467 12773
rect 25409 12764 25421 12767
rect 25280 12736 25421 12764
rect 25280 12724 25286 12736
rect 25409 12733 25421 12736
rect 25455 12733 25467 12767
rect 27172 12764 27200 12795
rect 27246 12792 27252 12844
rect 27304 12792 27310 12844
rect 27522 12792 27528 12844
rect 27580 12792 27586 12844
rect 27617 12835 27675 12841
rect 27617 12801 27629 12835
rect 27663 12830 27675 12835
rect 27706 12830 27712 12844
rect 27663 12802 27712 12830
rect 27663 12801 27675 12802
rect 27617 12795 27675 12801
rect 27706 12792 27712 12802
rect 27764 12792 27770 12844
rect 27890 12764 27896 12776
rect 27172 12736 27896 12764
rect 25409 12727 25467 12733
rect 27890 12724 27896 12736
rect 27948 12724 27954 12776
rect 14277 12699 14335 12705
rect 13464 12668 14228 12696
rect 5868 12600 5948 12628
rect 5997 12631 6055 12637
rect 5868 12588 5874 12600
rect 5997 12597 6009 12631
rect 6043 12628 6055 12631
rect 6178 12628 6184 12640
rect 6043 12600 6184 12628
rect 6043 12597 6055 12600
rect 5997 12591 6055 12597
rect 6178 12588 6184 12600
rect 6236 12588 6242 12640
rect 6362 12588 6368 12640
rect 6420 12628 6426 12640
rect 8018 12628 8024 12640
rect 6420 12600 8024 12628
rect 6420 12588 6426 12600
rect 8018 12588 8024 12600
rect 8076 12588 8082 12640
rect 8110 12588 8116 12640
rect 8168 12588 8174 12640
rect 11606 12588 11612 12640
rect 11664 12628 11670 12640
rect 12342 12628 12348 12640
rect 11664 12600 12348 12628
rect 11664 12588 11670 12600
rect 12342 12588 12348 12600
rect 12400 12588 12406 12640
rect 12989 12631 13047 12637
rect 12989 12597 13001 12631
rect 13035 12628 13047 12631
rect 13262 12628 13268 12640
rect 13035 12600 13268 12628
rect 13035 12597 13047 12600
rect 12989 12591 13047 12597
rect 13262 12588 13268 12600
rect 13320 12588 13326 12640
rect 14090 12588 14096 12640
rect 14148 12588 14154 12640
rect 14200 12628 14228 12668
rect 14277 12665 14289 12699
rect 14323 12696 14335 12699
rect 15194 12696 15200 12708
rect 14323 12668 15200 12696
rect 14323 12665 14335 12668
rect 14277 12659 14335 12665
rect 15194 12656 15200 12668
rect 15252 12656 15258 12708
rect 17402 12696 17408 12708
rect 17052 12668 17408 12696
rect 14461 12631 14519 12637
rect 14461 12628 14473 12631
rect 14200 12600 14473 12628
rect 14461 12597 14473 12600
rect 14507 12597 14519 12631
rect 14461 12591 14519 12597
rect 16666 12588 16672 12640
rect 16724 12588 16730 12640
rect 17052 12637 17080 12668
rect 17402 12656 17408 12668
rect 17460 12656 17466 12708
rect 17954 12656 17960 12708
rect 18012 12656 18018 12708
rect 22649 12699 22707 12705
rect 22649 12696 22661 12699
rect 18248 12668 22661 12696
rect 17037 12631 17095 12637
rect 17037 12597 17049 12631
rect 17083 12597 17095 12631
rect 17037 12591 17095 12597
rect 17218 12588 17224 12640
rect 17276 12628 17282 12640
rect 18248 12628 18276 12668
rect 22649 12665 22661 12668
rect 22695 12665 22707 12699
rect 23382 12696 23388 12708
rect 22649 12659 22707 12665
rect 22756 12668 23388 12696
rect 17276 12600 18276 12628
rect 17276 12588 17282 12600
rect 18322 12588 18328 12640
rect 18380 12588 18386 12640
rect 18877 12631 18935 12637
rect 18877 12597 18889 12631
rect 18923 12628 18935 12631
rect 19794 12628 19800 12640
rect 18923 12600 19800 12628
rect 18923 12597 18935 12600
rect 18877 12591 18935 12597
rect 19794 12588 19800 12600
rect 19852 12588 19858 12640
rect 21453 12631 21511 12637
rect 21453 12597 21465 12631
rect 21499 12628 21511 12631
rect 21542 12628 21548 12640
rect 21499 12600 21548 12628
rect 21499 12597 21511 12600
rect 21453 12591 21511 12597
rect 21542 12588 21548 12600
rect 21600 12588 21606 12640
rect 21726 12588 21732 12640
rect 21784 12628 21790 12640
rect 22189 12631 22247 12637
rect 22189 12628 22201 12631
rect 21784 12600 22201 12628
rect 21784 12588 21790 12600
rect 22189 12597 22201 12600
rect 22235 12628 22247 12631
rect 22756 12628 22784 12668
rect 23382 12656 23388 12668
rect 23440 12656 23446 12708
rect 24029 12699 24087 12705
rect 23584 12668 23980 12696
rect 22235 12600 22784 12628
rect 23017 12631 23075 12637
rect 22235 12597 22247 12600
rect 22189 12591 22247 12597
rect 23017 12597 23029 12631
rect 23063 12628 23075 12631
rect 23584 12628 23612 12668
rect 23063 12600 23612 12628
rect 23661 12631 23719 12637
rect 23063 12597 23075 12600
rect 23017 12591 23075 12597
rect 23661 12597 23673 12631
rect 23707 12628 23719 12631
rect 23842 12628 23848 12640
rect 23707 12600 23848 12628
rect 23707 12597 23719 12600
rect 23661 12591 23719 12597
rect 23842 12588 23848 12600
rect 23900 12588 23906 12640
rect 23952 12628 23980 12668
rect 24029 12665 24041 12699
rect 24075 12696 24087 12699
rect 24305 12699 24363 12705
rect 24305 12696 24317 12699
rect 24075 12668 24317 12696
rect 24075 12665 24087 12668
rect 24029 12659 24087 12665
rect 24305 12665 24317 12668
rect 24351 12665 24363 12699
rect 24305 12659 24363 12665
rect 27522 12656 27528 12708
rect 27580 12696 27586 12708
rect 28000 12696 28028 12872
rect 29196 12844 29224 12872
rect 29270 12860 29276 12912
rect 29328 12900 29334 12912
rect 29328 12872 29500 12900
rect 29328 12860 29334 12872
rect 28074 12792 28080 12844
rect 28132 12792 28138 12844
rect 28169 12835 28227 12841
rect 28169 12801 28181 12835
rect 28215 12832 28227 12835
rect 28258 12832 28264 12844
rect 28215 12804 28264 12832
rect 28215 12801 28227 12804
rect 28169 12795 28227 12801
rect 27580 12668 28028 12696
rect 27580 12656 27586 12668
rect 28074 12656 28080 12708
rect 28132 12696 28138 12708
rect 28184 12696 28212 12795
rect 28258 12792 28264 12804
rect 28316 12792 28322 12844
rect 28350 12792 28356 12844
rect 28408 12792 28414 12844
rect 28537 12835 28595 12841
rect 28537 12801 28549 12835
rect 28583 12801 28595 12835
rect 28537 12795 28595 12801
rect 28552 12764 28580 12795
rect 28718 12792 28724 12844
rect 28776 12792 28782 12844
rect 28810 12792 28816 12844
rect 28868 12832 28874 12844
rect 28997 12835 29055 12841
rect 28997 12832 29009 12835
rect 28868 12804 29009 12832
rect 28868 12792 28874 12804
rect 28997 12801 29009 12804
rect 29043 12801 29055 12835
rect 28997 12795 29055 12801
rect 29178 12792 29184 12844
rect 29236 12792 29242 12844
rect 29472 12832 29500 12872
rect 29914 12860 29920 12912
rect 29972 12900 29978 12912
rect 29972 12872 30696 12900
rect 29972 12860 29978 12872
rect 30009 12835 30067 12841
rect 30009 12832 30021 12835
rect 29472 12804 30021 12832
rect 30009 12801 30021 12804
rect 30055 12801 30067 12835
rect 30009 12795 30067 12801
rect 30098 12792 30104 12844
rect 30156 12832 30162 12844
rect 30193 12835 30251 12841
rect 30193 12832 30205 12835
rect 30156 12804 30205 12832
rect 30156 12792 30162 12804
rect 30193 12801 30205 12804
rect 30239 12801 30251 12835
rect 30193 12795 30251 12801
rect 30466 12792 30472 12844
rect 30524 12792 30530 12844
rect 30561 12835 30619 12841
rect 30561 12801 30573 12835
rect 30607 12801 30619 12835
rect 30561 12795 30619 12801
rect 30668 12822 30696 12872
rect 30926 12860 30932 12912
rect 30984 12900 30990 12912
rect 30984 12872 31340 12900
rect 30984 12860 30990 12872
rect 30745 12835 30803 12841
rect 30745 12822 30757 12835
rect 30668 12801 30757 12822
rect 30791 12801 30803 12835
rect 30668 12795 30803 12801
rect 28276 12736 28580 12764
rect 28276 12708 28304 12736
rect 29730 12724 29736 12776
rect 29788 12724 29794 12776
rect 30282 12724 30288 12776
rect 30340 12764 30346 12776
rect 30576 12764 30604 12795
rect 30668 12794 30782 12795
rect 30834 12792 30840 12844
rect 30892 12792 30898 12844
rect 31036 12841 31064 12872
rect 31312 12841 31340 12872
rect 31386 12860 31392 12912
rect 31444 12900 31450 12912
rect 35161 12903 35219 12909
rect 35161 12900 35173 12903
rect 31444 12872 35173 12900
rect 31444 12860 31450 12872
rect 35161 12869 35173 12872
rect 35207 12869 35219 12903
rect 35161 12863 35219 12869
rect 35342 12860 35348 12912
rect 35400 12900 35406 12912
rect 35526 12900 35532 12912
rect 35400 12872 35532 12900
rect 35400 12860 35406 12872
rect 35526 12860 35532 12872
rect 35584 12860 35590 12912
rect 38672 12900 38700 12928
rect 38672 12872 38976 12900
rect 31021 12835 31079 12841
rect 31021 12801 31033 12835
rect 31067 12801 31079 12835
rect 31021 12795 31079 12801
rect 31119 12835 31177 12841
rect 31119 12801 31131 12835
rect 31165 12822 31177 12835
rect 31297 12835 31355 12841
rect 31165 12801 31202 12822
rect 31119 12795 31202 12801
rect 31297 12801 31309 12835
rect 31343 12801 31355 12835
rect 31754 12832 31760 12844
rect 31297 12795 31355 12801
rect 31404 12804 31760 12832
rect 31128 12794 31202 12795
rect 30340 12736 30604 12764
rect 30929 12767 30987 12773
rect 30340 12724 30346 12736
rect 30929 12733 30941 12767
rect 30975 12733 30987 12767
rect 31174 12764 31202 12794
rect 31404 12764 31432 12804
rect 31754 12792 31760 12804
rect 31812 12792 31818 12844
rect 31846 12792 31852 12844
rect 31904 12832 31910 12844
rect 32125 12835 32183 12841
rect 32125 12832 32137 12835
rect 31904 12804 32137 12832
rect 31904 12792 31910 12804
rect 32125 12801 32137 12804
rect 32171 12801 32183 12835
rect 32125 12795 32183 12801
rect 32214 12792 32220 12844
rect 32272 12832 32278 12844
rect 32309 12835 32367 12841
rect 32309 12832 32321 12835
rect 32272 12804 32321 12832
rect 32272 12792 32278 12804
rect 32309 12801 32321 12804
rect 32355 12801 32367 12835
rect 32309 12795 32367 12801
rect 32401 12835 32459 12841
rect 32401 12801 32413 12835
rect 32447 12801 32459 12835
rect 32401 12795 32459 12801
rect 31174 12736 31432 12764
rect 30929 12727 30987 12733
rect 28132 12668 28212 12696
rect 28132 12656 28138 12668
rect 28258 12656 28264 12708
rect 28316 12656 28322 12708
rect 28350 12656 28356 12708
rect 28408 12696 28414 12708
rect 28408 12668 28994 12696
rect 28408 12656 28414 12668
rect 24486 12628 24492 12640
rect 23952 12600 24492 12628
rect 24486 12588 24492 12600
rect 24544 12588 24550 12640
rect 24854 12588 24860 12640
rect 24912 12588 24918 12640
rect 25133 12631 25191 12637
rect 25133 12597 25145 12631
rect 25179 12628 25191 12631
rect 25314 12628 25320 12640
rect 25179 12600 25320 12628
rect 25179 12597 25191 12600
rect 25133 12591 25191 12597
rect 25314 12588 25320 12600
rect 25372 12588 25378 12640
rect 25593 12631 25651 12637
rect 25593 12597 25605 12631
rect 25639 12628 25651 12631
rect 25866 12628 25872 12640
rect 25639 12600 25872 12628
rect 25639 12597 25651 12600
rect 25593 12591 25651 12597
rect 25866 12588 25872 12600
rect 25924 12588 25930 12640
rect 27798 12588 27804 12640
rect 27856 12628 27862 12640
rect 27893 12631 27951 12637
rect 27893 12628 27905 12631
rect 27856 12600 27905 12628
rect 27856 12588 27862 12600
rect 27893 12597 27905 12600
rect 27939 12597 27951 12631
rect 27893 12591 27951 12597
rect 27982 12588 27988 12640
rect 28040 12628 28046 12640
rect 28810 12628 28816 12640
rect 28040 12600 28816 12628
rect 28040 12588 28046 12600
rect 28810 12588 28816 12600
rect 28868 12588 28874 12640
rect 28966 12628 28994 12668
rect 30006 12656 30012 12708
rect 30064 12696 30070 12708
rect 30300 12696 30328 12724
rect 30944 12696 30972 12727
rect 30064 12668 30328 12696
rect 30392 12668 30972 12696
rect 30064 12656 30070 12668
rect 30392 12640 30420 12668
rect 31202 12656 31208 12708
rect 31260 12696 31266 12708
rect 32416 12696 32444 12795
rect 32490 12792 32496 12844
rect 32548 12832 32554 12844
rect 32950 12832 32956 12844
rect 32548 12804 32956 12832
rect 32548 12792 32554 12804
rect 32950 12792 32956 12804
rect 33008 12832 33014 12844
rect 33226 12832 33232 12844
rect 33008 12804 33232 12832
rect 33008 12792 33014 12804
rect 33226 12792 33232 12804
rect 33284 12792 33290 12844
rect 34790 12792 34796 12844
rect 34848 12792 34854 12844
rect 34886 12835 34944 12841
rect 34886 12801 34898 12835
rect 34932 12801 34944 12835
rect 34886 12795 34944 12801
rect 35069 12835 35127 12841
rect 35069 12801 35081 12835
rect 35115 12801 35127 12835
rect 35069 12795 35127 12801
rect 35258 12835 35316 12841
rect 35258 12801 35270 12835
rect 35304 12832 35316 12835
rect 35360 12832 35388 12860
rect 35304 12804 35388 12832
rect 35304 12801 35316 12804
rect 35258 12795 35316 12801
rect 33502 12724 33508 12776
rect 33560 12764 33566 12776
rect 34606 12764 34612 12776
rect 33560 12736 34612 12764
rect 33560 12724 33566 12736
rect 34606 12724 34612 12736
rect 34664 12764 34670 12776
rect 34901 12764 34929 12795
rect 34664 12736 34929 12764
rect 35084 12764 35112 12795
rect 38654 12792 38660 12844
rect 38712 12792 38718 12844
rect 38948 12841 38976 12872
rect 38933 12835 38991 12841
rect 38933 12801 38945 12835
rect 38979 12801 38991 12835
rect 38933 12795 38991 12801
rect 36078 12764 36084 12776
rect 35084 12736 36084 12764
rect 34664 12724 34670 12736
rect 36078 12724 36084 12736
rect 36136 12724 36142 12776
rect 38562 12724 38568 12776
rect 38620 12764 38626 12776
rect 38749 12767 38807 12773
rect 38749 12764 38761 12767
rect 38620 12736 38761 12764
rect 38620 12724 38626 12736
rect 38749 12733 38761 12736
rect 38795 12733 38807 12767
rect 38749 12727 38807 12733
rect 39482 12696 39488 12708
rect 31260 12668 32444 12696
rect 38948 12668 39488 12696
rect 31260 12656 31266 12668
rect 29086 12628 29092 12640
rect 28966 12600 29092 12628
rect 29086 12588 29092 12600
rect 29144 12628 29150 12640
rect 30101 12631 30159 12637
rect 30101 12628 30113 12631
rect 29144 12600 30113 12628
rect 29144 12588 29150 12600
rect 30101 12597 30113 12600
rect 30147 12597 30159 12631
rect 30101 12591 30159 12597
rect 30285 12631 30343 12637
rect 30285 12597 30297 12631
rect 30331 12628 30343 12631
rect 30374 12628 30380 12640
rect 30331 12600 30380 12628
rect 30331 12597 30343 12600
rect 30285 12591 30343 12597
rect 30374 12588 30380 12600
rect 30432 12588 30438 12640
rect 30466 12588 30472 12640
rect 30524 12628 30530 12640
rect 38948 12637 38976 12668
rect 39482 12656 39488 12668
rect 39540 12656 39546 12708
rect 30745 12631 30803 12637
rect 30745 12628 30757 12631
rect 30524 12600 30757 12628
rect 30524 12588 30530 12600
rect 30745 12597 30757 12600
rect 30791 12597 30803 12631
rect 30745 12591 30803 12597
rect 38933 12631 38991 12637
rect 38933 12597 38945 12631
rect 38979 12597 38991 12631
rect 38933 12591 38991 12597
rect 39114 12588 39120 12640
rect 39172 12588 39178 12640
rect 1104 12538 40572 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 40572 12538
rect 1104 12464 40572 12486
rect 4433 12427 4491 12433
rect 4433 12393 4445 12427
rect 4479 12424 4491 12427
rect 4706 12424 4712 12436
rect 4479 12396 4712 12424
rect 4479 12393 4491 12396
rect 4433 12387 4491 12393
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 5442 12424 5448 12436
rect 4816 12396 5448 12424
rect 4341 12359 4399 12365
rect 4341 12325 4353 12359
rect 4387 12356 4399 12359
rect 4614 12356 4620 12368
rect 4387 12328 4620 12356
rect 4387 12325 4399 12328
rect 4341 12319 4399 12325
rect 4614 12316 4620 12328
rect 4672 12316 4678 12368
rect 4065 12291 4123 12297
rect 4065 12257 4077 12291
rect 4111 12288 4123 12291
rect 4706 12288 4712 12300
rect 4111 12260 4712 12288
rect 4111 12257 4123 12260
rect 4065 12251 4123 12257
rect 4706 12248 4712 12260
rect 4764 12248 4770 12300
rect 4816 12297 4844 12396
rect 5442 12384 5448 12396
rect 5500 12384 5506 12436
rect 6362 12384 6368 12436
rect 6420 12384 6426 12436
rect 6454 12384 6460 12436
rect 6512 12424 6518 12436
rect 7009 12427 7067 12433
rect 7009 12424 7021 12427
rect 6512 12396 7021 12424
rect 6512 12384 6518 12396
rect 5902 12356 5908 12368
rect 4908 12328 5908 12356
rect 4801 12291 4859 12297
rect 4801 12257 4813 12291
rect 4847 12257 4859 12291
rect 4801 12251 4859 12257
rect 3970 12180 3976 12232
rect 4028 12180 4034 12232
rect 4617 12223 4675 12229
rect 4617 12189 4629 12223
rect 4663 12220 4675 12223
rect 4908 12220 4936 12328
rect 5902 12316 5908 12328
rect 5960 12356 5966 12368
rect 6270 12356 6276 12368
rect 5960 12328 6276 12356
rect 5960 12316 5966 12328
rect 6270 12316 6276 12328
rect 6328 12316 6334 12368
rect 5534 12248 5540 12300
rect 5592 12288 5598 12300
rect 6086 12288 6092 12300
rect 5592 12260 6092 12288
rect 5592 12248 5598 12260
rect 6086 12248 6092 12260
rect 6144 12248 6150 12300
rect 6564 12297 6592 12396
rect 7009 12393 7021 12396
rect 7055 12393 7067 12427
rect 7009 12387 7067 12393
rect 7653 12427 7711 12433
rect 7653 12393 7665 12427
rect 7699 12424 7711 12427
rect 7834 12424 7840 12436
rect 7699 12396 7840 12424
rect 7699 12393 7711 12396
rect 7653 12387 7711 12393
rect 7834 12384 7840 12396
rect 7892 12384 7898 12436
rect 12989 12427 13047 12433
rect 12989 12393 13001 12427
rect 13035 12424 13047 12427
rect 13078 12424 13084 12436
rect 13035 12396 13084 12424
rect 13035 12393 13047 12396
rect 12989 12387 13047 12393
rect 13078 12384 13084 12396
rect 13136 12384 13142 12436
rect 17954 12384 17960 12436
rect 18012 12384 18018 12436
rect 18966 12424 18972 12436
rect 18616 12396 18972 12424
rect 17034 12316 17040 12368
rect 17092 12316 17098 12368
rect 18230 12316 18236 12368
rect 18288 12356 18294 12368
rect 18616 12356 18644 12396
rect 18966 12384 18972 12396
rect 19024 12384 19030 12436
rect 19242 12384 19248 12436
rect 19300 12384 19306 12436
rect 19334 12384 19340 12436
rect 19392 12384 19398 12436
rect 19518 12384 19524 12436
rect 19576 12384 19582 12436
rect 19702 12384 19708 12436
rect 19760 12424 19766 12436
rect 19797 12427 19855 12433
rect 19797 12424 19809 12427
rect 19760 12396 19809 12424
rect 19760 12384 19766 12396
rect 19797 12393 19809 12396
rect 19843 12393 19855 12427
rect 19797 12387 19855 12393
rect 19886 12384 19892 12436
rect 19944 12424 19950 12436
rect 20165 12427 20223 12433
rect 20165 12424 20177 12427
rect 19944 12396 20177 12424
rect 19944 12384 19950 12396
rect 20165 12393 20177 12396
rect 20211 12393 20223 12427
rect 20165 12387 20223 12393
rect 20257 12427 20315 12433
rect 20257 12393 20269 12427
rect 20303 12424 20315 12427
rect 20346 12424 20352 12436
rect 20303 12396 20352 12424
rect 20303 12393 20315 12396
rect 20257 12387 20315 12393
rect 20346 12384 20352 12396
rect 20404 12384 20410 12436
rect 21266 12384 21272 12436
rect 21324 12424 21330 12436
rect 21726 12424 21732 12436
rect 21324 12396 21732 12424
rect 21324 12384 21330 12396
rect 21726 12384 21732 12396
rect 21784 12384 21790 12436
rect 26237 12427 26295 12433
rect 26237 12424 26249 12427
rect 23952 12396 26249 12424
rect 18288 12328 18644 12356
rect 18288 12316 18294 12328
rect 18690 12316 18696 12368
rect 18748 12356 18754 12368
rect 19260 12356 19288 12384
rect 18748 12328 19288 12356
rect 18748 12316 18754 12328
rect 23382 12316 23388 12368
rect 23440 12356 23446 12368
rect 23842 12356 23848 12368
rect 23440 12328 23848 12356
rect 23440 12316 23446 12328
rect 23842 12316 23848 12328
rect 23900 12316 23906 12368
rect 6549 12291 6607 12297
rect 6549 12257 6561 12291
rect 6595 12257 6607 12291
rect 6549 12251 6607 12257
rect 7006 12248 7012 12300
rect 7064 12288 7070 12300
rect 7193 12291 7251 12297
rect 7193 12288 7205 12291
rect 7064 12260 7205 12288
rect 7064 12248 7070 12260
rect 7193 12257 7205 12260
rect 7239 12257 7251 12291
rect 7193 12251 7251 12257
rect 7282 12248 7288 12300
rect 7340 12288 7346 12300
rect 7340 12260 7788 12288
rect 7340 12248 7346 12260
rect 7760 12232 7788 12260
rect 14550 12248 14556 12300
rect 14608 12288 14614 12300
rect 16761 12291 16819 12297
rect 16761 12288 16773 12291
rect 14608 12260 16773 12288
rect 14608 12248 14614 12260
rect 16761 12257 16773 12260
rect 16807 12257 16819 12291
rect 17052 12288 17080 12316
rect 19426 12288 19432 12300
rect 17052 12260 19432 12288
rect 16761 12251 16819 12257
rect 4663 12192 4936 12220
rect 5629 12223 5687 12229
rect 4663 12189 4675 12192
rect 4617 12183 4675 12189
rect 5629 12189 5641 12223
rect 5675 12220 5687 12223
rect 5675 12192 6132 12220
rect 5675 12189 5687 12192
rect 5629 12183 5687 12189
rect 5718 12112 5724 12164
rect 5776 12112 5782 12164
rect 5813 12155 5871 12161
rect 5813 12121 5825 12155
rect 5859 12121 5871 12155
rect 5813 12115 5871 12121
rect 3786 12044 3792 12096
rect 3844 12084 3850 12096
rect 5445 12087 5503 12093
rect 5445 12084 5457 12087
rect 3844 12056 5457 12084
rect 3844 12044 3850 12056
rect 5445 12053 5457 12056
rect 5491 12053 5503 12087
rect 5828 12084 5856 12115
rect 5902 12112 5908 12164
rect 5960 12161 5966 12164
rect 5960 12155 5989 12161
rect 5977 12121 5989 12155
rect 6104 12152 6132 12192
rect 6178 12180 6184 12232
rect 6236 12180 6242 12232
rect 6638 12180 6644 12232
rect 6696 12180 6702 12232
rect 6730 12180 6736 12232
rect 6788 12220 6794 12232
rect 6917 12223 6975 12229
rect 6917 12220 6929 12223
rect 6788 12192 6929 12220
rect 6788 12180 6794 12192
rect 6917 12189 6929 12192
rect 6963 12189 6975 12223
rect 6917 12183 6975 12189
rect 7558 12180 7564 12232
rect 7616 12180 7622 12232
rect 7742 12180 7748 12232
rect 7800 12180 7806 12232
rect 12618 12180 12624 12232
rect 12676 12220 12682 12232
rect 12805 12223 12863 12229
rect 12805 12220 12817 12223
rect 12676 12192 12817 12220
rect 12676 12180 12682 12192
rect 12805 12189 12817 12192
rect 12851 12189 12863 12223
rect 12805 12183 12863 12189
rect 12894 12180 12900 12232
rect 12952 12180 12958 12232
rect 13906 12180 13912 12232
rect 13964 12220 13970 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13964 12192 14105 12220
rect 13964 12180 13970 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14093 12183 14151 12189
rect 14737 12223 14795 12229
rect 14737 12189 14749 12223
rect 14783 12220 14795 12223
rect 14829 12223 14887 12229
rect 14829 12220 14841 12223
rect 14783 12192 14841 12220
rect 14783 12189 14795 12192
rect 14737 12183 14795 12189
rect 14829 12189 14841 12192
rect 14875 12189 14887 12223
rect 14829 12183 14887 12189
rect 15194 12180 15200 12232
rect 15252 12180 15258 12232
rect 17037 12223 17095 12229
rect 17037 12189 17049 12223
rect 17083 12220 17095 12223
rect 17310 12220 17316 12232
rect 17083 12192 17316 12220
rect 17083 12189 17095 12192
rect 17037 12183 17095 12189
rect 17310 12180 17316 12192
rect 17368 12180 17374 12232
rect 17512 12229 17540 12260
rect 19426 12248 19432 12260
rect 19484 12248 19490 12300
rect 20162 12248 20168 12300
rect 20220 12288 20226 12300
rect 20349 12291 20407 12297
rect 20349 12288 20361 12291
rect 20220 12260 20361 12288
rect 20220 12248 20226 12260
rect 20349 12257 20361 12260
rect 20395 12288 20407 12291
rect 23952 12288 23980 12396
rect 26237 12393 26249 12396
rect 26283 12424 26295 12427
rect 26283 12396 28994 12424
rect 26283 12393 26295 12396
rect 26237 12387 26295 12393
rect 27893 12359 27951 12365
rect 27893 12325 27905 12359
rect 27939 12356 27951 12359
rect 28074 12356 28080 12368
rect 27939 12328 28080 12356
rect 27939 12325 27951 12328
rect 27893 12319 27951 12325
rect 28074 12316 28080 12328
rect 28132 12316 28138 12368
rect 28966 12356 28994 12396
rect 29454 12384 29460 12436
rect 29512 12424 29518 12436
rect 30101 12427 30159 12433
rect 30101 12424 30113 12427
rect 29512 12396 30113 12424
rect 29512 12384 29518 12396
rect 30101 12393 30113 12396
rect 30147 12393 30159 12427
rect 30101 12387 30159 12393
rect 30745 12427 30803 12433
rect 30745 12393 30757 12427
rect 30791 12424 30803 12427
rect 30926 12424 30932 12436
rect 30791 12396 30932 12424
rect 30791 12393 30803 12396
rect 30745 12387 30803 12393
rect 30926 12384 30932 12396
rect 30984 12384 30990 12436
rect 33413 12427 33471 12433
rect 33413 12393 33425 12427
rect 33459 12424 33471 12427
rect 33778 12424 33784 12436
rect 33459 12396 33784 12424
rect 33459 12393 33471 12396
rect 33413 12387 33471 12393
rect 33778 12384 33784 12396
rect 33836 12384 33842 12436
rect 34790 12384 34796 12436
rect 34848 12424 34854 12436
rect 35345 12427 35403 12433
rect 35345 12424 35357 12427
rect 34848 12396 35357 12424
rect 34848 12384 34854 12396
rect 35345 12393 35357 12396
rect 35391 12393 35403 12427
rect 35345 12387 35403 12393
rect 37182 12384 37188 12436
rect 37240 12424 37246 12436
rect 38105 12427 38163 12433
rect 38105 12424 38117 12427
rect 37240 12396 38117 12424
rect 37240 12384 37246 12396
rect 38105 12393 38117 12396
rect 38151 12393 38163 12427
rect 38105 12387 38163 12393
rect 38565 12427 38623 12433
rect 38565 12393 38577 12427
rect 38611 12424 38623 12427
rect 38654 12424 38660 12436
rect 38611 12396 38660 12424
rect 38611 12393 38623 12396
rect 38565 12387 38623 12393
rect 38654 12384 38660 12396
rect 38712 12384 38718 12436
rect 33870 12356 33876 12368
rect 28966 12328 33876 12356
rect 33870 12316 33876 12328
rect 33928 12316 33934 12368
rect 37826 12356 37832 12368
rect 34440 12328 37832 12356
rect 30006 12288 30012 12300
rect 20395 12260 23980 12288
rect 26160 12260 30012 12288
rect 20395 12257 20407 12260
rect 20349 12251 20407 12257
rect 17497 12223 17555 12229
rect 17497 12189 17509 12223
rect 17543 12189 17555 12223
rect 17497 12183 17555 12189
rect 17865 12223 17923 12229
rect 17865 12189 17877 12223
rect 17911 12189 17923 12223
rect 17865 12183 17923 12189
rect 18141 12223 18199 12229
rect 18141 12189 18153 12223
rect 18187 12220 18199 12223
rect 18506 12220 18512 12232
rect 18187 12192 18512 12220
rect 18187 12189 18199 12192
rect 18141 12183 18199 12189
rect 8110 12152 8116 12164
rect 6104 12124 8116 12152
rect 5960 12115 5989 12121
rect 5960 12112 5966 12115
rect 8110 12112 8116 12124
rect 8168 12112 8174 12164
rect 10502 12112 10508 12164
rect 10560 12152 10566 12164
rect 15013 12155 15071 12161
rect 15013 12152 15025 12155
rect 10560 12124 15025 12152
rect 10560 12112 10566 12124
rect 14844 12096 14872 12124
rect 15013 12121 15025 12124
rect 15059 12121 15071 12155
rect 15013 12115 15071 12121
rect 15102 12112 15108 12164
rect 15160 12112 15166 12164
rect 17880 12152 17908 12183
rect 18506 12180 18512 12192
rect 18564 12220 18570 12232
rect 18601 12223 18659 12229
rect 18601 12220 18613 12223
rect 18564 12192 18613 12220
rect 18564 12180 18570 12192
rect 18601 12189 18613 12192
rect 18647 12189 18659 12223
rect 18601 12183 18659 12189
rect 18785 12223 18843 12229
rect 18785 12189 18797 12223
rect 18831 12220 18843 12223
rect 18874 12220 18880 12232
rect 18831 12192 18880 12220
rect 18831 12189 18843 12192
rect 18785 12183 18843 12189
rect 18874 12180 18880 12192
rect 18932 12180 18938 12232
rect 18966 12180 18972 12232
rect 19024 12220 19030 12232
rect 19024 12192 19748 12220
rect 19024 12180 19030 12192
rect 18325 12155 18383 12161
rect 18325 12152 18337 12155
rect 17880 12124 18337 12152
rect 18325 12121 18337 12124
rect 18371 12152 18383 12155
rect 19334 12152 19340 12164
rect 18371 12124 19340 12152
rect 18371 12121 18383 12124
rect 18325 12115 18383 12121
rect 19334 12112 19340 12124
rect 19392 12112 19398 12164
rect 19720 12161 19748 12192
rect 19794 12180 19800 12232
rect 19852 12220 19858 12232
rect 20073 12223 20131 12229
rect 20073 12220 20085 12223
rect 19852 12192 20085 12220
rect 19852 12180 19858 12192
rect 20073 12189 20085 12192
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 19705 12155 19763 12161
rect 19705 12121 19717 12155
rect 19751 12121 19763 12155
rect 20088 12152 20116 12183
rect 20530 12180 20536 12232
rect 20588 12180 20594 12232
rect 20625 12223 20683 12229
rect 20625 12189 20637 12223
rect 20671 12220 20683 12223
rect 22370 12220 22376 12232
rect 20671 12192 22376 12220
rect 20671 12189 20683 12192
rect 20625 12183 20683 12189
rect 21008 12164 21036 12192
rect 22370 12180 22376 12192
rect 22428 12220 22434 12232
rect 22922 12220 22928 12232
rect 22428 12192 22928 12220
rect 22428 12180 22434 12192
rect 22922 12180 22928 12192
rect 22980 12180 22986 12232
rect 26050 12180 26056 12232
rect 26108 12220 26114 12232
rect 26160 12220 26188 12260
rect 30006 12248 30012 12260
rect 30064 12248 30070 12300
rect 33502 12288 33508 12300
rect 33152 12260 33508 12288
rect 26108 12192 26188 12220
rect 26237 12223 26295 12229
rect 26108 12180 26114 12192
rect 26237 12189 26249 12223
rect 26283 12220 26295 12223
rect 26326 12220 26332 12232
rect 26283 12192 26332 12220
rect 26283 12189 26295 12192
rect 26237 12183 26295 12189
rect 26326 12180 26332 12192
rect 26384 12180 26390 12232
rect 27890 12180 27896 12232
rect 27948 12180 27954 12232
rect 28077 12223 28135 12229
rect 28077 12189 28089 12223
rect 28123 12189 28135 12223
rect 28077 12183 28135 12189
rect 20088 12124 20852 12152
rect 19705 12115 19763 12121
rect 6825 12087 6883 12093
rect 6825 12084 6837 12087
rect 5828 12056 6837 12084
rect 5445 12047 5503 12053
rect 6825 12053 6837 12056
rect 6871 12053 6883 12087
rect 6825 12047 6883 12053
rect 7466 12044 7472 12096
rect 7524 12044 7530 12096
rect 8570 12044 8576 12096
rect 8628 12084 8634 12096
rect 9490 12084 9496 12096
rect 8628 12056 9496 12084
rect 8628 12044 8634 12056
rect 9490 12044 9496 12056
rect 9548 12084 9554 12096
rect 12802 12084 12808 12096
rect 9548 12056 12808 12084
rect 9548 12044 9554 12056
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 14826 12044 14832 12096
rect 14884 12044 14890 12096
rect 15194 12044 15200 12096
rect 15252 12084 15258 12096
rect 15381 12087 15439 12093
rect 15381 12084 15393 12087
rect 15252 12056 15393 12084
rect 15252 12044 15258 12056
rect 15381 12053 15393 12056
rect 15427 12053 15439 12087
rect 15381 12047 15439 12053
rect 18598 12044 18604 12096
rect 18656 12084 18662 12096
rect 19150 12084 19156 12096
rect 18656 12056 19156 12084
rect 18656 12044 18662 12056
rect 19150 12044 19156 12056
rect 19208 12044 19214 12096
rect 19521 12087 19579 12093
rect 19521 12053 19533 12087
rect 19567 12084 19579 12087
rect 20714 12084 20720 12096
rect 19567 12056 20720 12084
rect 19567 12053 19579 12056
rect 19521 12047 19579 12053
rect 20714 12044 20720 12056
rect 20772 12044 20778 12096
rect 20824 12093 20852 12124
rect 20990 12112 20996 12164
rect 21048 12112 21054 12164
rect 26418 12112 26424 12164
rect 26476 12152 26482 12164
rect 28092 12152 28120 12183
rect 28534 12180 28540 12232
rect 28592 12220 28598 12232
rect 29914 12220 29920 12232
rect 28592 12192 29920 12220
rect 28592 12180 28598 12192
rect 29914 12180 29920 12192
rect 29972 12180 29978 12232
rect 30098 12180 30104 12232
rect 30156 12180 30162 12232
rect 30653 12223 30711 12229
rect 30653 12189 30665 12223
rect 30699 12189 30711 12223
rect 30653 12183 30711 12189
rect 26476 12124 28994 12152
rect 26476 12112 26482 12124
rect 20809 12087 20867 12093
rect 20809 12053 20821 12087
rect 20855 12053 20867 12087
rect 20809 12047 20867 12053
rect 22186 12044 22192 12096
rect 22244 12084 22250 12096
rect 25130 12084 25136 12096
rect 22244 12056 25136 12084
rect 22244 12044 22250 12056
rect 25130 12044 25136 12056
rect 25188 12084 25194 12096
rect 28718 12084 28724 12096
rect 25188 12056 28724 12084
rect 25188 12044 25194 12056
rect 28718 12044 28724 12056
rect 28776 12044 28782 12096
rect 28966 12084 28994 12124
rect 29454 12084 29460 12096
rect 28966 12056 29460 12084
rect 29454 12044 29460 12056
rect 29512 12044 29518 12096
rect 29932 12084 29960 12180
rect 30668 12152 30696 12183
rect 30742 12180 30748 12232
rect 30800 12180 30806 12232
rect 33152 12229 33180 12260
rect 33502 12248 33508 12260
rect 33560 12248 33566 12300
rect 33781 12291 33839 12297
rect 33781 12257 33793 12291
rect 33827 12288 33839 12291
rect 34440 12288 34468 12328
rect 37826 12316 37832 12328
rect 37884 12316 37890 12368
rect 33827 12260 34468 12288
rect 33827 12257 33839 12260
rect 33781 12251 33839 12257
rect 33137 12223 33195 12229
rect 33137 12189 33149 12223
rect 33183 12189 33195 12223
rect 33137 12183 33195 12189
rect 33226 12180 33232 12232
rect 33284 12220 33290 12232
rect 33597 12223 33655 12229
rect 33597 12220 33609 12223
rect 33284 12192 33609 12220
rect 33284 12180 33290 12192
rect 33597 12189 33609 12192
rect 33643 12189 33655 12223
rect 33597 12183 33655 12189
rect 30834 12152 30840 12164
rect 30668 12124 30840 12152
rect 30834 12112 30840 12124
rect 30892 12152 30898 12164
rect 33796 12152 33824 12251
rect 34606 12248 34612 12300
rect 34664 12288 34670 12300
rect 34701 12291 34759 12297
rect 34701 12288 34713 12291
rect 34664 12260 34713 12288
rect 34664 12248 34670 12260
rect 34701 12257 34713 12260
rect 34747 12257 34759 12291
rect 36630 12288 36636 12300
rect 34701 12251 34759 12257
rect 35084 12260 36636 12288
rect 33962 12180 33968 12232
rect 34020 12220 34026 12232
rect 34859 12223 34917 12229
rect 34859 12220 34871 12223
rect 34020 12192 34871 12220
rect 34020 12180 34026 12192
rect 34859 12189 34871 12192
rect 34905 12220 34917 12223
rect 35084 12220 35112 12260
rect 36630 12248 36636 12260
rect 36688 12248 36694 12300
rect 38289 12291 38347 12297
rect 38289 12257 38301 12291
rect 38335 12288 38347 12291
rect 39574 12288 39580 12300
rect 38335 12260 39580 12288
rect 38335 12257 38347 12260
rect 38289 12251 38347 12257
rect 39574 12248 39580 12260
rect 39632 12248 39638 12300
rect 34905 12192 35112 12220
rect 35161 12223 35219 12229
rect 34905 12189 34917 12192
rect 34859 12183 34917 12189
rect 35161 12189 35173 12223
rect 35207 12220 35219 12223
rect 35342 12220 35348 12232
rect 35207 12192 35348 12220
rect 35207 12189 35219 12192
rect 35161 12183 35219 12189
rect 35342 12180 35348 12192
rect 35400 12180 35406 12232
rect 35526 12180 35532 12232
rect 35584 12220 35590 12232
rect 35713 12223 35771 12229
rect 35713 12220 35725 12223
rect 35584 12192 35725 12220
rect 35584 12180 35590 12192
rect 35713 12189 35725 12192
rect 35759 12189 35771 12223
rect 35713 12183 35771 12189
rect 38378 12180 38384 12232
rect 38436 12180 38442 12232
rect 30892 12124 33824 12152
rect 30892 12112 30898 12124
rect 34514 12112 34520 12164
rect 34572 12152 34578 12164
rect 34698 12152 34704 12164
rect 34572 12124 34704 12152
rect 34572 12112 34578 12124
rect 34698 12112 34704 12124
rect 34756 12112 34762 12164
rect 34977 12155 35035 12161
rect 34977 12121 34989 12155
rect 35023 12121 35035 12155
rect 34977 12115 35035 12121
rect 31294 12084 31300 12096
rect 29932 12056 31300 12084
rect 31294 12044 31300 12056
rect 31352 12084 31358 12096
rect 31754 12084 31760 12096
rect 31352 12056 31760 12084
rect 31352 12044 31358 12056
rect 31754 12044 31760 12056
rect 31812 12044 31818 12096
rect 34238 12044 34244 12096
rect 34296 12084 34302 12096
rect 34882 12084 34888 12096
rect 34296 12056 34888 12084
rect 34296 12044 34302 12056
rect 34882 12044 34888 12056
rect 34940 12044 34946 12096
rect 34992 12084 35020 12115
rect 35066 12112 35072 12164
rect 35124 12112 35130 12164
rect 35360 12152 35388 12180
rect 35360 12124 35572 12152
rect 35250 12084 35256 12096
rect 34992 12056 35256 12084
rect 35250 12044 35256 12056
rect 35308 12084 35314 12096
rect 35434 12084 35440 12096
rect 35308 12056 35440 12084
rect 35308 12044 35314 12056
rect 35434 12044 35440 12056
rect 35492 12044 35498 12096
rect 35544 12093 35572 12124
rect 38102 12112 38108 12164
rect 38160 12112 38166 12164
rect 35529 12087 35587 12093
rect 35529 12053 35541 12087
rect 35575 12053 35587 12087
rect 35529 12047 35587 12053
rect 1104 11994 40572 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 40572 11994
rect 1104 11920 40572 11942
rect 4154 11840 4160 11892
rect 4212 11880 4218 11892
rect 4706 11880 4712 11892
rect 4212 11852 4712 11880
rect 4212 11840 4218 11852
rect 4706 11840 4712 11852
rect 4764 11840 4770 11892
rect 5261 11883 5319 11889
rect 5261 11849 5273 11883
rect 5307 11880 5319 11883
rect 5534 11880 5540 11892
rect 5307 11852 5540 11880
rect 5307 11849 5319 11852
rect 5261 11843 5319 11849
rect 5534 11840 5540 11852
rect 5592 11840 5598 11892
rect 5718 11840 5724 11892
rect 5776 11880 5782 11892
rect 6365 11883 6423 11889
rect 6365 11880 6377 11883
rect 5776 11852 6377 11880
rect 5776 11840 5782 11852
rect 6365 11849 6377 11852
rect 6411 11849 6423 11883
rect 6365 11843 6423 11849
rect 6546 11840 6552 11892
rect 6604 11880 6610 11892
rect 10502 11880 10508 11892
rect 6604 11852 10508 11880
rect 6604 11840 6610 11852
rect 10502 11840 10508 11852
rect 10560 11840 10566 11892
rect 14458 11880 14464 11892
rect 13924 11852 14464 11880
rect 3786 11772 3792 11824
rect 3844 11772 3850 11824
rect 4172 11812 4200 11840
rect 4172 11784 4278 11812
rect 7650 11772 7656 11824
rect 7708 11812 7714 11824
rect 7708 11784 8616 11812
rect 7708 11772 7714 11784
rect 6640 11747 6698 11753
rect 6640 11713 6652 11747
rect 6686 11713 6698 11747
rect 6640 11707 6698 11713
rect 3234 11636 3240 11688
rect 3292 11676 3298 11688
rect 3510 11676 3516 11688
rect 3292 11648 3516 11676
rect 3292 11636 3298 11648
rect 3510 11636 3516 11648
rect 3568 11636 3574 11688
rect 6656 11676 6684 11707
rect 6730 11704 6736 11756
rect 6788 11704 6794 11756
rect 8294 11704 8300 11756
rect 8352 11744 8358 11756
rect 8588 11753 8616 11784
rect 8846 11772 8852 11824
rect 8904 11772 8910 11824
rect 9493 11815 9551 11821
rect 9493 11781 9505 11815
rect 9539 11812 9551 11815
rect 9582 11812 9588 11824
rect 9539 11784 9588 11812
rect 9539 11781 9551 11784
rect 9493 11775 9551 11781
rect 9582 11772 9588 11784
rect 9640 11812 9646 11824
rect 9640 11784 10180 11812
rect 9640 11772 9646 11784
rect 8481 11747 8539 11753
rect 8481 11744 8493 11747
rect 8352 11716 8493 11744
rect 8352 11704 8358 11716
rect 8481 11713 8493 11716
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 8574 11747 8632 11753
rect 8574 11713 8586 11747
rect 8620 11713 8632 11747
rect 8574 11707 8632 11713
rect 8754 11704 8760 11756
rect 8812 11704 8818 11756
rect 8987 11747 9045 11753
rect 8987 11713 8999 11747
rect 9033 11744 9045 11747
rect 9306 11744 9312 11756
rect 9033 11716 9312 11744
rect 9033 11713 9045 11716
rect 8987 11707 9045 11713
rect 9306 11704 9312 11716
rect 9364 11704 9370 11756
rect 10152 11753 10180 11784
rect 10962 11772 10968 11824
rect 11020 11812 11026 11824
rect 12986 11812 12992 11824
rect 11020 11784 12992 11812
rect 11020 11772 11026 11784
rect 12986 11772 12992 11784
rect 13044 11812 13050 11824
rect 13924 11812 13952 11852
rect 14458 11840 14464 11852
rect 14516 11880 14522 11892
rect 15657 11883 15715 11889
rect 15657 11880 15669 11883
rect 14516 11852 15669 11880
rect 14516 11840 14522 11852
rect 15657 11849 15669 11852
rect 15703 11849 15715 11883
rect 15657 11843 15715 11849
rect 16850 11840 16856 11892
rect 16908 11840 16914 11892
rect 17221 11883 17279 11889
rect 17221 11849 17233 11883
rect 17267 11880 17279 11883
rect 18966 11880 18972 11892
rect 17267 11852 18972 11880
rect 17267 11849 17279 11852
rect 17221 11843 17279 11849
rect 18966 11840 18972 11852
rect 19024 11840 19030 11892
rect 19150 11840 19156 11892
rect 19208 11880 19214 11892
rect 25501 11883 25559 11889
rect 19208 11852 25452 11880
rect 19208 11840 19214 11852
rect 13044 11784 13952 11812
rect 13044 11772 13050 11784
rect 15194 11772 15200 11824
rect 15252 11772 15258 11824
rect 17402 11772 17408 11824
rect 17460 11812 17466 11824
rect 17770 11812 17776 11824
rect 17460 11784 17776 11812
rect 17460 11772 17466 11784
rect 17770 11772 17776 11784
rect 17828 11772 17834 11824
rect 18984 11812 19012 11840
rect 20990 11812 20996 11824
rect 18984 11784 20996 11812
rect 10045 11747 10103 11753
rect 10045 11744 10057 11747
rect 9784 11716 10057 11744
rect 7742 11676 7748 11688
rect 6656 11648 7748 11676
rect 7742 11636 7748 11648
rect 7800 11636 7806 11688
rect 8772 11676 8800 11704
rect 9582 11676 9588 11688
rect 8772 11648 9588 11676
rect 9582 11636 9588 11648
rect 9640 11636 9646 11688
rect 8846 11568 8852 11620
rect 8904 11608 8910 11620
rect 9784 11617 9812 11716
rect 10045 11713 10057 11716
rect 10091 11713 10103 11747
rect 10045 11707 10103 11713
rect 10138 11747 10196 11753
rect 10138 11713 10150 11747
rect 10184 11713 10196 11747
rect 10138 11707 10196 11713
rect 13078 11704 13084 11756
rect 13136 11704 13142 11756
rect 9858 11636 9864 11688
rect 9916 11676 9922 11688
rect 9953 11679 10011 11685
rect 9953 11676 9965 11679
rect 9916 11648 9965 11676
rect 9916 11636 9922 11648
rect 9953 11645 9965 11648
rect 9999 11645 10011 11679
rect 9953 11639 10011 11645
rect 10318 11636 10324 11688
rect 10376 11676 10382 11688
rect 10962 11676 10968 11688
rect 10376 11648 10968 11676
rect 10376 11636 10382 11648
rect 10962 11636 10968 11648
rect 11020 11636 11026 11688
rect 11882 11636 11888 11688
rect 11940 11676 11946 11688
rect 12250 11676 12256 11688
rect 11940 11648 12256 11676
rect 11940 11636 11946 11648
rect 12250 11636 12256 11648
rect 12308 11636 12314 11688
rect 12526 11636 12532 11688
rect 12584 11676 12590 11688
rect 13173 11679 13231 11685
rect 13173 11676 13185 11679
rect 12584 11648 13185 11676
rect 12584 11636 12590 11648
rect 13173 11645 13185 11648
rect 13219 11676 13231 11679
rect 13446 11676 13452 11688
rect 13219 11648 13452 11676
rect 13219 11645 13231 11648
rect 13173 11639 13231 11645
rect 13446 11636 13452 11648
rect 13504 11636 13510 11688
rect 13725 11679 13783 11685
rect 13725 11645 13737 11679
rect 13771 11676 13783 11679
rect 13906 11676 13912 11688
rect 13771 11648 13912 11676
rect 13771 11645 13783 11648
rect 13725 11639 13783 11645
rect 13906 11636 13912 11648
rect 13964 11636 13970 11688
rect 14108 11676 14136 11730
rect 15470 11704 15476 11756
rect 15528 11704 15534 11756
rect 15749 11747 15807 11753
rect 15749 11713 15761 11747
rect 15795 11713 15807 11747
rect 15749 11707 15807 11713
rect 15933 11747 15991 11753
rect 15933 11713 15945 11747
rect 15979 11744 15991 11747
rect 16114 11744 16120 11756
rect 15979 11716 16120 11744
rect 15979 11713 15991 11716
rect 15933 11707 15991 11713
rect 15764 11676 15792 11707
rect 16114 11704 16120 11716
rect 16172 11704 16178 11756
rect 17034 11704 17040 11756
rect 17092 11704 17098 11756
rect 17313 11747 17371 11753
rect 17313 11713 17325 11747
rect 17359 11744 17371 11747
rect 17678 11744 17684 11756
rect 17359 11716 17684 11744
rect 17359 11713 17371 11716
rect 17313 11707 17371 11713
rect 17678 11704 17684 11716
rect 17736 11744 17742 11756
rect 19518 11744 19524 11756
rect 17736 11716 19524 11744
rect 17736 11704 17742 11716
rect 19518 11704 19524 11716
rect 19576 11704 19582 11756
rect 20070 11704 20076 11756
rect 20128 11704 20134 11756
rect 20165 11747 20223 11753
rect 20165 11713 20177 11747
rect 20211 11744 20223 11747
rect 20254 11744 20260 11756
rect 20211 11716 20260 11744
rect 20211 11713 20223 11716
rect 20165 11707 20223 11713
rect 20254 11704 20260 11716
rect 20312 11704 20318 11756
rect 20548 11753 20576 11784
rect 20990 11772 20996 11784
rect 21048 11772 21054 11824
rect 22002 11772 22008 11824
rect 22060 11812 22066 11824
rect 24029 11815 24087 11821
rect 24029 11812 24041 11815
rect 22060 11784 24041 11812
rect 22060 11772 22066 11784
rect 24029 11781 24041 11784
rect 24075 11812 24087 11815
rect 24854 11812 24860 11824
rect 24075 11784 24860 11812
rect 24075 11781 24087 11784
rect 24029 11775 24087 11781
rect 24854 11772 24860 11784
rect 24912 11772 24918 11824
rect 25424 11812 25452 11852
rect 25501 11849 25513 11883
rect 25547 11880 25559 11883
rect 25590 11880 25596 11892
rect 25547 11852 25596 11880
rect 25547 11849 25559 11852
rect 25501 11843 25559 11849
rect 25590 11840 25596 11852
rect 25648 11840 25654 11892
rect 25682 11840 25688 11892
rect 25740 11880 25746 11892
rect 31202 11880 31208 11892
rect 25740 11852 31208 11880
rect 25740 11840 25746 11852
rect 31202 11840 31208 11852
rect 31260 11840 31266 11892
rect 33042 11840 33048 11892
rect 33100 11880 33106 11892
rect 33594 11880 33600 11892
rect 33100 11852 33600 11880
rect 33100 11840 33106 11852
rect 33594 11840 33600 11852
rect 33652 11880 33658 11892
rect 33652 11852 34718 11880
rect 33652 11840 33658 11852
rect 25869 11815 25927 11821
rect 25424 11784 25820 11812
rect 20349 11747 20407 11753
rect 20349 11713 20361 11747
rect 20395 11713 20407 11747
rect 20349 11707 20407 11713
rect 20533 11747 20591 11753
rect 20533 11713 20545 11747
rect 20579 11713 20591 11747
rect 20533 11707 20591 11713
rect 20809 11747 20867 11753
rect 20809 11713 20821 11747
rect 20855 11744 20867 11747
rect 20898 11744 20904 11756
rect 20855 11716 20904 11744
rect 20855 11713 20867 11716
rect 20809 11707 20867 11713
rect 18230 11676 18236 11688
rect 14108 11648 15700 11676
rect 15764 11648 18236 11676
rect 9769 11611 9827 11617
rect 9769 11608 9781 11611
rect 8904 11580 9781 11608
rect 8904 11568 8910 11580
rect 9769 11577 9781 11580
rect 9815 11577 9827 11611
rect 9769 11571 9827 11577
rect 9876 11580 10364 11608
rect 8662 11500 8668 11552
rect 8720 11540 8726 11552
rect 9125 11543 9183 11549
rect 9125 11540 9137 11543
rect 8720 11512 9137 11540
rect 8720 11500 8726 11512
rect 9125 11509 9137 11512
rect 9171 11509 9183 11543
rect 9125 11503 9183 11509
rect 9582 11500 9588 11552
rect 9640 11540 9646 11552
rect 9876 11540 9904 11580
rect 9640 11512 9904 11540
rect 9640 11500 9646 11512
rect 10042 11500 10048 11552
rect 10100 11540 10106 11552
rect 10229 11543 10287 11549
rect 10229 11540 10241 11543
rect 10100 11512 10241 11540
rect 10100 11500 10106 11512
rect 10229 11509 10241 11512
rect 10275 11509 10287 11543
rect 10336 11540 10364 11580
rect 12158 11568 12164 11620
rect 12216 11608 12222 11620
rect 12342 11608 12348 11620
rect 12216 11580 12348 11608
rect 12216 11568 12222 11580
rect 12342 11568 12348 11580
rect 12400 11608 12406 11620
rect 15672 11608 15700 11648
rect 18230 11636 18236 11648
rect 18288 11636 18294 11688
rect 20364 11676 20392 11707
rect 20898 11704 20904 11716
rect 20956 11704 20962 11756
rect 21085 11747 21143 11753
rect 21085 11713 21097 11747
rect 21131 11744 21143 11747
rect 21542 11744 21548 11756
rect 21131 11716 21548 11744
rect 21131 11713 21143 11716
rect 21085 11707 21143 11713
rect 21542 11704 21548 11716
rect 21600 11744 21606 11756
rect 22738 11744 22744 11756
rect 21600 11716 22744 11744
rect 21600 11704 21606 11716
rect 22738 11704 22744 11716
rect 22796 11744 22802 11756
rect 23382 11744 23388 11756
rect 22796 11716 23388 11744
rect 22796 11704 22802 11716
rect 23382 11704 23388 11716
rect 23440 11704 23446 11756
rect 24121 11747 24179 11753
rect 24121 11713 24133 11747
rect 24167 11744 24179 11747
rect 24210 11744 24216 11756
rect 24167 11716 24216 11744
rect 24167 11713 24179 11716
rect 24121 11707 24179 11713
rect 24210 11704 24216 11716
rect 24268 11704 24274 11756
rect 24486 11704 24492 11756
rect 24544 11704 24550 11756
rect 24946 11704 24952 11756
rect 25004 11704 25010 11756
rect 25130 11704 25136 11756
rect 25188 11704 25194 11756
rect 25225 11747 25283 11753
rect 25225 11713 25237 11747
rect 25271 11744 25283 11747
rect 25314 11744 25320 11756
rect 25271 11716 25320 11744
rect 25271 11713 25283 11716
rect 25225 11707 25283 11713
rect 25314 11704 25320 11716
rect 25372 11704 25378 11756
rect 25424 11744 25452 11784
rect 25501 11747 25559 11753
rect 25501 11744 25513 11747
rect 25424 11716 25513 11744
rect 25501 11713 25513 11716
rect 25547 11713 25559 11747
rect 25501 11707 25559 11713
rect 25685 11747 25743 11753
rect 25685 11713 25697 11747
rect 25731 11713 25743 11747
rect 25685 11707 25743 11713
rect 20180 11648 20392 11676
rect 20180 11620 20208 11648
rect 20714 11636 20720 11688
rect 20772 11676 20778 11688
rect 20993 11679 21051 11685
rect 20993 11676 21005 11679
rect 20772 11648 21005 11676
rect 20772 11636 20778 11648
rect 20993 11645 21005 11648
rect 21039 11676 21051 11679
rect 21266 11676 21272 11688
rect 21039 11648 21272 11676
rect 21039 11645 21051 11648
rect 20993 11639 21051 11645
rect 21266 11636 21272 11648
rect 21324 11636 21330 11688
rect 22094 11636 22100 11688
rect 22152 11676 22158 11688
rect 23198 11676 23204 11688
rect 22152 11648 23204 11676
rect 22152 11636 22158 11648
rect 23198 11636 23204 11648
rect 23256 11636 23262 11688
rect 24673 11679 24731 11685
rect 24673 11645 24685 11679
rect 24719 11645 24731 11679
rect 24673 11639 24731 11645
rect 16758 11608 16764 11620
rect 12400 11580 14228 11608
rect 15672 11580 16764 11608
rect 12400 11568 12406 11580
rect 12250 11540 12256 11552
rect 10336 11512 12256 11540
rect 10229 11503 10287 11509
rect 12250 11500 12256 11512
rect 12308 11500 12314 11552
rect 13446 11500 13452 11552
rect 13504 11500 13510 11552
rect 14200 11540 14228 11580
rect 16758 11568 16764 11580
rect 16816 11568 16822 11620
rect 17770 11568 17776 11620
rect 17828 11608 17834 11620
rect 19794 11608 19800 11620
rect 17828 11580 19800 11608
rect 17828 11568 17834 11580
rect 19794 11568 19800 11580
rect 19852 11568 19858 11620
rect 20162 11568 20168 11620
rect 20220 11568 20226 11620
rect 20257 11611 20315 11617
rect 20257 11577 20269 11611
rect 20303 11608 20315 11611
rect 20625 11611 20683 11617
rect 20625 11608 20637 11611
rect 20303 11580 20637 11608
rect 20303 11577 20315 11580
rect 20257 11571 20315 11577
rect 20625 11577 20637 11580
rect 20671 11577 20683 11611
rect 24688 11608 24716 11639
rect 25406 11636 25412 11688
rect 25464 11676 25470 11688
rect 25700 11676 25728 11707
rect 25464 11648 25728 11676
rect 25792 11676 25820 11784
rect 25869 11781 25881 11815
rect 25915 11812 25927 11815
rect 25958 11812 25964 11824
rect 25915 11784 25964 11812
rect 25915 11781 25927 11784
rect 25869 11775 25927 11781
rect 25958 11772 25964 11784
rect 26016 11772 26022 11824
rect 26053 11815 26111 11821
rect 26053 11781 26065 11815
rect 26099 11812 26111 11815
rect 26326 11812 26332 11824
rect 26099 11784 26332 11812
rect 26099 11781 26111 11784
rect 26053 11775 26111 11781
rect 26326 11772 26332 11784
rect 26384 11812 26390 11824
rect 30190 11812 30196 11824
rect 26384 11784 26740 11812
rect 26384 11772 26390 11784
rect 26145 11747 26203 11753
rect 26145 11713 26157 11747
rect 26191 11744 26203 11747
rect 26234 11744 26240 11756
rect 26191 11716 26240 11744
rect 26191 11713 26203 11716
rect 26145 11707 26203 11713
rect 26050 11676 26056 11688
rect 25792 11648 26056 11676
rect 25464 11636 25470 11648
rect 26050 11636 26056 11648
rect 26108 11636 26114 11688
rect 25041 11611 25099 11617
rect 25041 11608 25053 11611
rect 24688 11580 25053 11608
rect 20625 11571 20683 11577
rect 25041 11577 25053 11580
rect 25087 11608 25099 11611
rect 25222 11608 25228 11620
rect 25087 11580 25228 11608
rect 25087 11577 25099 11580
rect 25041 11571 25099 11577
rect 25222 11568 25228 11580
rect 25280 11608 25286 11620
rect 25682 11608 25688 11620
rect 25280 11580 25688 11608
rect 25280 11568 25286 11580
rect 25682 11568 25688 11580
rect 25740 11568 25746 11620
rect 25958 11568 25964 11620
rect 26016 11608 26022 11620
rect 26160 11608 26188 11707
rect 26234 11704 26240 11716
rect 26292 11704 26298 11756
rect 26418 11704 26424 11756
rect 26476 11704 26482 11756
rect 26712 11753 26740 11784
rect 27816 11784 30196 11812
rect 26605 11747 26663 11753
rect 26605 11713 26617 11747
rect 26651 11713 26663 11747
rect 26605 11707 26663 11713
rect 26697 11747 26755 11753
rect 26697 11713 26709 11747
rect 26743 11713 26755 11747
rect 26697 11707 26755 11713
rect 26620 11676 26648 11707
rect 27816 11676 27844 11784
rect 30190 11772 30196 11784
rect 30248 11772 30254 11824
rect 33321 11815 33379 11821
rect 33321 11781 33333 11815
rect 33367 11812 33379 11815
rect 33502 11812 33508 11824
rect 33367 11784 33508 11812
rect 33367 11781 33379 11784
rect 33321 11775 33379 11781
rect 33502 11772 33508 11784
rect 33560 11772 33566 11824
rect 34690 11821 34718 11852
rect 34790 11840 34796 11892
rect 34848 11880 34854 11892
rect 35066 11880 35072 11892
rect 34848 11852 35072 11880
rect 34848 11840 34854 11852
rect 35066 11840 35072 11852
rect 35124 11840 35130 11892
rect 37093 11883 37151 11889
rect 37093 11849 37105 11883
rect 37139 11880 37151 11883
rect 38102 11880 38108 11892
rect 37139 11852 38108 11880
rect 37139 11849 37151 11852
rect 37093 11843 37151 11849
rect 38102 11840 38108 11852
rect 38160 11840 38166 11892
rect 38473 11883 38531 11889
rect 38473 11849 38485 11883
rect 38519 11880 38531 11883
rect 38519 11852 39068 11880
rect 38519 11849 38531 11852
rect 38473 11843 38531 11849
rect 34675 11815 34733 11821
rect 34675 11781 34687 11815
rect 34721 11781 34733 11815
rect 34675 11775 34733 11781
rect 34882 11772 34888 11824
rect 34940 11772 34946 11824
rect 39040 11821 39068 11852
rect 39025 11815 39083 11821
rect 39025 11781 39037 11815
rect 39071 11781 39083 11815
rect 39025 11775 39083 11781
rect 27982 11704 27988 11756
rect 28040 11744 28046 11756
rect 28442 11744 28448 11756
rect 28040 11716 28448 11744
rect 28040 11704 28046 11716
rect 28442 11704 28448 11716
rect 28500 11744 28506 11756
rect 28629 11747 28687 11753
rect 28629 11744 28641 11747
rect 28500 11716 28641 11744
rect 28500 11704 28506 11716
rect 28629 11713 28641 11716
rect 28675 11713 28687 11747
rect 28629 11707 28687 11713
rect 29454 11704 29460 11756
rect 29512 11744 29518 11756
rect 30098 11744 30104 11756
rect 29512 11716 30104 11744
rect 29512 11704 29518 11716
rect 30098 11704 30104 11716
rect 30156 11704 30162 11756
rect 32493 11747 32551 11753
rect 32493 11713 32505 11747
rect 32539 11744 32551 11747
rect 32858 11744 32864 11756
rect 32539 11716 32864 11744
rect 32539 11713 32551 11716
rect 32493 11707 32551 11713
rect 32858 11704 32864 11716
rect 32916 11704 32922 11756
rect 33594 11704 33600 11756
rect 33652 11704 33658 11756
rect 34054 11704 34060 11756
rect 34112 11744 34118 11756
rect 34793 11747 34851 11753
rect 34793 11744 34805 11747
rect 34112 11716 34805 11744
rect 34112 11704 34118 11716
rect 34793 11713 34805 11716
rect 34839 11713 34851 11747
rect 34793 11707 34851 11713
rect 34977 11747 35035 11753
rect 34977 11713 34989 11747
rect 35023 11744 35035 11747
rect 35342 11744 35348 11756
rect 35023 11716 35348 11744
rect 35023 11713 35035 11716
rect 34977 11707 35035 11713
rect 35342 11704 35348 11716
rect 35400 11704 35406 11756
rect 36262 11704 36268 11756
rect 36320 11744 36326 11756
rect 36449 11747 36507 11753
rect 36449 11744 36461 11747
rect 36320 11716 36461 11744
rect 36320 11704 36326 11716
rect 36449 11713 36461 11716
rect 36495 11713 36507 11747
rect 36449 11707 36507 11713
rect 36538 11704 36544 11756
rect 36596 11704 36602 11756
rect 36630 11704 36636 11756
rect 36688 11744 36694 11756
rect 36725 11747 36783 11753
rect 36725 11744 36737 11747
rect 36688 11716 36737 11744
rect 36688 11704 36694 11716
rect 36725 11713 36737 11716
rect 36771 11713 36783 11747
rect 36725 11707 36783 11713
rect 36814 11704 36820 11756
rect 36872 11704 36878 11756
rect 36914 11747 36972 11753
rect 36914 11713 36926 11747
rect 36960 11713 36972 11747
rect 36914 11707 36972 11713
rect 26620 11648 27844 11676
rect 28537 11679 28595 11685
rect 28537 11645 28549 11679
rect 28583 11676 28595 11679
rect 29546 11676 29552 11688
rect 28583 11648 29552 11676
rect 28583 11645 28595 11648
rect 28537 11639 28595 11645
rect 29546 11636 29552 11648
rect 29604 11636 29610 11688
rect 30558 11636 30564 11688
rect 30616 11676 30622 11688
rect 31665 11679 31723 11685
rect 31665 11676 31677 11679
rect 30616 11648 31677 11676
rect 30616 11636 30622 11648
rect 31665 11645 31677 11648
rect 31711 11676 31723 11679
rect 31846 11676 31852 11688
rect 31711 11648 31852 11676
rect 31711 11645 31723 11648
rect 31665 11639 31723 11645
rect 31846 11636 31852 11648
rect 31904 11636 31910 11688
rect 31941 11679 31999 11685
rect 31941 11645 31953 11679
rect 31987 11676 31999 11679
rect 33502 11676 33508 11688
rect 31987 11648 33508 11676
rect 31987 11645 31999 11648
rect 31941 11639 31999 11645
rect 33502 11636 33508 11648
rect 33560 11636 33566 11688
rect 34517 11679 34575 11685
rect 34517 11645 34529 11679
rect 34563 11645 34575 11679
rect 35360 11676 35388 11704
rect 36929 11676 36957 11707
rect 38010 11704 38016 11756
rect 38068 11704 38074 11756
rect 38286 11704 38292 11756
rect 38344 11704 38350 11756
rect 38746 11704 38752 11756
rect 38804 11704 38810 11756
rect 35360 11648 36957 11676
rect 34517 11639 34575 11645
rect 26016 11580 26188 11608
rect 26421 11611 26479 11617
rect 26016 11568 26022 11580
rect 26421 11577 26433 11611
rect 26467 11608 26479 11611
rect 26510 11608 26516 11620
rect 26467 11580 26516 11608
rect 26467 11577 26479 11580
rect 26421 11571 26479 11577
rect 26510 11568 26516 11580
rect 26568 11568 26574 11620
rect 26878 11568 26884 11620
rect 26936 11608 26942 11620
rect 28261 11611 28319 11617
rect 28261 11608 28273 11611
rect 26936 11580 28273 11608
rect 26936 11568 26942 11580
rect 28261 11577 28273 11580
rect 28307 11577 28319 11611
rect 28261 11571 28319 11577
rect 19889 11543 19947 11549
rect 19889 11540 19901 11543
rect 14200 11512 19901 11540
rect 19889 11509 19901 11512
rect 19935 11509 19947 11543
rect 19889 11503 19947 11509
rect 20070 11500 20076 11552
rect 20128 11540 20134 11552
rect 20438 11540 20444 11552
rect 20128 11512 20444 11540
rect 20128 11500 20134 11512
rect 20438 11500 20444 11512
rect 20496 11500 20502 11552
rect 21358 11500 21364 11552
rect 21416 11540 21422 11552
rect 24213 11543 24271 11549
rect 24213 11540 24225 11543
rect 21416 11512 24225 11540
rect 21416 11500 21422 11512
rect 24213 11509 24225 11512
rect 24259 11509 24271 11543
rect 24213 11503 24271 11509
rect 24762 11500 24768 11552
rect 24820 11500 24826 11552
rect 24946 11500 24952 11552
rect 25004 11540 25010 11552
rect 25866 11540 25872 11552
rect 25004 11512 25872 11540
rect 25004 11500 25010 11512
rect 25866 11500 25872 11512
rect 25924 11500 25930 11552
rect 26234 11500 26240 11552
rect 26292 11540 26298 11552
rect 27614 11540 27620 11552
rect 26292 11512 27620 11540
rect 26292 11500 26298 11512
rect 27614 11500 27620 11512
rect 27672 11500 27678 11552
rect 28350 11500 28356 11552
rect 28408 11540 28414 11552
rect 28626 11540 28632 11552
rect 28408 11512 28632 11540
rect 28408 11500 28414 11512
rect 28626 11500 28632 11512
rect 28684 11500 28690 11552
rect 31938 11500 31944 11552
rect 31996 11540 32002 11552
rect 33410 11540 33416 11552
rect 31996 11512 33416 11540
rect 31996 11500 32002 11512
rect 33410 11500 33416 11512
rect 33468 11540 33474 11552
rect 33689 11543 33747 11549
rect 33689 11540 33701 11543
rect 33468 11512 33701 11540
rect 33468 11500 33474 11512
rect 33689 11509 33701 11512
rect 33735 11509 33747 11543
rect 34532 11540 34560 11639
rect 37366 11636 37372 11688
rect 37424 11676 37430 11688
rect 38105 11679 38163 11685
rect 38105 11676 38117 11679
rect 37424 11648 38117 11676
rect 37424 11636 37430 11648
rect 38105 11645 38117 11648
rect 38151 11645 38163 11679
rect 38105 11639 38163 11645
rect 38930 11636 38936 11688
rect 38988 11636 38994 11688
rect 34606 11540 34612 11552
rect 34532 11512 34612 11540
rect 33689 11503 33747 11509
rect 34606 11500 34612 11512
rect 34664 11500 34670 11552
rect 35161 11543 35219 11549
rect 35161 11509 35173 11543
rect 35207 11540 35219 11543
rect 38013 11543 38071 11549
rect 38013 11540 38025 11543
rect 35207 11512 38025 11540
rect 35207 11509 35219 11512
rect 35161 11503 35219 11509
rect 38013 11509 38025 11512
rect 38059 11540 38071 11543
rect 38378 11540 38384 11552
rect 38059 11512 38384 11540
rect 38059 11509 38071 11512
rect 38013 11503 38071 11509
rect 38378 11500 38384 11512
rect 38436 11500 38442 11552
rect 38562 11500 38568 11552
rect 38620 11500 38626 11552
rect 39025 11543 39083 11549
rect 39025 11509 39037 11543
rect 39071 11540 39083 11543
rect 39298 11540 39304 11552
rect 39071 11512 39304 11540
rect 39071 11509 39083 11512
rect 39025 11503 39083 11509
rect 39298 11500 39304 11512
rect 39356 11500 39362 11552
rect 1104 11450 40572 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 40572 11450
rect 1104 11376 40572 11398
rect 8662 11296 8668 11348
rect 8720 11296 8726 11348
rect 9306 11296 9312 11348
rect 9364 11336 9370 11348
rect 12158 11336 12164 11348
rect 9364 11308 12164 11336
rect 9364 11296 9370 11308
rect 7098 11228 7104 11280
rect 7156 11268 7162 11280
rect 8113 11271 8171 11277
rect 8113 11268 8125 11271
rect 7156 11240 8125 11268
rect 7156 11228 7162 11240
rect 8113 11237 8125 11240
rect 8159 11237 8171 11271
rect 8113 11231 8171 11237
rect 10229 11271 10287 11277
rect 10229 11237 10241 11271
rect 10275 11237 10287 11271
rect 10229 11231 10287 11237
rect 8757 11203 8815 11209
rect 8757 11169 8769 11203
rect 8803 11200 8815 11203
rect 9033 11203 9091 11209
rect 9033 11200 9045 11203
rect 8803 11172 9045 11200
rect 8803 11169 8815 11172
rect 8757 11163 8815 11169
rect 9033 11169 9045 11172
rect 9079 11169 9091 11203
rect 9033 11163 9091 11169
rect 9582 11160 9588 11212
rect 9640 11200 9646 11212
rect 9640 11172 9812 11200
rect 9640 11160 9646 11172
rect 2041 11135 2099 11141
rect 2041 11101 2053 11135
rect 2087 11132 2099 11135
rect 3510 11132 3516 11144
rect 2087 11104 3516 11132
rect 2087 11101 2099 11104
rect 2041 11095 2099 11101
rect 3510 11092 3516 11104
rect 3568 11092 3574 11144
rect 7650 11092 7656 11144
rect 7708 11132 7714 11144
rect 7837 11135 7895 11141
rect 7837 11132 7849 11135
rect 7708 11104 7849 11132
rect 7708 11092 7714 11104
rect 7837 11101 7849 11104
rect 7883 11101 7895 11135
rect 7837 11095 7895 11101
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11132 8079 11135
rect 8294 11135 8352 11141
rect 8294 11132 8306 11135
rect 8067 11104 8306 11132
rect 8067 11101 8079 11104
rect 8021 11095 8079 11101
rect 8294 11101 8306 11104
rect 8340 11132 8352 11135
rect 8386 11132 8392 11144
rect 8340 11104 8392 11132
rect 8340 11101 8352 11104
rect 8294 11095 8352 11101
rect 8386 11092 8392 11104
rect 8444 11092 8450 11144
rect 8941 11135 8999 11141
rect 8941 11101 8953 11135
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11132 9183 11135
rect 9306 11132 9312 11144
rect 9171 11104 9312 11132
rect 9171 11101 9183 11104
rect 9125 11095 9183 11101
rect 7926 11024 7932 11076
rect 7984 11064 7990 11076
rect 8202 11064 8208 11076
rect 7984 11036 8208 11064
rect 7984 11024 7990 11036
rect 8202 11024 8208 11036
rect 8260 11064 8266 11076
rect 8956 11064 8984 11095
rect 9306 11092 9312 11104
rect 9364 11092 9370 11144
rect 9490 11092 9496 11144
rect 9548 11132 9554 11144
rect 9784 11141 9812 11172
rect 9769 11135 9827 11141
rect 9548 11104 9720 11132
rect 9548 11092 9554 11104
rect 8260 11036 8984 11064
rect 8260 11024 8266 11036
rect 9398 11024 9404 11076
rect 9456 11064 9462 11076
rect 9585 11067 9643 11073
rect 9585 11064 9597 11067
rect 9456 11036 9597 11064
rect 9456 11024 9462 11036
rect 9585 11033 9597 11036
rect 9631 11033 9643 11067
rect 9692 11064 9720 11104
rect 9769 11101 9781 11135
rect 9815 11101 9827 11135
rect 9769 11095 9827 11101
rect 9861 11135 9919 11141
rect 9861 11101 9873 11135
rect 9907 11132 9919 11135
rect 9950 11132 9956 11144
rect 9907 11104 9956 11132
rect 9907 11101 9919 11104
rect 9861 11095 9919 11101
rect 9950 11092 9956 11104
rect 10008 11092 10014 11144
rect 10042 11092 10048 11144
rect 10100 11092 10106 11144
rect 10137 11135 10195 11141
rect 10137 11101 10149 11135
rect 10183 11132 10195 11135
rect 10244 11132 10272 11231
rect 10183 11104 10272 11132
rect 10336 11132 10364 11308
rect 12158 11296 12164 11308
rect 12216 11296 12222 11348
rect 12342 11296 12348 11348
rect 12400 11336 12406 11348
rect 13814 11336 13820 11348
rect 12400 11308 13820 11336
rect 12400 11296 12406 11308
rect 11701 11271 11759 11277
rect 11701 11237 11713 11271
rect 11747 11268 11759 11271
rect 11747 11240 12112 11268
rect 11747 11237 11759 11240
rect 11701 11231 11759 11237
rect 11057 11203 11115 11209
rect 11057 11200 11069 11203
rect 10520 11172 11069 11200
rect 10520 11141 10548 11172
rect 11057 11169 11069 11172
rect 11103 11169 11115 11203
rect 11057 11163 11115 11169
rect 11348 11172 11836 11200
rect 10408 11135 10466 11141
rect 10408 11132 10420 11135
rect 10336 11104 10420 11132
rect 10183 11101 10195 11104
rect 10137 11095 10195 11101
rect 10408 11101 10420 11104
rect 10454 11101 10466 11135
rect 10408 11095 10466 11101
rect 10505 11135 10563 11141
rect 10505 11101 10517 11135
rect 10551 11101 10563 11135
rect 10725 11135 10783 11141
rect 10725 11132 10737 11135
rect 10505 11095 10563 11101
rect 10704 11101 10737 11132
rect 10771 11101 10783 11135
rect 10704 11095 10783 11101
rect 10318 11064 10324 11076
rect 9692 11036 10324 11064
rect 9585 11027 9643 11033
rect 10318 11024 10324 11036
rect 10376 11064 10382 11076
rect 10597 11067 10655 11073
rect 10597 11064 10609 11067
rect 10376 11036 10609 11064
rect 10376 11024 10382 11036
rect 10597 11033 10609 11036
rect 10643 11033 10655 11067
rect 10597 11027 10655 11033
rect 10704 11008 10732 11095
rect 10870 11092 10876 11144
rect 10928 11092 10934 11144
rect 11146 11092 11152 11144
rect 11204 11132 11210 11144
rect 11348 11141 11376 11172
rect 11333 11135 11391 11141
rect 11333 11132 11345 11135
rect 11204 11104 11345 11132
rect 11204 11092 11210 11104
rect 11333 11101 11345 11104
rect 11379 11101 11391 11135
rect 11333 11095 11391 11101
rect 11422 11092 11428 11144
rect 11480 11132 11486 11144
rect 11808 11141 11836 11172
rect 11517 11135 11575 11141
rect 11517 11132 11529 11135
rect 11480 11104 11529 11132
rect 11480 11092 11486 11104
rect 11517 11101 11529 11104
rect 11563 11101 11575 11135
rect 11517 11095 11575 11101
rect 11793 11135 11851 11141
rect 11793 11101 11805 11135
rect 11839 11101 11851 11135
rect 11793 11095 11851 11101
rect 11977 11135 12035 11141
rect 11977 11101 11989 11135
rect 12023 11101 12035 11135
rect 11977 11095 12035 11101
rect 11532 11064 11560 11095
rect 11992 11064 12020 11095
rect 11532 11036 12020 11064
rect 12084 11064 12112 11240
rect 12176 11132 12204 11296
rect 12253 11271 12311 11277
rect 12253 11237 12265 11271
rect 12299 11268 12311 11271
rect 12434 11268 12440 11280
rect 12299 11240 12440 11268
rect 12299 11237 12311 11240
rect 12253 11231 12311 11237
rect 12434 11228 12440 11240
rect 12492 11228 12498 11280
rect 12391 11135 12449 11141
rect 12391 11132 12403 11135
rect 12176 11104 12403 11132
rect 12391 11101 12403 11104
rect 12437 11101 12449 11135
rect 12391 11095 12449 11101
rect 12526 11092 12532 11144
rect 12584 11092 12590 11144
rect 12636 11141 12664 11308
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 14185 11339 14243 11345
rect 14185 11305 14197 11339
rect 14231 11336 14243 11339
rect 15102 11336 15108 11348
rect 14231 11308 15108 11336
rect 14231 11305 14243 11308
rect 14185 11299 14243 11305
rect 15102 11296 15108 11308
rect 15160 11296 15166 11348
rect 17310 11296 17316 11348
rect 17368 11296 17374 11348
rect 17589 11339 17647 11345
rect 17589 11305 17601 11339
rect 17635 11336 17647 11339
rect 17862 11336 17868 11348
rect 17635 11308 17868 11336
rect 17635 11305 17647 11308
rect 17589 11299 17647 11305
rect 17862 11296 17868 11308
rect 17920 11296 17926 11348
rect 18230 11296 18236 11348
rect 18288 11296 18294 11348
rect 19242 11296 19248 11348
rect 19300 11336 19306 11348
rect 19889 11339 19947 11345
rect 19889 11336 19901 11339
rect 19300 11308 19901 11336
rect 19300 11296 19306 11308
rect 19889 11305 19901 11308
rect 19935 11336 19947 11339
rect 20990 11336 20996 11348
rect 19935 11308 20996 11336
rect 19935 11305 19947 11308
rect 19889 11299 19947 11305
rect 20990 11296 20996 11308
rect 21048 11296 21054 11348
rect 21082 11296 21088 11348
rect 21140 11336 21146 11348
rect 21266 11336 21272 11348
rect 21140 11308 21272 11336
rect 21140 11296 21146 11308
rect 21266 11296 21272 11308
rect 21324 11296 21330 11348
rect 21729 11339 21787 11345
rect 21729 11305 21741 11339
rect 21775 11336 21787 11339
rect 22186 11336 22192 11348
rect 21775 11308 22192 11336
rect 21775 11305 21787 11308
rect 21729 11299 21787 11305
rect 22186 11296 22192 11308
rect 22244 11336 22250 11348
rect 22462 11336 22468 11348
rect 22244 11308 22468 11336
rect 22244 11296 22250 11308
rect 22462 11296 22468 11308
rect 22520 11296 22526 11348
rect 24394 11296 24400 11348
rect 24452 11296 24458 11348
rect 24581 11339 24639 11345
rect 24581 11305 24593 11339
rect 24627 11336 24639 11339
rect 24762 11336 24768 11348
rect 24627 11308 24768 11336
rect 24627 11305 24639 11308
rect 24581 11299 24639 11305
rect 12802 11228 12808 11280
rect 12860 11268 12866 11280
rect 17129 11271 17187 11277
rect 17129 11268 17141 11271
rect 12860 11240 17141 11268
rect 12860 11228 12866 11240
rect 13004 11200 13032 11240
rect 17129 11237 17141 11240
rect 17175 11237 17187 11271
rect 17129 11231 17187 11237
rect 20073 11271 20131 11277
rect 20073 11237 20085 11271
rect 20119 11237 20131 11271
rect 20530 11268 20536 11280
rect 20073 11231 20131 11237
rect 20272 11240 20536 11268
rect 12912 11172 13032 11200
rect 12912 11141 12940 11172
rect 15194 11160 15200 11212
rect 15252 11200 15258 11212
rect 15473 11203 15531 11209
rect 15473 11200 15485 11203
rect 15252 11172 15485 11200
rect 15252 11160 15258 11172
rect 15473 11169 15485 11172
rect 15519 11200 15531 11203
rect 16114 11200 16120 11212
rect 15519 11172 16120 11200
rect 15519 11169 15531 11172
rect 15473 11163 15531 11169
rect 16114 11160 16120 11172
rect 16172 11160 16178 11212
rect 17586 11160 17592 11212
rect 17644 11200 17650 11212
rect 20088 11200 20116 11231
rect 20272 11209 20300 11240
rect 20530 11228 20536 11240
rect 20588 11268 20594 11280
rect 24596 11268 24624 11299
rect 24762 11296 24768 11308
rect 24820 11296 24826 11348
rect 26050 11296 26056 11348
rect 26108 11336 26114 11348
rect 26786 11336 26792 11348
rect 26108 11308 26792 11336
rect 26108 11296 26114 11308
rect 26786 11296 26792 11308
rect 26844 11296 26850 11348
rect 27065 11339 27123 11345
rect 27065 11305 27077 11339
rect 27111 11336 27123 11339
rect 27982 11336 27988 11348
rect 27111 11308 27988 11336
rect 27111 11305 27123 11308
rect 27065 11299 27123 11305
rect 27982 11296 27988 11308
rect 28040 11296 28046 11348
rect 28077 11339 28135 11345
rect 28077 11305 28089 11339
rect 28123 11336 28135 11339
rect 28258 11336 28264 11348
rect 28123 11308 28264 11336
rect 28123 11305 28135 11308
rect 28077 11299 28135 11305
rect 28258 11296 28264 11308
rect 28316 11336 28322 11348
rect 28445 11339 28503 11345
rect 28445 11336 28457 11339
rect 28316 11308 28457 11336
rect 28316 11296 28322 11308
rect 28445 11305 28457 11308
rect 28491 11305 28503 11339
rect 28445 11299 28503 11305
rect 29546 11296 29552 11348
rect 29604 11336 29610 11348
rect 30926 11336 30932 11348
rect 29604 11308 30932 11336
rect 29604 11296 29610 11308
rect 30926 11296 30932 11308
rect 30984 11296 30990 11348
rect 37185 11339 37243 11345
rect 37185 11305 37197 11339
rect 37231 11336 37243 11339
rect 37274 11336 37280 11348
rect 37231 11308 37280 11336
rect 37231 11305 37243 11308
rect 37185 11299 37243 11305
rect 37274 11296 37280 11308
rect 37332 11296 37338 11348
rect 20588 11240 21864 11268
rect 20588 11228 20594 11240
rect 17644 11172 20116 11200
rect 20257 11203 20315 11209
rect 17644 11160 17650 11172
rect 12621 11135 12679 11141
rect 12621 11101 12633 11135
rect 12667 11101 12679 11135
rect 12621 11095 12679 11101
rect 12804 11135 12862 11141
rect 12804 11101 12816 11135
rect 12850 11101 12862 11135
rect 12804 11095 12862 11101
rect 12897 11135 12955 11141
rect 12897 11101 12909 11135
rect 12943 11101 12955 11135
rect 12897 11095 12955 11101
rect 12989 11135 13047 11141
rect 12989 11101 13001 11135
rect 13035 11132 13047 11135
rect 13035 11104 13216 11132
rect 13035 11101 13047 11104
rect 12989 11095 13047 11101
rect 12250 11064 12256 11076
rect 12084 11036 12256 11064
rect 12250 11024 12256 11036
rect 12308 11064 12314 11076
rect 12820 11064 12848 11095
rect 13081 11067 13139 11073
rect 13081 11064 13093 11067
rect 12308 11036 12756 11064
rect 12820 11036 13093 11064
rect 12308 11024 12314 11036
rect 1854 10956 1860 11008
rect 1912 10956 1918 11008
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 9490 10996 9496 11008
rect 8352 10968 9496 10996
rect 8352 10956 8358 10968
rect 9490 10956 9496 10968
rect 9548 10956 9554 11008
rect 9766 10956 9772 11008
rect 9824 10996 9830 11008
rect 10686 10996 10692 11008
rect 9824 10968 10692 10996
rect 9824 10956 9830 10968
rect 10686 10956 10692 10968
rect 10744 10956 10750 11008
rect 11885 10999 11943 11005
rect 11885 10965 11897 10999
rect 11931 10996 11943 10999
rect 12342 10996 12348 11008
rect 11931 10968 12348 10996
rect 11931 10965 11943 10968
rect 11885 10959 11943 10965
rect 12342 10956 12348 10968
rect 12400 10956 12406 11008
rect 12728 10996 12756 11036
rect 13081 11033 13093 11036
rect 13127 11033 13139 11067
rect 13081 11027 13139 11033
rect 13188 10996 13216 11104
rect 13446 11092 13452 11144
rect 13504 11132 13510 11144
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13504 11104 14105 11132
rect 13504 11092 13510 11104
rect 14093 11101 14105 11104
rect 14139 11101 14151 11135
rect 14093 11095 14151 11101
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11132 14335 11135
rect 14366 11132 14372 11144
rect 14323 11104 14372 11132
rect 14323 11101 14335 11104
rect 14277 11095 14335 11101
rect 14366 11092 14372 11104
rect 14424 11092 14430 11144
rect 15657 11135 15715 11141
rect 15657 11101 15669 11135
rect 15703 11132 15715 11135
rect 16574 11132 16580 11144
rect 15703 11104 16580 11132
rect 15703 11101 15715 11104
rect 15657 11095 15715 11101
rect 16574 11092 16580 11104
rect 16632 11132 16638 11144
rect 16942 11132 16948 11144
rect 16632 11104 16948 11132
rect 16632 11092 16638 11104
rect 16942 11092 16948 11104
rect 17000 11092 17006 11144
rect 17770 11132 17776 11144
rect 17420 11104 17776 11132
rect 17297 11067 17355 11073
rect 17297 11033 17309 11067
rect 17343 11064 17355 11067
rect 17420 11064 17448 11104
rect 17770 11092 17776 11104
rect 17828 11092 17834 11144
rect 18064 11141 18092 11172
rect 20257 11169 20269 11203
rect 20303 11169 20315 11203
rect 20257 11163 20315 11169
rect 20346 11160 20352 11212
rect 20404 11160 20410 11212
rect 20806 11160 20812 11212
rect 20864 11200 20870 11212
rect 20864 11172 21772 11200
rect 20864 11160 20870 11172
rect 17865 11135 17923 11141
rect 17865 11101 17877 11135
rect 17911 11101 17923 11135
rect 17865 11095 17923 11101
rect 18049 11135 18107 11141
rect 18049 11101 18061 11135
rect 18095 11101 18107 11135
rect 18049 11095 18107 11101
rect 18141 11135 18199 11141
rect 18141 11101 18153 11135
rect 18187 11132 18199 11135
rect 18233 11135 18291 11141
rect 18233 11132 18245 11135
rect 18187 11104 18245 11132
rect 18187 11101 18199 11104
rect 18141 11095 18199 11101
rect 18233 11101 18245 11104
rect 18279 11101 18291 11135
rect 18233 11095 18291 11101
rect 17343 11036 17448 11064
rect 17497 11067 17555 11073
rect 17343 11033 17355 11036
rect 17297 11027 17355 11033
rect 17497 11033 17509 11067
rect 17543 11064 17555 11067
rect 17880 11064 17908 11095
rect 18248 11064 18276 11095
rect 18506 11092 18512 11144
rect 18564 11092 18570 11144
rect 21744 11141 21772 11172
rect 20533 11135 20591 11141
rect 20533 11101 20545 11135
rect 20579 11101 20591 11135
rect 20533 11095 20591 11101
rect 20717 11135 20775 11141
rect 20717 11101 20729 11135
rect 20763 11132 20775 11135
rect 21545 11135 21603 11141
rect 21545 11132 21557 11135
rect 20763 11104 21557 11132
rect 20763 11101 20775 11104
rect 20717 11095 20775 11101
rect 21545 11101 21557 11104
rect 21591 11101 21603 11135
rect 21545 11095 21603 11101
rect 21729 11135 21787 11141
rect 21729 11101 21741 11135
rect 21775 11101 21787 11135
rect 21729 11095 21787 11101
rect 19334 11064 19340 11076
rect 17543 11036 18184 11064
rect 18248 11036 19340 11064
rect 17543 11033 17555 11036
rect 17497 11027 17555 11033
rect 12728 10968 13216 10996
rect 17402 10956 17408 11008
rect 17460 10996 17466 11008
rect 17512 10996 17540 11027
rect 17460 10968 17540 10996
rect 18156 10996 18184 11036
rect 19334 11024 19340 11036
rect 19392 11024 19398 11076
rect 19702 11064 19708 11076
rect 19444 11036 19708 11064
rect 18417 10999 18475 11005
rect 18417 10996 18429 10999
rect 18156 10968 18429 10996
rect 17460 10956 17466 10968
rect 18417 10965 18429 10968
rect 18463 10996 18475 10999
rect 19444 10996 19472 11036
rect 19702 11024 19708 11036
rect 19760 11024 19766 11076
rect 19921 11067 19979 11073
rect 19921 11033 19933 11067
rect 19967 11064 19979 11067
rect 20254 11064 20260 11076
rect 19967 11036 20260 11064
rect 19967 11033 19979 11036
rect 19921 11027 19979 11033
rect 20254 11024 20260 11036
rect 20312 11024 20318 11076
rect 18463 10968 19472 10996
rect 20548 10996 20576 11095
rect 21269 11067 21327 11073
rect 21269 11033 21281 11067
rect 21315 11064 21327 11067
rect 21450 11064 21456 11076
rect 21315 11036 21456 11064
rect 21315 11033 21327 11036
rect 21269 11027 21327 11033
rect 21450 11024 21456 11036
rect 21508 11024 21514 11076
rect 21836 11064 21864 11240
rect 22664 11240 24624 11268
rect 22278 11160 22284 11212
rect 22336 11160 22342 11212
rect 22462 11092 22468 11144
rect 22520 11092 22526 11144
rect 22664 11141 22692 11240
rect 25406 11228 25412 11280
rect 25464 11268 25470 11280
rect 25464 11240 28488 11268
rect 25464 11228 25470 11240
rect 28000 11212 28028 11240
rect 24673 11203 24731 11209
rect 24673 11200 24685 11203
rect 22940 11172 24685 11200
rect 22940 11141 22968 11172
rect 24673 11169 24685 11172
rect 24719 11200 24731 11203
rect 27525 11203 27583 11209
rect 27525 11200 27537 11203
rect 24719 11172 27537 11200
rect 24719 11169 24731 11172
rect 24673 11163 24731 11169
rect 27525 11169 27537 11172
rect 27571 11169 27583 11203
rect 27525 11163 27583 11169
rect 27982 11160 27988 11212
rect 28040 11160 28046 11212
rect 28460 11200 28488 11240
rect 33244 11240 33640 11268
rect 30190 11200 30196 11212
rect 28460 11172 29040 11200
rect 22649 11135 22707 11141
rect 22649 11101 22661 11135
rect 22695 11101 22707 11135
rect 22649 11095 22707 11101
rect 22925 11135 22983 11141
rect 22925 11101 22937 11135
rect 22971 11101 22983 11135
rect 22925 11095 22983 11101
rect 23198 11092 23204 11144
rect 23256 11092 23262 11144
rect 24762 11092 24768 11144
rect 24820 11092 24826 11144
rect 25130 11092 25136 11144
rect 25188 11132 25194 11144
rect 25869 11135 25927 11141
rect 25869 11132 25881 11135
rect 25188 11104 25881 11132
rect 25188 11092 25194 11104
rect 25869 11101 25881 11104
rect 25915 11101 25927 11135
rect 25869 11095 25927 11101
rect 26145 11135 26203 11141
rect 26145 11101 26157 11135
rect 26191 11132 26203 11135
rect 26326 11132 26332 11144
rect 26191 11104 26332 11132
rect 26191 11101 26203 11104
rect 26145 11095 26203 11101
rect 25884 11064 25912 11095
rect 26326 11092 26332 11104
rect 26384 11092 26390 11144
rect 26786 11092 26792 11144
rect 26844 11092 26850 11144
rect 26881 11135 26939 11141
rect 26881 11101 26893 11135
rect 26927 11132 26939 11135
rect 26970 11132 26976 11144
rect 26927 11104 26976 11132
rect 26927 11101 26939 11104
rect 26881 11095 26939 11101
rect 26970 11092 26976 11104
rect 27028 11132 27034 11144
rect 27028 11104 27644 11132
rect 27028 11092 27034 11104
rect 26418 11064 26424 11076
rect 21836 11036 23060 11064
rect 25884 11036 26424 11064
rect 23032 11008 23060 11036
rect 26418 11024 26424 11036
rect 26476 11064 26482 11076
rect 27065 11067 27123 11073
rect 27065 11064 27077 11067
rect 26476 11036 27077 11064
rect 26476 11024 26482 11036
rect 27065 11033 27077 11036
rect 27111 11033 27123 11067
rect 27065 11027 27123 11033
rect 20714 10996 20720 11008
rect 20548 10968 20720 10996
rect 18463 10965 18475 10968
rect 18417 10959 18475 10965
rect 20714 10956 20720 10968
rect 20772 10956 20778 11008
rect 21910 10956 21916 11008
rect 21968 10956 21974 11008
rect 23014 10956 23020 11008
rect 23072 10996 23078 11008
rect 25961 10999 26019 11005
rect 25961 10996 25973 10999
rect 23072 10968 25973 10996
rect 23072 10956 23078 10968
rect 25961 10965 25973 10968
rect 26007 10965 26019 10999
rect 27616 10996 27644 11104
rect 27706 11092 27712 11144
rect 27764 11132 27770 11144
rect 27801 11135 27859 11141
rect 27801 11132 27813 11135
rect 27764 11104 27813 11132
rect 27764 11092 27770 11104
rect 27801 11101 27813 11104
rect 27847 11101 27859 11135
rect 27801 11095 27859 11101
rect 27890 11092 27896 11144
rect 27948 11092 27954 11144
rect 28261 11135 28319 11141
rect 28261 11101 28273 11135
rect 28307 11132 28319 11135
rect 28350 11132 28356 11144
rect 28307 11104 28356 11132
rect 28307 11101 28319 11104
rect 28261 11095 28319 11101
rect 28350 11092 28356 11104
rect 28408 11092 28414 11144
rect 28460 11141 28488 11172
rect 28445 11135 28503 11141
rect 28445 11101 28457 11135
rect 28491 11101 28503 11135
rect 28445 11095 28503 11101
rect 28721 11135 28779 11141
rect 28721 11101 28733 11135
rect 28767 11132 28779 11135
rect 28810 11132 28816 11144
rect 28767 11104 28816 11132
rect 28767 11101 28779 11104
rect 28721 11095 28779 11101
rect 28810 11092 28816 11104
rect 28868 11092 28874 11144
rect 29012 11141 29040 11172
rect 29748 11172 30196 11200
rect 28997 11135 29055 11141
rect 28997 11101 29009 11135
rect 29043 11101 29055 11135
rect 28997 11095 29055 11101
rect 29178 11092 29184 11144
rect 29236 11092 29242 11144
rect 29454 11092 29460 11144
rect 29512 11132 29518 11144
rect 29748 11141 29776 11172
rect 30190 11160 30196 11172
rect 30248 11160 30254 11212
rect 32214 11160 32220 11212
rect 32272 11200 32278 11212
rect 33042 11200 33048 11212
rect 32272 11172 33048 11200
rect 32272 11160 32278 11172
rect 33042 11160 33048 11172
rect 33100 11200 33106 11212
rect 33244 11209 33272 11240
rect 33612 11212 33640 11240
rect 33962 11228 33968 11280
rect 34020 11268 34026 11280
rect 38470 11268 38476 11280
rect 34020 11240 36584 11268
rect 34020 11228 34026 11240
rect 33137 11203 33195 11209
rect 33137 11200 33149 11203
rect 33100 11172 33149 11200
rect 33100 11160 33106 11172
rect 33137 11169 33149 11172
rect 33183 11169 33195 11203
rect 33137 11163 33195 11169
rect 33229 11203 33287 11209
rect 33229 11169 33241 11203
rect 33275 11169 33287 11203
rect 33229 11163 33287 11169
rect 33318 11160 33324 11212
rect 33376 11160 33382 11212
rect 33594 11160 33600 11212
rect 33652 11200 33658 11212
rect 35342 11200 35348 11212
rect 33652 11172 34100 11200
rect 33652 11160 33658 11172
rect 29549 11135 29607 11141
rect 29549 11132 29561 11135
rect 29512 11104 29561 11132
rect 29512 11092 29518 11104
rect 29549 11101 29561 11104
rect 29595 11101 29607 11135
rect 29549 11095 29607 11101
rect 29733 11135 29791 11141
rect 29733 11101 29745 11135
rect 29779 11101 29791 11135
rect 29733 11095 29791 11101
rect 29825 11135 29883 11141
rect 29825 11101 29837 11135
rect 29871 11129 29883 11135
rect 29932 11129 30512 11132
rect 29871 11104 30512 11129
rect 29871 11101 29960 11104
rect 29825 11095 29883 11101
rect 28629 11067 28687 11073
rect 28629 11033 28641 11067
rect 28675 11064 28687 11067
rect 29196 11064 29224 11092
rect 28675 11036 29224 11064
rect 28675 11033 28687 11036
rect 28629 11027 28687 11033
rect 28534 10996 28540 11008
rect 27616 10968 28540 10996
rect 25961 10959 26019 10965
rect 28534 10956 28540 10968
rect 28592 10956 28598 11008
rect 29086 10956 29092 11008
rect 29144 10996 29150 11008
rect 29273 10999 29331 11005
rect 29273 10996 29285 10999
rect 29144 10968 29285 10996
rect 29144 10956 29150 10968
rect 29273 10965 29285 10968
rect 29319 10996 29331 10999
rect 29454 10996 29460 11008
rect 29319 10968 29460 10996
rect 29319 10965 29331 10968
rect 29273 10959 29331 10965
rect 29454 10956 29460 10968
rect 29512 10956 29518 11008
rect 29822 10956 29828 11008
rect 29880 10996 29886 11008
rect 29932 10996 29960 11101
rect 30006 11024 30012 11076
rect 30064 11064 30070 11076
rect 30282 11064 30288 11076
rect 30064 11036 30288 11064
rect 30064 11024 30070 11036
rect 30282 11024 30288 11036
rect 30340 11024 30346 11076
rect 30484 11064 30512 11104
rect 30558 11092 30564 11144
rect 30616 11132 30622 11144
rect 30834 11132 30840 11144
rect 30616 11104 30840 11132
rect 30616 11092 30622 11104
rect 30834 11092 30840 11104
rect 30892 11092 30898 11144
rect 31757 11135 31815 11141
rect 31757 11101 31769 11135
rect 31803 11132 31815 11135
rect 32033 11135 32091 11141
rect 32033 11132 32045 11135
rect 31803 11104 32045 11132
rect 31803 11101 31815 11104
rect 31757 11095 31815 11101
rect 32033 11101 32045 11104
rect 32079 11101 32091 11135
rect 32033 11095 32091 11101
rect 30742 11064 30748 11076
rect 30484 11036 30748 11064
rect 30742 11024 30748 11036
rect 30800 11064 30806 11076
rect 30800 11036 31617 11064
rect 30800 11024 30806 11036
rect 29880 10968 29960 10996
rect 29880 10956 29886 10968
rect 30466 10956 30472 11008
rect 30524 10996 30530 11008
rect 31110 10996 31116 11008
rect 30524 10968 31116 10996
rect 30524 10956 30530 10968
rect 31110 10956 31116 10968
rect 31168 10956 31174 11008
rect 31589 10996 31617 11036
rect 31662 11024 31668 11076
rect 31720 11064 31726 11076
rect 31772 11064 31800 11095
rect 32858 11092 32864 11144
rect 32916 11092 32922 11144
rect 33410 11092 33416 11144
rect 33468 11092 33474 11144
rect 33870 11141 33876 11144
rect 33689 11135 33747 11141
rect 33689 11101 33701 11135
rect 33735 11101 33747 11135
rect 33689 11095 33747 11101
rect 33847 11135 33876 11141
rect 33847 11101 33859 11135
rect 33847 11095 33876 11101
rect 33318 11064 33324 11076
rect 31720 11036 31800 11064
rect 32048 11036 33324 11064
rect 31720 11024 31726 11036
rect 32048 10996 32076 11036
rect 33318 11024 33324 11036
rect 33376 11024 33382 11076
rect 33704 11064 33732 11095
rect 33870 11092 33876 11095
rect 33928 11092 33934 11144
rect 34072 11141 34100 11172
rect 34900 11172 35348 11200
rect 34057 11135 34115 11141
rect 34057 11101 34069 11135
rect 34103 11101 34115 11135
rect 34057 11095 34115 11101
rect 34149 11135 34207 11141
rect 34149 11101 34161 11135
rect 34195 11101 34207 11135
rect 34149 11095 34207 11101
rect 33704 11036 33824 11064
rect 31589 10968 32076 10996
rect 32122 10956 32128 11008
rect 32180 10996 32186 11008
rect 32674 10996 32680 11008
rect 32180 10968 32680 10996
rect 32180 10956 32186 10968
rect 32674 10956 32680 10968
rect 32732 10956 32738 11008
rect 32766 10956 32772 11008
rect 32824 10996 32830 11008
rect 32953 10999 33011 11005
rect 32953 10996 32965 10999
rect 32824 10968 32965 10996
rect 32824 10956 32830 10968
rect 32953 10965 32965 10968
rect 32999 10965 33011 10999
rect 33796 10996 33824 11036
rect 33962 11024 33968 11076
rect 34020 11024 34026 11076
rect 34164 11064 34192 11095
rect 34330 11092 34336 11144
rect 34388 11092 34394 11144
rect 34606 11092 34612 11144
rect 34664 11132 34670 11144
rect 34900 11141 34928 11172
rect 35342 11160 35348 11172
rect 35400 11200 35406 11212
rect 36265 11203 36323 11209
rect 36265 11200 36277 11203
rect 35400 11172 36277 11200
rect 35400 11160 35406 11172
rect 36265 11169 36277 11172
rect 36311 11169 36323 11203
rect 36265 11163 36323 11169
rect 34885 11135 34943 11141
rect 34885 11132 34897 11135
rect 34664 11104 34897 11132
rect 34664 11092 34670 11104
rect 34885 11101 34897 11104
rect 34931 11101 34943 11135
rect 34885 11095 34943 11101
rect 34974 11092 34980 11144
rect 35032 11092 35038 11144
rect 35253 11135 35311 11141
rect 35253 11101 35265 11135
rect 35299 11132 35311 11135
rect 35986 11132 35992 11144
rect 35299 11104 35992 11132
rect 35299 11101 35311 11104
rect 35253 11095 35311 11101
rect 35986 11092 35992 11104
rect 36044 11092 36050 11144
rect 36403 11135 36461 11141
rect 36403 11132 36415 11135
rect 36188 11104 36415 11132
rect 35069 11067 35127 11073
rect 35069 11064 35081 11067
rect 34164 11036 35081 11064
rect 35069 11033 35081 11036
rect 35115 11064 35127 11067
rect 36078 11064 36084 11076
rect 35115 11036 36084 11064
rect 35115 11033 35127 11036
rect 35069 11027 35127 11033
rect 36078 11024 36084 11036
rect 36136 11024 36142 11076
rect 34606 10996 34612 11008
rect 33796 10968 34612 10996
rect 32953 10959 33011 10965
rect 34606 10956 34612 10968
rect 34664 10956 34670 11008
rect 34698 10956 34704 11008
rect 34756 10956 34762 11008
rect 34882 10956 34888 11008
rect 34940 10996 34946 11008
rect 36188 10996 36216 11104
rect 36403 11101 36415 11104
rect 36449 11101 36461 11135
rect 36403 11095 36461 11101
rect 36556 11073 36584 11240
rect 36648 11240 38476 11268
rect 36648 11144 36676 11240
rect 38470 11228 38476 11240
rect 38528 11228 38534 11280
rect 37090 11160 37096 11212
rect 37148 11160 37154 11212
rect 39666 11200 39672 11212
rect 37200 11172 39672 11200
rect 36630 11092 36636 11144
rect 36688 11092 36694 11144
rect 36722 11092 36728 11144
rect 36780 11092 36786 11144
rect 37200 11132 37228 11172
rect 39666 11160 39672 11172
rect 39724 11160 39730 11212
rect 36832 11104 37228 11132
rect 36541 11067 36599 11073
rect 36541 11033 36553 11067
rect 36587 11064 36599 11067
rect 36832 11064 36860 11104
rect 37274 11092 37280 11144
rect 37332 11092 37338 11144
rect 36587 11036 36860 11064
rect 36909 11067 36967 11073
rect 36587 11033 36599 11036
rect 36541 11027 36599 11033
rect 36909 11033 36921 11067
rect 36955 11064 36967 11067
rect 37001 11067 37059 11073
rect 37001 11064 37013 11067
rect 36955 11036 37013 11064
rect 36955 11033 36967 11036
rect 36909 11027 36967 11033
rect 37001 11033 37013 11036
rect 37047 11033 37059 11067
rect 37001 11027 37059 11033
rect 34940 10968 36216 10996
rect 37461 10999 37519 11005
rect 34940 10956 34946 10968
rect 37461 10965 37473 10999
rect 37507 10996 37519 10999
rect 38286 10996 38292 11008
rect 37507 10968 38292 10996
rect 37507 10965 37519 10968
rect 37461 10959 37519 10965
rect 38286 10956 38292 10968
rect 38344 10956 38350 11008
rect 1104 10906 40572 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 40572 10906
rect 1104 10832 40572 10854
rect 7374 10752 7380 10804
rect 7432 10792 7438 10804
rect 7432 10764 7604 10792
rect 7432 10752 7438 10764
rect 5718 10684 5724 10736
rect 5776 10724 5782 10736
rect 7576 10733 7604 10764
rect 8404 10764 9168 10792
rect 8404 10736 8432 10764
rect 6641 10727 6699 10733
rect 6641 10724 6653 10727
rect 5776 10696 6653 10724
rect 5776 10684 5782 10696
rect 6641 10693 6653 10696
rect 6687 10693 6699 10727
rect 6641 10687 6699 10693
rect 7561 10727 7619 10733
rect 7561 10693 7573 10727
rect 7607 10724 7619 10727
rect 7650 10724 7656 10736
rect 7607 10696 7656 10724
rect 7607 10693 7619 10696
rect 7561 10687 7619 10693
rect 7650 10684 7656 10696
rect 7708 10724 7714 10736
rect 7708 10696 8064 10724
rect 7708 10684 7714 10696
rect 6546 10616 6552 10668
rect 6604 10616 6610 10668
rect 6730 10616 6736 10668
rect 6788 10616 6794 10668
rect 6914 10616 6920 10668
rect 6972 10616 6978 10668
rect 7193 10659 7251 10665
rect 7193 10625 7205 10659
rect 7239 10625 7251 10659
rect 7193 10619 7251 10625
rect 7208 10588 7236 10619
rect 7466 10616 7472 10668
rect 7524 10616 7530 10668
rect 7745 10659 7803 10665
rect 7745 10625 7757 10659
rect 7791 10656 7803 10659
rect 7926 10656 7932 10668
rect 7791 10628 7932 10656
rect 7791 10625 7803 10628
rect 7745 10619 7803 10625
rect 7760 10588 7788 10619
rect 7926 10616 7932 10628
rect 7984 10616 7990 10668
rect 8036 10665 8064 10696
rect 8386 10684 8392 10736
rect 8444 10684 8450 10736
rect 8589 10727 8647 10733
rect 8589 10724 8601 10727
rect 8588 10693 8601 10724
rect 8635 10693 8647 10727
rect 8588 10687 8647 10693
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 8202 10616 8208 10668
rect 8260 10616 8266 10668
rect 8588 10588 8616 10687
rect 8754 10684 8760 10736
rect 8812 10724 8818 10736
rect 9140 10733 9168 10764
rect 10042 10752 10048 10804
rect 10100 10792 10106 10804
rect 10137 10795 10195 10801
rect 10137 10792 10149 10795
rect 10100 10764 10149 10792
rect 10100 10752 10106 10764
rect 10137 10761 10149 10764
rect 10183 10761 10195 10795
rect 10137 10755 10195 10761
rect 10410 10752 10416 10804
rect 10468 10792 10474 10804
rect 14461 10795 14519 10801
rect 14461 10792 14473 10795
rect 10468 10764 14473 10792
rect 10468 10752 10474 10764
rect 14461 10761 14473 10764
rect 14507 10761 14519 10795
rect 14461 10755 14519 10761
rect 16942 10752 16948 10804
rect 17000 10752 17006 10804
rect 21818 10792 21824 10804
rect 21192 10764 21824 10792
rect 8941 10727 8999 10733
rect 8941 10724 8953 10727
rect 8812 10696 8953 10724
rect 8812 10684 8818 10696
rect 8941 10693 8953 10696
rect 8987 10693 8999 10727
rect 8941 10687 8999 10693
rect 9125 10727 9183 10733
rect 9125 10693 9137 10727
rect 9171 10724 9183 10727
rect 9585 10727 9643 10733
rect 9585 10724 9597 10727
rect 9171 10696 9597 10724
rect 9171 10693 9183 10696
rect 9125 10687 9183 10693
rect 9585 10693 9597 10696
rect 9631 10724 9643 10727
rect 10870 10724 10876 10736
rect 9631 10696 10088 10724
rect 9631 10693 9643 10696
rect 9585 10687 9643 10693
rect 8849 10659 8907 10665
rect 8849 10625 8861 10659
rect 8895 10625 8907 10659
rect 9858 10656 9864 10668
rect 9819 10628 9864 10656
rect 8849 10619 8907 10625
rect 8864 10588 8892 10619
rect 9858 10616 9864 10628
rect 9916 10616 9922 10668
rect 10060 10665 10088 10696
rect 10152 10696 10876 10724
rect 10152 10668 10180 10696
rect 10870 10684 10876 10696
rect 10928 10684 10934 10736
rect 12342 10684 12348 10736
rect 12400 10724 12406 10736
rect 12713 10727 12771 10733
rect 12713 10724 12725 10727
rect 12400 10696 12725 10724
rect 12400 10684 12406 10696
rect 12713 10693 12725 10696
rect 12759 10693 12771 10727
rect 12713 10687 12771 10693
rect 14734 10684 14740 10736
rect 14792 10724 14798 10736
rect 21082 10724 21088 10736
rect 14792 10696 15148 10724
rect 14792 10684 14798 10696
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 10045 10659 10103 10665
rect 10045 10625 10057 10659
rect 10091 10625 10103 10659
rect 10045 10619 10103 10625
rect 7208 10560 7788 10588
rect 8036 10560 8892 10588
rect 6362 10412 6368 10464
rect 6420 10412 6426 10464
rect 7006 10412 7012 10464
rect 7064 10412 7070 10464
rect 7374 10412 7380 10464
rect 7432 10452 7438 10464
rect 7929 10455 7987 10461
rect 7929 10452 7941 10455
rect 7432 10424 7941 10452
rect 7432 10412 7438 10424
rect 7929 10421 7941 10424
rect 7975 10452 7987 10455
rect 8036 10452 8064 10560
rect 9766 10548 9772 10600
rect 9824 10588 9830 10600
rect 9968 10588 9996 10619
rect 10134 10616 10140 10668
rect 10192 10616 10198 10668
rect 10229 10659 10287 10665
rect 10229 10625 10241 10659
rect 10275 10656 10287 10659
rect 11882 10656 11888 10668
rect 10275 10628 11888 10656
rect 10275 10625 10287 10628
rect 10229 10619 10287 10625
rect 9824 10560 9996 10588
rect 9824 10548 9830 10560
rect 9306 10480 9312 10532
rect 9364 10520 9370 10532
rect 10244 10520 10272 10619
rect 11882 10616 11888 10628
rect 11940 10616 11946 10668
rect 12434 10616 12440 10668
rect 12492 10616 12498 10668
rect 12618 10616 12624 10668
rect 12676 10616 12682 10668
rect 12805 10659 12863 10665
rect 12805 10625 12817 10659
rect 12851 10656 12863 10659
rect 12986 10656 12992 10668
rect 12851 10628 12992 10656
rect 12851 10625 12863 10628
rect 12805 10619 12863 10625
rect 12986 10616 12992 10628
rect 13044 10616 13050 10668
rect 14458 10616 14464 10668
rect 14516 10656 14522 10668
rect 15120 10665 15148 10696
rect 16960 10696 21088 10724
rect 14829 10659 14887 10665
rect 14829 10656 14841 10659
rect 14516 10628 14841 10656
rect 14516 10616 14522 10628
rect 14829 10625 14841 10628
rect 14875 10625 14887 10659
rect 14829 10619 14887 10625
rect 14921 10659 14979 10665
rect 14921 10625 14933 10659
rect 14967 10625 14979 10659
rect 14921 10619 14979 10625
rect 15105 10659 15163 10665
rect 15105 10625 15117 10659
rect 15151 10656 15163 10659
rect 15378 10656 15384 10668
rect 15151 10628 15384 10656
rect 15151 10625 15163 10628
rect 15105 10619 15163 10625
rect 14737 10591 14795 10597
rect 14737 10557 14749 10591
rect 14783 10588 14795 10591
rect 14936 10588 14964 10619
rect 15378 10616 15384 10628
rect 15436 10616 15442 10668
rect 16960 10665 16988 10696
rect 21082 10684 21088 10696
rect 21140 10684 21146 10736
rect 16945 10659 17003 10665
rect 16945 10625 16957 10659
rect 16991 10625 17003 10659
rect 16945 10619 17003 10625
rect 17129 10659 17187 10665
rect 17129 10625 17141 10659
rect 17175 10656 17187 10659
rect 20806 10656 20812 10668
rect 17175 10628 20812 10656
rect 17175 10625 17187 10628
rect 17129 10619 17187 10625
rect 20806 10616 20812 10628
rect 20864 10616 20870 10668
rect 20990 10616 20996 10668
rect 21048 10616 21054 10668
rect 21192 10665 21220 10764
rect 21818 10752 21824 10764
rect 21876 10752 21882 10804
rect 22462 10752 22468 10804
rect 22520 10792 22526 10804
rect 22557 10795 22615 10801
rect 22557 10792 22569 10795
rect 22520 10764 22569 10792
rect 22520 10752 22526 10764
rect 22557 10761 22569 10764
rect 22603 10761 22615 10795
rect 22557 10755 22615 10761
rect 23106 10752 23112 10804
rect 23164 10752 23170 10804
rect 24026 10752 24032 10804
rect 24084 10752 24090 10804
rect 25222 10792 25228 10804
rect 24228 10764 25228 10792
rect 22094 10684 22100 10736
rect 22152 10724 22158 10736
rect 24228 10733 24256 10764
rect 25222 10752 25228 10764
rect 25280 10792 25286 10804
rect 25280 10764 26004 10792
rect 25280 10752 25286 10764
rect 24213 10727 24271 10733
rect 24213 10724 24225 10727
rect 22152 10696 24225 10724
rect 22152 10684 22158 10696
rect 24213 10693 24225 10696
rect 24259 10693 24271 10727
rect 24213 10687 24271 10693
rect 24302 10684 24308 10736
rect 24360 10724 24366 10736
rect 24397 10727 24455 10733
rect 24397 10724 24409 10727
rect 24360 10696 24409 10724
rect 24360 10684 24366 10696
rect 24397 10693 24409 10696
rect 24443 10693 24455 10727
rect 24397 10687 24455 10693
rect 24486 10684 24492 10736
rect 24544 10724 24550 10736
rect 24544 10696 25176 10724
rect 24544 10684 24550 10696
rect 21177 10659 21235 10665
rect 21177 10625 21189 10659
rect 21223 10625 21235 10659
rect 21177 10619 21235 10625
rect 21266 10616 21272 10668
rect 21324 10616 21330 10668
rect 21361 10659 21419 10665
rect 21361 10625 21373 10659
rect 21407 10656 21419 10659
rect 21542 10656 21548 10668
rect 21407 10628 21548 10656
rect 21407 10625 21419 10628
rect 21361 10619 21419 10625
rect 21542 10616 21548 10628
rect 21600 10616 21606 10668
rect 21818 10616 21824 10668
rect 21876 10616 21882 10668
rect 22005 10659 22063 10665
rect 22005 10625 22017 10659
rect 22051 10656 22063 10659
rect 22462 10656 22468 10668
rect 22051 10628 22468 10656
rect 22051 10625 22063 10628
rect 22005 10619 22063 10625
rect 22462 10616 22468 10628
rect 22520 10616 22526 10668
rect 23014 10616 23020 10668
rect 23072 10616 23078 10668
rect 23293 10659 23351 10665
rect 23293 10625 23305 10659
rect 23339 10656 23351 10659
rect 23382 10656 23388 10668
rect 23339 10628 23388 10656
rect 23339 10625 23351 10628
rect 23293 10619 23351 10625
rect 23382 10616 23388 10628
rect 23440 10616 23446 10668
rect 23477 10659 23535 10665
rect 23477 10625 23489 10659
rect 23523 10656 23535 10659
rect 24762 10656 24768 10668
rect 23523 10628 24768 10656
rect 23523 10625 23535 10628
rect 23477 10619 23535 10625
rect 24762 10616 24768 10628
rect 24820 10616 24826 10668
rect 15194 10588 15200 10600
rect 14783 10560 15200 10588
rect 14783 10557 14795 10560
rect 14737 10551 14795 10557
rect 15194 10548 15200 10560
rect 15252 10548 15258 10600
rect 21284 10588 21312 10616
rect 21726 10588 21732 10600
rect 21284 10560 21732 10588
rect 21726 10548 21732 10560
rect 21784 10548 21790 10600
rect 21910 10548 21916 10600
rect 21968 10588 21974 10600
rect 22281 10591 22339 10597
rect 22281 10588 22293 10591
rect 21968 10560 22293 10588
rect 21968 10548 21974 10560
rect 22281 10557 22293 10560
rect 22327 10557 22339 10591
rect 22281 10551 22339 10557
rect 24673 10591 24731 10597
rect 24673 10557 24685 10591
rect 24719 10588 24731 10591
rect 24854 10588 24860 10600
rect 24719 10560 24860 10588
rect 24719 10557 24731 10560
rect 24673 10551 24731 10557
rect 24854 10548 24860 10560
rect 24912 10548 24918 10600
rect 25148 10588 25176 10696
rect 25406 10684 25412 10736
rect 25464 10684 25470 10736
rect 25314 10616 25320 10668
rect 25372 10656 25378 10668
rect 25777 10659 25835 10665
rect 25777 10656 25789 10659
rect 25372 10628 25789 10656
rect 25372 10616 25378 10628
rect 25777 10625 25789 10628
rect 25823 10625 25835 10659
rect 25777 10619 25835 10625
rect 25976 10588 26004 10764
rect 26050 10752 26056 10804
rect 26108 10792 26114 10804
rect 27798 10792 27804 10804
rect 26108 10764 27804 10792
rect 26108 10752 26114 10764
rect 27798 10752 27804 10764
rect 27856 10752 27862 10804
rect 27890 10752 27896 10804
rect 27948 10792 27954 10804
rect 28077 10795 28135 10801
rect 28077 10792 28089 10795
rect 27948 10764 28089 10792
rect 27948 10752 27954 10764
rect 28077 10761 28089 10764
rect 28123 10761 28135 10795
rect 28077 10755 28135 10761
rect 28350 10752 28356 10804
rect 28408 10792 28414 10804
rect 30653 10795 30711 10801
rect 30653 10792 30665 10795
rect 28408 10764 30665 10792
rect 28408 10752 28414 10764
rect 30653 10761 30665 10764
rect 30699 10761 30711 10795
rect 30653 10755 30711 10761
rect 31202 10752 31208 10804
rect 31260 10752 31266 10804
rect 31757 10795 31815 10801
rect 31757 10761 31769 10795
rect 31803 10761 31815 10795
rect 31757 10755 31815 10761
rect 26237 10727 26295 10733
rect 26237 10693 26249 10727
rect 26283 10724 26295 10727
rect 26418 10724 26424 10736
rect 26283 10696 26424 10724
rect 26283 10693 26295 10696
rect 26237 10687 26295 10693
rect 26418 10684 26424 10696
rect 26476 10684 26482 10736
rect 28534 10724 28540 10736
rect 27816 10696 28540 10724
rect 26050 10616 26056 10668
rect 26108 10656 26114 10668
rect 27525 10659 27583 10665
rect 27525 10656 27537 10659
rect 26108 10628 27537 10656
rect 26108 10616 26114 10628
rect 27525 10625 27537 10628
rect 27571 10625 27583 10659
rect 27525 10619 27583 10625
rect 27614 10616 27620 10668
rect 27672 10656 27678 10668
rect 27816 10665 27844 10696
rect 28534 10684 28540 10696
rect 28592 10684 28598 10736
rect 29638 10684 29644 10736
rect 29696 10684 29702 10736
rect 31772 10724 31800 10755
rect 32858 10752 32864 10804
rect 32916 10752 32922 10804
rect 37550 10792 37556 10804
rect 37292 10764 37556 10792
rect 31036 10696 31800 10724
rect 27709 10659 27767 10665
rect 27709 10656 27721 10659
rect 27672 10628 27721 10656
rect 27672 10616 27678 10628
rect 27709 10625 27721 10628
rect 27755 10625 27767 10659
rect 27709 10619 27767 10625
rect 27801 10659 27859 10665
rect 27801 10625 27813 10659
rect 27847 10625 27859 10659
rect 27801 10619 27859 10625
rect 27893 10659 27951 10665
rect 27893 10625 27905 10659
rect 27939 10625 27951 10659
rect 27893 10619 27951 10625
rect 27908 10588 27936 10619
rect 27982 10616 27988 10668
rect 28040 10656 28046 10668
rect 28169 10659 28227 10665
rect 28169 10656 28181 10659
rect 28040 10628 28181 10656
rect 28040 10616 28046 10628
rect 28169 10625 28181 10628
rect 28215 10625 28227 10659
rect 28169 10619 28227 10625
rect 28258 10616 28264 10668
rect 28316 10656 28322 10668
rect 28353 10659 28411 10665
rect 28353 10656 28365 10659
rect 28316 10628 28365 10656
rect 28316 10616 28322 10628
rect 28353 10625 28365 10628
rect 28399 10656 28411 10659
rect 28810 10656 28816 10668
rect 28399 10628 28816 10656
rect 28399 10625 28411 10628
rect 28353 10619 28411 10625
rect 28810 10616 28816 10628
rect 28868 10616 28874 10668
rect 29178 10616 29184 10668
rect 29236 10656 29242 10668
rect 29822 10656 29828 10668
rect 29236 10628 29828 10656
rect 29236 10616 29242 10628
rect 29822 10616 29828 10628
rect 29880 10616 29886 10668
rect 30282 10616 30288 10668
rect 30340 10616 30346 10668
rect 30834 10616 30840 10668
rect 30892 10616 30898 10668
rect 31036 10597 31064 10696
rect 32214 10684 32220 10736
rect 32272 10724 32278 10736
rect 32401 10727 32459 10733
rect 32401 10724 32413 10727
rect 32272 10696 32413 10724
rect 32272 10684 32278 10696
rect 32401 10693 32413 10696
rect 32447 10693 32459 10727
rect 32401 10687 32459 10693
rect 32493 10727 32551 10733
rect 32493 10693 32505 10727
rect 32539 10724 32551 10727
rect 33962 10724 33968 10736
rect 32539 10696 33968 10724
rect 32539 10693 32551 10696
rect 32493 10687 32551 10693
rect 33962 10684 33968 10696
rect 34020 10684 34026 10736
rect 34330 10684 34336 10736
rect 34388 10724 34394 10736
rect 37292 10733 37320 10764
rect 37550 10752 37556 10764
rect 37608 10752 37614 10804
rect 37277 10727 37335 10733
rect 37277 10724 37289 10727
rect 34388 10696 37289 10724
rect 34388 10684 34394 10696
rect 37277 10693 37289 10696
rect 37323 10693 37335 10727
rect 37277 10687 37335 10693
rect 38841 10727 38899 10733
rect 38841 10693 38853 10727
rect 38887 10724 38899 10727
rect 39114 10724 39120 10736
rect 38887 10696 39120 10724
rect 38887 10693 38899 10696
rect 38841 10687 38899 10693
rect 39114 10684 39120 10696
rect 39172 10684 39178 10736
rect 31110 10616 31116 10668
rect 31168 10656 31174 10668
rect 31389 10659 31447 10665
rect 31389 10656 31401 10659
rect 31168 10628 31401 10656
rect 31168 10616 31174 10628
rect 31389 10625 31401 10628
rect 31435 10656 31447 10659
rect 31435 10628 31708 10656
rect 31435 10625 31447 10628
rect 31389 10619 31447 10625
rect 31021 10591 31079 10597
rect 31021 10588 31033 10591
rect 25148 10560 25268 10588
rect 25976 10560 31033 10588
rect 9364 10492 10272 10520
rect 9364 10480 9370 10492
rect 11882 10480 11888 10532
rect 11940 10520 11946 10532
rect 18690 10520 18696 10532
rect 11940 10492 18696 10520
rect 11940 10480 11946 10492
rect 18690 10480 18696 10492
rect 18748 10480 18754 10532
rect 21637 10523 21695 10529
rect 21637 10489 21649 10523
rect 21683 10520 21695 10523
rect 22189 10523 22247 10529
rect 22189 10520 22201 10523
rect 21683 10492 22201 10520
rect 21683 10489 21695 10492
rect 21637 10483 21695 10489
rect 22189 10489 22201 10492
rect 22235 10489 22247 10523
rect 22189 10483 22247 10489
rect 24118 10480 24124 10532
rect 24176 10520 24182 10532
rect 25240 10520 25268 10560
rect 31021 10557 31033 10560
rect 31067 10557 31079 10591
rect 31573 10591 31631 10597
rect 31573 10588 31585 10591
rect 31021 10551 31079 10557
rect 31404 10560 31585 10588
rect 31404 10532 31432 10560
rect 31573 10557 31585 10560
rect 31619 10557 31631 10591
rect 31573 10551 31631 10557
rect 24176 10492 25160 10520
rect 25240 10492 28028 10520
rect 24176 10480 24182 10492
rect 7975 10424 8064 10452
rect 7975 10421 7987 10424
rect 7929 10415 7987 10421
rect 8110 10412 8116 10464
rect 8168 10412 8174 10464
rect 8478 10412 8484 10464
rect 8536 10452 8542 10464
rect 8573 10455 8631 10461
rect 8573 10452 8585 10455
rect 8536 10424 8585 10452
rect 8536 10412 8542 10424
rect 8573 10421 8585 10424
rect 8619 10421 8631 10455
rect 8573 10415 8631 10421
rect 8754 10412 8760 10464
rect 8812 10412 8818 10464
rect 9125 10455 9183 10461
rect 9125 10421 9137 10455
rect 9171 10452 9183 10455
rect 10226 10452 10232 10464
rect 9171 10424 10232 10452
rect 9171 10421 9183 10424
rect 9125 10415 9183 10421
rect 10226 10412 10232 10424
rect 10284 10412 10290 10464
rect 12989 10455 13047 10461
rect 12989 10421 13001 10455
rect 13035 10452 13047 10455
rect 13446 10452 13452 10464
rect 13035 10424 13452 10452
rect 13035 10421 13047 10424
rect 12989 10415 13047 10421
rect 13446 10412 13452 10424
rect 13504 10412 13510 10464
rect 14734 10412 14740 10464
rect 14792 10412 14798 10464
rect 15010 10412 15016 10464
rect 15068 10452 15074 10464
rect 15105 10455 15163 10461
rect 15105 10452 15117 10455
rect 15068 10424 15117 10452
rect 15068 10412 15074 10424
rect 15105 10421 15117 10424
rect 15151 10421 15163 10455
rect 15105 10415 15163 10421
rect 17034 10412 17040 10464
rect 17092 10452 17098 10464
rect 19518 10452 19524 10464
rect 17092 10424 19524 10452
rect 17092 10412 17098 10424
rect 19518 10412 19524 10424
rect 19576 10452 19582 10464
rect 20346 10452 20352 10464
rect 19576 10424 20352 10452
rect 19576 10412 19582 10424
rect 20346 10412 20352 10424
rect 20404 10412 20410 10464
rect 20990 10412 20996 10464
rect 21048 10452 21054 10464
rect 21818 10452 21824 10464
rect 21048 10424 21824 10452
rect 21048 10412 21054 10424
rect 21818 10412 21824 10424
rect 21876 10452 21882 10464
rect 22002 10452 22008 10464
rect 21876 10424 22008 10452
rect 21876 10412 21882 10424
rect 22002 10412 22008 10424
rect 22060 10412 22066 10464
rect 22097 10455 22155 10461
rect 22097 10421 22109 10455
rect 22143 10452 22155 10455
rect 22370 10452 22376 10464
rect 22143 10424 22376 10452
rect 22143 10421 22155 10424
rect 22097 10415 22155 10421
rect 22370 10412 22376 10424
rect 22428 10412 22434 10464
rect 24213 10455 24271 10461
rect 24213 10421 24225 10455
rect 24259 10452 24271 10455
rect 25038 10452 25044 10464
rect 24259 10424 25044 10452
rect 24259 10421 24271 10424
rect 24213 10415 24271 10421
rect 25038 10412 25044 10424
rect 25096 10412 25102 10464
rect 25132 10452 25160 10492
rect 26053 10455 26111 10461
rect 26053 10452 26065 10455
rect 25132 10424 26065 10452
rect 26053 10421 26065 10424
rect 26099 10421 26111 10455
rect 28000 10452 28028 10492
rect 28074 10480 28080 10532
rect 28132 10520 28138 10532
rect 28353 10523 28411 10529
rect 28353 10520 28365 10523
rect 28132 10492 28365 10520
rect 28132 10480 28138 10492
rect 28353 10489 28365 10492
rect 28399 10489 28411 10523
rect 28353 10483 28411 10489
rect 31386 10480 31392 10532
rect 31444 10480 31450 10532
rect 31680 10520 31708 10628
rect 31846 10616 31852 10668
rect 31904 10656 31910 10668
rect 31941 10659 31999 10665
rect 31941 10656 31953 10659
rect 31904 10628 31953 10656
rect 31904 10616 31910 10628
rect 31941 10625 31953 10628
rect 31987 10625 31999 10659
rect 31941 10619 31999 10625
rect 32306 10616 32312 10668
rect 32364 10616 32370 10668
rect 32582 10616 32588 10668
rect 32640 10656 32646 10668
rect 32677 10659 32735 10665
rect 32677 10656 32689 10659
rect 32640 10628 32689 10656
rect 32640 10616 32646 10628
rect 32677 10625 32689 10628
rect 32723 10625 32735 10659
rect 32677 10619 32735 10625
rect 32769 10659 32827 10665
rect 32769 10625 32781 10659
rect 32815 10656 32827 10659
rect 32858 10656 32864 10668
rect 32815 10628 32864 10656
rect 32815 10625 32827 10628
rect 32769 10619 32827 10625
rect 32858 10616 32864 10628
rect 32916 10616 32922 10668
rect 32950 10616 32956 10668
rect 33008 10656 33014 10668
rect 33045 10659 33103 10665
rect 33045 10656 33057 10659
rect 33008 10628 33057 10656
rect 33008 10616 33014 10628
rect 33045 10625 33057 10628
rect 33091 10625 33103 10659
rect 33045 10619 33103 10625
rect 33321 10659 33379 10665
rect 33321 10625 33333 10659
rect 33367 10656 33379 10659
rect 34698 10656 34704 10668
rect 33367 10628 34704 10656
rect 33367 10625 33379 10628
rect 33321 10619 33379 10625
rect 34698 10616 34704 10628
rect 34756 10616 34762 10668
rect 37550 10616 37556 10668
rect 37608 10616 37614 10668
rect 38286 10616 38292 10668
rect 38344 10616 38350 10668
rect 38473 10659 38531 10665
rect 38473 10625 38485 10659
rect 38519 10656 38531 10659
rect 39025 10659 39083 10665
rect 39025 10656 39037 10659
rect 38519 10628 39037 10656
rect 38519 10625 38531 10628
rect 38473 10619 38531 10625
rect 39025 10625 39037 10628
rect 39071 10656 39083 10659
rect 39206 10656 39212 10668
rect 39071 10628 39212 10656
rect 39071 10625 39083 10628
rect 39025 10619 39083 10625
rect 39206 10616 39212 10628
rect 39264 10616 39270 10668
rect 32122 10548 32128 10600
rect 32180 10588 32186 10600
rect 33137 10591 33195 10597
rect 33137 10588 33149 10591
rect 32180 10560 33149 10588
rect 32180 10548 32186 10560
rect 33137 10557 33149 10560
rect 33183 10557 33195 10591
rect 33137 10551 33195 10557
rect 31938 10520 31944 10532
rect 31680 10492 31944 10520
rect 31938 10480 31944 10492
rect 31996 10480 32002 10532
rect 33152 10520 33180 10551
rect 33226 10548 33232 10600
rect 33284 10548 33290 10600
rect 37461 10591 37519 10597
rect 37461 10557 37473 10591
rect 37507 10588 37519 10591
rect 37734 10588 37740 10600
rect 37507 10560 37740 10588
rect 37507 10557 37519 10560
rect 37461 10551 37519 10557
rect 37734 10548 37740 10560
rect 37792 10548 37798 10600
rect 34054 10520 34060 10532
rect 33152 10492 34060 10520
rect 34054 10480 34060 10492
rect 34112 10520 34118 10532
rect 36078 10520 36084 10532
rect 34112 10492 36084 10520
rect 34112 10480 34118 10492
rect 36078 10480 36084 10492
rect 36136 10480 36142 10532
rect 38746 10520 38752 10532
rect 38488 10492 38752 10520
rect 31110 10452 31116 10464
rect 28000 10424 31116 10452
rect 26053 10415 26111 10421
rect 31110 10412 31116 10424
rect 31168 10412 31174 10464
rect 32125 10455 32183 10461
rect 32125 10421 32137 10455
rect 32171 10452 32183 10455
rect 34698 10452 34704 10464
rect 32171 10424 34704 10452
rect 32171 10421 32183 10424
rect 32125 10415 32183 10421
rect 34698 10412 34704 10424
rect 34756 10412 34762 10464
rect 35342 10412 35348 10464
rect 35400 10452 35406 10464
rect 38488 10461 38516 10492
rect 38746 10480 38752 10492
rect 38804 10480 38810 10532
rect 37277 10455 37335 10461
rect 37277 10452 37289 10455
rect 35400 10424 37289 10452
rect 35400 10412 35406 10424
rect 37277 10421 37289 10424
rect 37323 10421 37335 10455
rect 37277 10415 37335 10421
rect 37737 10455 37795 10461
rect 37737 10421 37749 10455
rect 37783 10452 37795 10455
rect 38473 10455 38531 10461
rect 38473 10452 38485 10455
rect 37783 10424 38485 10452
rect 37783 10421 37795 10424
rect 37737 10415 37795 10421
rect 38473 10421 38485 10424
rect 38519 10421 38531 10455
rect 38473 10415 38531 10421
rect 38654 10412 38660 10464
rect 38712 10412 38718 10464
rect 39209 10455 39267 10461
rect 39209 10421 39221 10455
rect 39255 10452 39267 10455
rect 39390 10452 39396 10464
rect 39255 10424 39396 10452
rect 39255 10421 39267 10424
rect 39209 10415 39267 10421
rect 39390 10412 39396 10424
rect 39448 10412 39454 10464
rect 1104 10362 40572 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 40572 10362
rect 1104 10288 40572 10310
rect 4236 10251 4294 10257
rect 4236 10217 4248 10251
rect 4282 10248 4294 10251
rect 6362 10248 6368 10260
rect 4282 10220 6368 10248
rect 4282 10217 4294 10220
rect 4236 10211 4294 10217
rect 6362 10208 6368 10220
rect 6420 10208 6426 10260
rect 6730 10208 6736 10260
rect 6788 10248 6794 10260
rect 8662 10248 8668 10260
rect 6788 10220 8668 10248
rect 6788 10208 6794 10220
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 8754 10208 8760 10260
rect 8812 10248 8818 10260
rect 10137 10251 10195 10257
rect 10137 10248 10149 10251
rect 8812 10220 10149 10248
rect 8812 10208 8818 10220
rect 10137 10217 10149 10220
rect 10183 10217 10195 10251
rect 10137 10211 10195 10217
rect 12618 10208 12624 10260
rect 12676 10208 12682 10260
rect 14461 10251 14519 10257
rect 14461 10217 14473 10251
rect 14507 10217 14519 10251
rect 14461 10211 14519 10217
rect 5718 10140 5724 10192
rect 5776 10140 5782 10192
rect 6104 10152 8432 10180
rect 3510 10072 3516 10124
rect 3568 10112 3574 10124
rect 3973 10115 4031 10121
rect 3973 10112 3985 10115
rect 3568 10084 3985 10112
rect 3568 10072 3574 10084
rect 3973 10081 3985 10084
rect 4019 10112 4031 10115
rect 4019 10084 5580 10112
rect 4019 10081 4031 10084
rect 3973 10075 4031 10081
rect 4706 9936 4712 9988
rect 4764 9936 4770 9988
rect 5552 9976 5580 10084
rect 6104 10053 6132 10152
rect 7285 10115 7343 10121
rect 7285 10081 7297 10115
rect 7331 10081 7343 10115
rect 8110 10112 8116 10124
rect 7285 10075 7343 10081
rect 7484 10084 8116 10112
rect 6089 10047 6147 10053
rect 6089 10013 6101 10047
rect 6135 10013 6147 10047
rect 6089 10007 6147 10013
rect 7098 10004 7104 10056
rect 7156 10004 7162 10056
rect 6822 9976 6828 9988
rect 5552 9948 6828 9976
rect 6822 9936 6828 9948
rect 6880 9936 6886 9988
rect 7300 9976 7328 10075
rect 7374 10004 7380 10056
rect 7432 10004 7438 10056
rect 7484 10053 7512 10084
rect 8110 10072 8116 10084
rect 8168 10072 8174 10124
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 7558 10004 7564 10056
rect 7616 10004 7622 10056
rect 7650 10004 7656 10056
rect 7708 10044 7714 10056
rect 7745 10047 7803 10053
rect 7745 10044 7757 10047
rect 7708 10016 7757 10044
rect 7708 10004 7714 10016
rect 7745 10013 7757 10016
rect 7791 10013 7803 10047
rect 7745 10007 7803 10013
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10044 7895 10047
rect 7926 10044 7932 10056
rect 7883 10016 7932 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 7926 10004 7932 10016
rect 7984 10004 7990 10056
rect 8294 10004 8300 10056
rect 8352 10004 8358 10056
rect 8404 10044 8432 10152
rect 9582 10140 9588 10192
rect 9640 10180 9646 10192
rect 9640 10152 10088 10180
rect 9640 10140 9646 10152
rect 9030 10072 9036 10124
rect 9088 10112 9094 10124
rect 9953 10115 10011 10121
rect 9953 10112 9965 10115
rect 9088 10084 9965 10112
rect 9088 10072 9094 10084
rect 9953 10081 9965 10084
rect 9999 10081 10011 10115
rect 10060 10112 10088 10152
rect 10318 10140 10324 10192
rect 10376 10180 10382 10192
rect 11790 10180 11796 10192
rect 10376 10152 11796 10180
rect 10376 10140 10382 10152
rect 11790 10140 11796 10152
rect 11848 10180 11854 10192
rect 14476 10180 14504 10211
rect 14550 10208 14556 10260
rect 14608 10248 14614 10260
rect 14918 10248 14924 10260
rect 14608 10220 14924 10248
rect 14608 10208 14614 10220
rect 14918 10208 14924 10220
rect 14976 10208 14982 10260
rect 16850 10208 16856 10260
rect 16908 10208 16914 10260
rect 18690 10208 18696 10260
rect 18748 10208 18754 10260
rect 19061 10251 19119 10257
rect 19061 10217 19073 10251
rect 19107 10217 19119 10251
rect 19061 10211 19119 10217
rect 11848 10152 14504 10180
rect 11848 10140 11854 10152
rect 12434 10112 12440 10124
rect 10060 10084 12440 10112
rect 9953 10075 10011 10081
rect 8941 10047 8999 10053
rect 8941 10044 8953 10047
rect 8404 10016 8953 10044
rect 8941 10013 8953 10016
rect 8987 10044 8999 10047
rect 9968 10044 9996 10075
rect 12434 10072 12440 10084
rect 12492 10112 12498 10124
rect 15105 10115 15163 10121
rect 15105 10112 15117 10115
rect 12492 10084 15117 10112
rect 12492 10072 12498 10084
rect 15105 10081 15117 10084
rect 15151 10081 15163 10115
rect 16868 10112 16896 10208
rect 19076 10180 19104 10211
rect 19518 10208 19524 10260
rect 19576 10208 19582 10260
rect 19628 10220 19840 10248
rect 19628 10180 19656 10220
rect 19076 10152 19656 10180
rect 19705 10183 19763 10189
rect 19705 10149 19717 10183
rect 19751 10149 19763 10183
rect 19812 10180 19840 10220
rect 20346 10208 20352 10260
rect 20404 10248 20410 10260
rect 25685 10251 25743 10257
rect 25685 10248 25697 10251
rect 20404 10220 25697 10248
rect 20404 10208 20410 10220
rect 25685 10217 25697 10220
rect 25731 10217 25743 10251
rect 25685 10211 25743 10217
rect 26602 10208 26608 10260
rect 26660 10248 26666 10260
rect 26697 10251 26755 10257
rect 26697 10248 26709 10251
rect 26660 10220 26709 10248
rect 26660 10208 26666 10220
rect 26697 10217 26709 10220
rect 26743 10217 26755 10251
rect 26697 10211 26755 10217
rect 27706 10208 27712 10260
rect 27764 10248 27770 10260
rect 28074 10248 28080 10260
rect 27764 10220 28080 10248
rect 27764 10208 27770 10220
rect 28074 10208 28080 10220
rect 28132 10208 28138 10260
rect 28537 10251 28595 10257
rect 28537 10217 28549 10251
rect 28583 10248 28595 10251
rect 29178 10248 29184 10260
rect 28583 10220 29184 10248
rect 28583 10217 28595 10220
rect 28537 10211 28595 10217
rect 29178 10208 29184 10220
rect 29236 10248 29242 10260
rect 29236 10220 29408 10248
rect 29236 10208 29242 10220
rect 19978 10180 19984 10192
rect 19812 10152 19984 10180
rect 19705 10143 19763 10149
rect 18969 10115 19027 10121
rect 16868 10084 18000 10112
rect 15105 10075 15163 10081
rect 10134 10044 10140 10056
rect 8987 10016 9812 10044
rect 9968 10016 10140 10044
rect 8987 10013 8999 10016
rect 8941 10007 8999 10013
rect 8312 9976 8340 10004
rect 9582 9976 9588 9988
rect 7300 9948 7788 9976
rect 8312 9948 9588 9976
rect 7760 9920 7788 9948
rect 9582 9936 9588 9948
rect 9640 9976 9646 9988
rect 9677 9979 9735 9985
rect 9677 9976 9689 9979
rect 9640 9948 9689 9976
rect 9640 9936 9646 9948
rect 9677 9945 9689 9948
rect 9723 9945 9735 9979
rect 9784 9976 9812 10016
rect 10134 10004 10140 10016
rect 10192 10004 10198 10056
rect 10226 10004 10232 10056
rect 10284 10004 10290 10056
rect 10686 10004 10692 10056
rect 10744 10044 10750 10056
rect 11333 10047 11391 10053
rect 11333 10044 11345 10047
rect 10744 10016 11345 10044
rect 10744 10004 10750 10016
rect 11333 10013 11345 10016
rect 11379 10013 11391 10047
rect 11333 10007 11391 10013
rect 11514 10004 11520 10056
rect 11572 10004 11578 10056
rect 11624 10016 12664 10044
rect 11624 9976 11652 10016
rect 9784 9948 11652 9976
rect 9677 9939 9735 9945
rect 11882 9936 11888 9988
rect 11940 9976 11946 9988
rect 12253 9979 12311 9985
rect 12253 9976 12265 9979
rect 11940 9948 12265 9976
rect 11940 9936 11946 9948
rect 12253 9945 12265 9948
rect 12299 9945 12311 9979
rect 12253 9939 12311 9945
rect 12437 9979 12495 9985
rect 12437 9945 12449 9979
rect 12483 9976 12495 9979
rect 12526 9976 12532 9988
rect 12483 9948 12532 9976
rect 12483 9945 12495 9948
rect 12437 9939 12495 9945
rect 12526 9936 12532 9948
rect 12584 9936 12590 9988
rect 12636 9976 12664 10016
rect 12710 10004 12716 10056
rect 12768 10004 12774 10056
rect 12802 10004 12808 10056
rect 12860 10044 12866 10056
rect 12897 10047 12955 10053
rect 12897 10044 12909 10047
rect 12860 10016 12909 10044
rect 12860 10004 12866 10016
rect 12897 10013 12909 10016
rect 12943 10013 12955 10047
rect 12897 10007 12955 10013
rect 14645 10047 14703 10053
rect 14645 10013 14657 10047
rect 14691 10044 14703 10047
rect 15010 10044 15016 10056
rect 14691 10016 15016 10044
rect 14691 10013 14703 10016
rect 14645 10007 14703 10013
rect 15010 10004 15016 10016
rect 15068 10004 15074 10056
rect 17218 10004 17224 10056
rect 17276 10004 17282 10056
rect 17586 10004 17592 10056
rect 17644 10004 17650 10056
rect 17972 10053 18000 10084
rect 18969 10081 18981 10115
rect 19015 10112 19027 10115
rect 19015 10084 19288 10112
rect 19015 10081 19027 10084
rect 18969 10075 19027 10081
rect 17681 10047 17739 10053
rect 17681 10013 17693 10047
rect 17727 10044 17739 10047
rect 17865 10047 17923 10053
rect 17865 10044 17877 10047
rect 17727 10016 17877 10044
rect 17727 10013 17739 10016
rect 17681 10007 17739 10013
rect 17865 10013 17877 10016
rect 17911 10013 17923 10047
rect 17865 10007 17923 10013
rect 17957 10047 18015 10053
rect 17957 10013 17969 10047
rect 18003 10013 18015 10047
rect 17957 10007 18015 10013
rect 12636 9948 12940 9976
rect 7193 9911 7251 9917
rect 7193 9877 7205 9911
rect 7239 9908 7251 9911
rect 7282 9908 7288 9920
rect 7239 9880 7288 9908
rect 7239 9877 7251 9880
rect 7193 9871 7251 9877
rect 7282 9868 7288 9880
rect 7340 9868 7346 9920
rect 7650 9868 7656 9920
rect 7708 9868 7714 9920
rect 7742 9868 7748 9920
rect 7800 9908 7806 9920
rect 9030 9908 9036 9920
rect 7800 9880 9036 9908
rect 7800 9868 7806 9880
rect 9030 9868 9036 9880
rect 9088 9868 9094 9920
rect 9306 9868 9312 9920
rect 9364 9908 9370 9920
rect 9953 9911 10011 9917
rect 9953 9908 9965 9911
rect 9364 9880 9965 9908
rect 9364 9868 9370 9880
rect 9953 9877 9965 9880
rect 9999 9877 10011 9911
rect 9953 9871 10011 9877
rect 11054 9868 11060 9920
rect 11112 9908 11118 9920
rect 11425 9911 11483 9917
rect 11425 9908 11437 9911
rect 11112 9880 11437 9908
rect 11112 9868 11118 9880
rect 11425 9877 11437 9880
rect 11471 9877 11483 9911
rect 11425 9871 11483 9877
rect 12802 9868 12808 9920
rect 12860 9868 12866 9920
rect 12912 9908 12940 9948
rect 14366 9936 14372 9988
rect 14424 9976 14430 9988
rect 14737 9979 14795 9985
rect 14737 9976 14749 9979
rect 14424 9948 14749 9976
rect 14424 9936 14430 9948
rect 14737 9945 14749 9948
rect 14783 9945 14795 9979
rect 14737 9939 14795 9945
rect 15378 9936 15384 9988
rect 15436 9936 15442 9988
rect 15488 9948 15870 9976
rect 14642 9908 14648 9920
rect 12912 9880 14648 9908
rect 14642 9868 14648 9880
rect 14700 9868 14706 9920
rect 14826 9868 14832 9920
rect 14884 9908 14890 9920
rect 15488 9908 15516 9948
rect 17310 9936 17316 9988
rect 17368 9936 17374 9988
rect 17402 9936 17408 9988
rect 17460 9936 17466 9988
rect 14884 9880 15516 9908
rect 14884 9868 14890 9880
rect 17034 9868 17040 9920
rect 17092 9868 17098 9920
rect 17328 9908 17356 9936
rect 17770 9908 17776 9920
rect 17328 9880 17776 9908
rect 17770 9868 17776 9880
rect 17828 9868 17834 9920
rect 17972 9908 18000 10007
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 19058 10044 19064 10056
rect 18380 10016 19064 10044
rect 18380 10004 18386 10016
rect 19058 10004 19064 10016
rect 19116 10004 19122 10056
rect 19260 10044 19288 10084
rect 19334 10072 19340 10124
rect 19392 10072 19398 10124
rect 19610 10072 19616 10124
rect 19668 10112 19674 10124
rect 19720 10112 19748 10143
rect 19978 10140 19984 10152
rect 20036 10140 20042 10192
rect 24302 10140 24308 10192
rect 24360 10180 24366 10192
rect 24360 10152 26004 10180
rect 24360 10140 24366 10152
rect 25130 10112 25136 10124
rect 19668 10084 19748 10112
rect 19904 10084 25136 10112
rect 19668 10072 19674 10084
rect 19260 10016 19472 10044
rect 19444 9988 19472 10016
rect 19518 10004 19524 10056
rect 19576 10004 19582 10056
rect 19904 10044 19932 10084
rect 19720 10016 19932 10044
rect 19242 9936 19248 9988
rect 19300 9936 19306 9988
rect 19426 9936 19432 9988
rect 19484 9976 19490 9988
rect 19720 9976 19748 10016
rect 19978 10004 19984 10056
rect 20036 10004 20042 10056
rect 20088 10053 20116 10084
rect 25130 10072 25136 10084
rect 25188 10072 25194 10124
rect 25774 10112 25780 10124
rect 25332 10084 25780 10112
rect 25332 10056 25360 10084
rect 25774 10072 25780 10084
rect 25832 10072 25838 10124
rect 20073 10047 20131 10053
rect 20073 10013 20085 10047
rect 20119 10013 20131 10047
rect 20073 10007 20131 10013
rect 23842 10004 23848 10056
rect 23900 10044 23906 10056
rect 24302 10044 24308 10056
rect 23900 10016 24308 10044
rect 23900 10004 23906 10016
rect 24302 10004 24308 10016
rect 24360 10004 24366 10056
rect 24854 10004 24860 10056
rect 24912 10004 24918 10056
rect 25314 10004 25320 10056
rect 25372 10004 25378 10056
rect 25590 10004 25596 10056
rect 25648 10004 25654 10056
rect 25976 10053 26004 10152
rect 26620 10112 26648 10208
rect 27798 10140 27804 10192
rect 27856 10180 27862 10192
rect 28905 10183 28963 10189
rect 28905 10180 28917 10183
rect 27856 10152 28917 10180
rect 27856 10140 27862 10152
rect 28905 10149 28917 10152
rect 28951 10149 28963 10183
rect 28905 10143 28963 10149
rect 28997 10183 29055 10189
rect 28997 10149 29009 10183
rect 29043 10149 29055 10183
rect 28997 10143 29055 10149
rect 26068 10084 26648 10112
rect 26068 10053 26096 10084
rect 27154 10072 27160 10124
rect 27212 10112 27218 10124
rect 27212 10084 28580 10112
rect 27212 10072 27218 10084
rect 25961 10047 26019 10053
rect 25961 10013 25973 10047
rect 26007 10013 26019 10047
rect 25961 10007 26019 10013
rect 26053 10047 26111 10053
rect 26053 10013 26065 10047
rect 26099 10013 26111 10047
rect 26053 10007 26111 10013
rect 26329 10047 26387 10053
rect 26329 10013 26341 10047
rect 26375 10013 26387 10047
rect 26329 10007 26387 10013
rect 19484 9948 19748 9976
rect 19484 9936 19490 9948
rect 19794 9936 19800 9988
rect 19852 9936 19858 9988
rect 19996 9976 20024 10004
rect 25406 9976 25412 9988
rect 19996 9948 25412 9976
rect 25406 9936 25412 9948
rect 25464 9936 25470 9988
rect 25501 9979 25559 9985
rect 25501 9945 25513 9979
rect 25547 9976 25559 9979
rect 26234 9976 26240 9988
rect 25547 9948 26240 9976
rect 25547 9945 25559 9948
rect 25501 9939 25559 9945
rect 26234 9936 26240 9948
rect 26292 9936 26298 9988
rect 24394 9908 24400 9920
rect 17972 9880 24400 9908
rect 24394 9868 24400 9880
rect 24452 9868 24458 9920
rect 25130 9868 25136 9920
rect 25188 9868 25194 9920
rect 26142 9868 26148 9920
rect 26200 9868 26206 9920
rect 26344 9908 26372 10007
rect 26418 10004 26424 10056
rect 26476 10004 26482 10056
rect 26513 10047 26571 10053
rect 26513 10013 26525 10047
rect 26559 10013 26571 10047
rect 26513 10007 26571 10013
rect 26697 10047 26755 10053
rect 26697 10013 26709 10047
rect 26743 10044 26755 10047
rect 27614 10044 27620 10056
rect 26743 10016 27620 10044
rect 26743 10013 26755 10016
rect 26697 10007 26755 10013
rect 26528 9976 26556 10007
rect 27614 10004 27620 10016
rect 27672 10004 27678 10056
rect 27724 10053 27752 10084
rect 27709 10047 27767 10053
rect 27709 10013 27721 10047
rect 27755 10013 27767 10047
rect 28077 10047 28135 10053
rect 28077 10044 28089 10047
rect 27709 10007 27767 10013
rect 27908 10016 28089 10044
rect 27338 9976 27344 9988
rect 26528 9948 27344 9976
rect 27338 9936 27344 9948
rect 27396 9936 27402 9988
rect 27908 9920 27936 10016
rect 28077 10013 28089 10016
rect 28123 10013 28135 10047
rect 28077 10007 28135 10013
rect 28442 10004 28448 10056
rect 28500 10004 28506 10056
rect 28552 9976 28580 10084
rect 28626 10004 28632 10056
rect 28684 10044 28690 10056
rect 28721 10047 28779 10053
rect 28721 10044 28733 10047
rect 28684 10016 28733 10044
rect 28684 10004 28690 10016
rect 28721 10013 28733 10016
rect 28767 10044 28779 10047
rect 29012 10044 29040 10143
rect 29380 10121 29408 10220
rect 30650 10208 30656 10260
rect 30708 10248 30714 10260
rect 30837 10251 30895 10257
rect 30837 10248 30849 10251
rect 30708 10220 30849 10248
rect 30708 10208 30714 10220
rect 30837 10217 30849 10220
rect 30883 10248 30895 10251
rect 30926 10248 30932 10260
rect 30883 10220 30932 10248
rect 30883 10217 30895 10220
rect 30837 10211 30895 10217
rect 30926 10208 30932 10220
rect 30984 10208 30990 10260
rect 31036 10220 31524 10248
rect 31036 10180 31064 10220
rect 29472 10152 31064 10180
rect 29365 10115 29423 10121
rect 29365 10081 29377 10115
rect 29411 10081 29423 10115
rect 29365 10075 29423 10081
rect 28767 10016 29040 10044
rect 28767 10013 28779 10016
rect 28721 10007 28779 10013
rect 29086 10004 29092 10056
rect 29144 10044 29150 10056
rect 29472 10044 29500 10152
rect 31110 10140 31116 10192
rect 31168 10180 31174 10192
rect 31386 10180 31392 10192
rect 31168 10152 31392 10180
rect 31168 10140 31174 10152
rect 31386 10140 31392 10152
rect 31444 10140 31450 10192
rect 31496 10180 31524 10220
rect 31754 10208 31760 10260
rect 31812 10248 31818 10260
rect 32309 10251 32367 10257
rect 32309 10248 32321 10251
rect 31812 10220 32321 10248
rect 31812 10208 31818 10220
rect 32309 10217 32321 10220
rect 32355 10217 32367 10251
rect 32309 10211 32367 10217
rect 32766 10208 32772 10260
rect 32824 10208 32830 10260
rect 33410 10248 33416 10260
rect 32876 10220 33416 10248
rect 32493 10183 32551 10189
rect 31496 10152 32444 10180
rect 29546 10072 29552 10124
rect 29604 10112 29610 10124
rect 29641 10115 29699 10121
rect 29641 10112 29653 10115
rect 29604 10084 29653 10112
rect 29604 10072 29610 10084
rect 29641 10081 29653 10084
rect 29687 10081 29699 10115
rect 32416 10112 32444 10152
rect 32493 10149 32505 10183
rect 32539 10180 32551 10183
rect 32876 10180 32904 10220
rect 33410 10208 33416 10220
rect 33468 10208 33474 10260
rect 34698 10208 34704 10260
rect 34756 10248 34762 10260
rect 36725 10251 36783 10257
rect 36725 10248 36737 10251
rect 34756 10220 36737 10248
rect 34756 10208 34762 10220
rect 36725 10217 36737 10220
rect 36771 10248 36783 10251
rect 37274 10248 37280 10260
rect 36771 10220 37280 10248
rect 36771 10217 36783 10220
rect 36725 10211 36783 10217
rect 37274 10208 37280 10220
rect 37332 10208 37338 10260
rect 32539 10152 32904 10180
rect 32953 10183 33011 10189
rect 32539 10149 32551 10152
rect 32493 10143 32551 10149
rect 32953 10149 32965 10183
rect 32999 10180 33011 10183
rect 32999 10152 35848 10180
rect 32999 10149 33011 10152
rect 32953 10143 33011 10149
rect 35158 10112 35164 10124
rect 29641 10075 29699 10081
rect 30484 10084 31156 10112
rect 32416 10084 35164 10112
rect 29144 10016 29500 10044
rect 29144 10004 29150 10016
rect 29822 10004 29828 10056
rect 29880 10004 29886 10056
rect 30009 10047 30067 10053
rect 30009 10013 30021 10047
rect 30055 10044 30067 10047
rect 30098 10044 30104 10056
rect 30055 10016 30104 10044
rect 30055 10013 30067 10016
rect 30009 10007 30067 10013
rect 30098 10004 30104 10016
rect 30156 10004 30162 10056
rect 30484 9976 30512 10084
rect 30561 10047 30619 10053
rect 30561 10013 30573 10047
rect 30607 10013 30619 10047
rect 30561 10007 30619 10013
rect 30653 10047 30711 10053
rect 30653 10013 30665 10047
rect 30699 10044 30711 10047
rect 30742 10044 30748 10056
rect 30699 10016 30748 10044
rect 30699 10013 30711 10016
rect 30653 10007 30711 10013
rect 28552 9948 30512 9976
rect 30576 9976 30604 10007
rect 30742 10004 30748 10016
rect 30800 10004 30806 10056
rect 31128 10053 31156 10084
rect 35158 10072 35164 10084
rect 35216 10072 35222 10124
rect 31113 10047 31171 10053
rect 31113 10013 31125 10047
rect 31159 10044 31171 10047
rect 31386 10044 31392 10056
rect 31159 10016 31392 10044
rect 31159 10013 31171 10016
rect 31113 10007 31171 10013
rect 31386 10004 31392 10016
rect 31444 10004 31450 10056
rect 32030 10004 32036 10056
rect 32088 10044 32094 10056
rect 32585 10047 32643 10053
rect 32585 10044 32597 10047
rect 32088 10016 32597 10044
rect 32088 10004 32094 10016
rect 32585 10013 32597 10016
rect 32631 10013 32643 10047
rect 32585 10007 32643 10013
rect 32674 10004 32680 10056
rect 32732 10044 32738 10056
rect 32769 10047 32827 10053
rect 32769 10044 32781 10047
rect 32732 10016 32781 10044
rect 32732 10004 32738 10016
rect 32769 10013 32781 10016
rect 32815 10013 32827 10047
rect 32769 10007 32827 10013
rect 33042 10004 33048 10056
rect 33100 10044 33106 10056
rect 34514 10044 34520 10056
rect 33100 10016 34520 10044
rect 33100 10004 33106 10016
rect 34514 10004 34520 10016
rect 34572 10004 34578 10056
rect 35066 10004 35072 10056
rect 35124 10044 35130 10056
rect 35820 10044 35848 10152
rect 36909 10115 36967 10121
rect 36909 10081 36921 10115
rect 36955 10112 36967 10115
rect 37182 10112 37188 10124
rect 36955 10084 37188 10112
rect 36955 10081 36967 10084
rect 36909 10075 36967 10081
rect 37182 10072 37188 10084
rect 37240 10072 37246 10124
rect 38194 10072 38200 10124
rect 38252 10112 38258 10124
rect 39669 10115 39727 10121
rect 39669 10112 39681 10115
rect 38252 10084 39681 10112
rect 38252 10072 38258 10084
rect 39669 10081 39681 10084
rect 39715 10081 39727 10115
rect 39669 10075 39727 10081
rect 37001 10047 37059 10053
rect 37001 10044 37013 10047
rect 35124 10016 35756 10044
rect 35820 10016 37013 10044
rect 35124 10004 35130 10016
rect 32122 9976 32128 9988
rect 30576 9948 32128 9976
rect 26878 9908 26884 9920
rect 26344 9880 26884 9908
rect 26878 9868 26884 9880
rect 26936 9868 26942 9920
rect 27890 9868 27896 9920
rect 27948 9868 27954 9920
rect 28258 9868 28264 9920
rect 28316 9868 28322 9920
rect 30466 9868 30472 9920
rect 30524 9908 30530 9920
rect 30576 9908 30604 9948
rect 32122 9936 32128 9948
rect 32180 9936 32186 9988
rect 32341 9979 32399 9985
rect 32341 9945 32353 9979
rect 32387 9976 32399 9979
rect 32950 9976 32956 9988
rect 32387 9948 32956 9976
rect 32387 9945 32399 9948
rect 32341 9939 32399 9945
rect 32950 9936 32956 9948
rect 33008 9936 33014 9988
rect 33778 9936 33784 9988
rect 33836 9976 33842 9988
rect 35621 9979 35679 9985
rect 35621 9976 35633 9979
rect 33836 9948 35633 9976
rect 33836 9936 33842 9948
rect 35621 9945 35633 9948
rect 35667 9945 35679 9979
rect 35728 9976 35756 10016
rect 37001 10013 37013 10016
rect 37047 10044 37059 10047
rect 37550 10044 37556 10056
rect 37047 10016 37556 10044
rect 37047 10013 37059 10016
rect 37001 10007 37059 10013
rect 37550 10004 37556 10016
rect 37608 10004 37614 10056
rect 37826 10004 37832 10056
rect 37884 10004 37890 10056
rect 37918 10004 37924 10056
rect 37976 10004 37982 10056
rect 36354 9976 36360 9988
rect 35728 9948 36360 9976
rect 35621 9939 35679 9945
rect 36354 9936 36360 9948
rect 36412 9976 36418 9988
rect 36630 9976 36636 9988
rect 36412 9948 36636 9976
rect 36412 9936 36418 9948
rect 36630 9936 36636 9948
rect 36688 9936 36694 9988
rect 36725 9979 36783 9985
rect 36725 9945 36737 9979
rect 36771 9976 36783 9979
rect 37936 9976 37964 10004
rect 36771 9948 37964 9976
rect 38962 9948 39068 9976
rect 36771 9945 36783 9948
rect 36725 9939 36783 9945
rect 39040 9920 39068 9948
rect 39390 9936 39396 9988
rect 39448 9936 39454 9988
rect 30524 9880 30604 9908
rect 30524 9868 30530 9880
rect 30926 9868 30932 9920
rect 30984 9868 30990 9920
rect 31386 9868 31392 9920
rect 31444 9908 31450 9920
rect 35250 9908 35256 9920
rect 31444 9880 35256 9908
rect 31444 9868 31450 9880
rect 35250 9868 35256 9880
rect 35308 9868 35314 9920
rect 35434 9868 35440 9920
rect 35492 9908 35498 9920
rect 35713 9911 35771 9917
rect 35713 9908 35725 9911
rect 35492 9880 35725 9908
rect 35492 9868 35498 9880
rect 35713 9877 35725 9880
rect 35759 9877 35771 9911
rect 35713 9871 35771 9877
rect 37185 9911 37243 9917
rect 37185 9877 37197 9911
rect 37231 9908 37243 9911
rect 37366 9908 37372 9920
rect 37231 9880 37372 9908
rect 37231 9877 37243 9880
rect 37185 9871 37243 9877
rect 37366 9868 37372 9880
rect 37424 9868 37430 9920
rect 37458 9868 37464 9920
rect 37516 9908 37522 9920
rect 37645 9911 37703 9917
rect 37645 9908 37657 9911
rect 37516 9880 37657 9908
rect 37516 9868 37522 9880
rect 37645 9877 37657 9880
rect 37691 9877 37703 9911
rect 37645 9871 37703 9877
rect 37918 9868 37924 9920
rect 37976 9868 37982 9920
rect 39022 9868 39028 9920
rect 39080 9868 39086 9920
rect 1104 9818 40572 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 40572 9818
rect 1104 9744 40572 9766
rect 8205 9707 8263 9713
rect 8205 9673 8217 9707
rect 8251 9704 8263 9707
rect 8478 9704 8484 9716
rect 8251 9676 8484 9704
rect 8251 9673 8263 9676
rect 8205 9667 8263 9673
rect 8478 9664 8484 9676
rect 8536 9664 8542 9716
rect 8662 9664 8668 9716
rect 8720 9704 8726 9716
rect 8941 9707 8999 9713
rect 8941 9704 8953 9707
rect 8720 9676 8953 9704
rect 8720 9664 8726 9676
rect 8941 9673 8953 9676
rect 8987 9673 8999 9707
rect 8941 9667 8999 9673
rect 9232 9676 9444 9704
rect 9232 9636 9260 9676
rect 8128 9608 9260 9636
rect 6822 9528 6828 9580
rect 6880 9528 6886 9580
rect 7006 9528 7012 9580
rect 7064 9528 7070 9580
rect 7193 9571 7251 9577
rect 7193 9537 7205 9571
rect 7239 9568 7251 9571
rect 7650 9568 7656 9580
rect 7239 9540 7656 9568
rect 7239 9537 7251 9540
rect 7193 9531 7251 9537
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 8128 9577 8156 9608
rect 9306 9596 9312 9648
rect 9364 9596 9370 9648
rect 9416 9636 9444 9676
rect 11514 9664 11520 9716
rect 11572 9704 11578 9716
rect 12342 9704 12348 9716
rect 11572 9676 12348 9704
rect 11572 9664 11578 9676
rect 12342 9664 12348 9676
rect 12400 9704 12406 9716
rect 12529 9707 12587 9713
rect 12529 9704 12541 9707
rect 12400 9676 12541 9704
rect 12400 9664 12406 9676
rect 12529 9673 12541 9676
rect 12575 9673 12587 9707
rect 12529 9667 12587 9673
rect 14458 9664 14464 9716
rect 14516 9664 14522 9716
rect 15010 9704 15016 9716
rect 14568 9676 15016 9704
rect 9493 9639 9551 9645
rect 9493 9636 9505 9639
rect 9416 9608 9505 9636
rect 9493 9605 9505 9608
rect 9539 9605 9551 9639
rect 9493 9599 9551 9605
rect 9677 9639 9735 9645
rect 9677 9605 9689 9639
rect 9723 9636 9735 9639
rect 9723 9608 9904 9636
rect 9723 9605 9735 9608
rect 9677 9599 9735 9605
rect 8113 9571 8171 9577
rect 8113 9537 8125 9571
rect 8159 9537 8171 9571
rect 8113 9531 8171 9537
rect 8369 9571 8427 9577
rect 8369 9537 8381 9571
rect 8415 9568 8427 9571
rect 8415 9537 8432 9568
rect 8369 9531 8432 9537
rect 7024 9500 7052 9528
rect 8128 9500 8156 9531
rect 7024 9472 8156 9500
rect 8404 9500 8432 9531
rect 9122 9528 9128 9580
rect 9180 9528 9186 9580
rect 9398 9528 9404 9580
rect 9456 9528 9462 9580
rect 9769 9571 9827 9577
rect 9769 9537 9781 9571
rect 9815 9537 9827 9571
rect 9769 9531 9827 9537
rect 9784 9500 9812 9531
rect 8404 9472 9812 9500
rect 8404 9444 8432 9472
rect 8386 9392 8392 9444
rect 8444 9392 8450 9444
rect 8478 9392 8484 9444
rect 8536 9432 8542 9444
rect 9876 9432 9904 9608
rect 10226 9596 10232 9648
rect 10284 9636 10290 9648
rect 10689 9639 10747 9645
rect 10689 9636 10701 9639
rect 10284 9608 10701 9636
rect 10284 9596 10290 9608
rect 10689 9605 10701 9608
rect 10735 9636 10747 9639
rect 10962 9636 10968 9648
rect 10735 9608 10968 9636
rect 10735 9605 10747 9608
rect 10689 9599 10747 9605
rect 10962 9596 10968 9608
rect 11020 9596 11026 9648
rect 11885 9639 11943 9645
rect 11885 9605 11897 9639
rect 11931 9636 11943 9639
rect 11931 9608 12204 9636
rect 11931 9605 11943 9608
rect 11885 9599 11943 9605
rect 11054 9528 11060 9580
rect 11112 9528 11118 9580
rect 11146 9528 11152 9580
rect 11204 9568 11210 9580
rect 11422 9568 11428 9580
rect 11204 9540 11428 9568
rect 11204 9528 11210 9540
rect 11422 9528 11428 9540
rect 11480 9528 11486 9580
rect 11698 9528 11704 9580
rect 11756 9528 11762 9580
rect 11977 9571 12035 9577
rect 11977 9537 11989 9571
rect 12023 9537 12035 9571
rect 12176 9568 12204 9608
rect 12250 9596 12256 9648
rect 12308 9636 12314 9648
rect 14568 9645 14596 9676
rect 15010 9664 15016 9676
rect 15068 9664 15074 9716
rect 15378 9664 15384 9716
rect 15436 9704 15442 9716
rect 15657 9707 15715 9713
rect 15657 9704 15669 9707
rect 15436 9676 15669 9704
rect 15436 9664 15442 9676
rect 15657 9673 15669 9676
rect 15703 9673 15715 9707
rect 15657 9667 15715 9673
rect 22370 9664 22376 9716
rect 22428 9704 22434 9716
rect 22649 9707 22707 9713
rect 22649 9704 22661 9707
rect 22428 9676 22661 9704
rect 22428 9664 22434 9676
rect 22649 9673 22661 9676
rect 22695 9673 22707 9707
rect 22649 9667 22707 9673
rect 24118 9664 24124 9716
rect 24176 9704 24182 9716
rect 24305 9707 24363 9713
rect 24305 9704 24317 9707
rect 24176 9676 24317 9704
rect 24176 9664 24182 9676
rect 24305 9673 24317 9676
rect 24351 9673 24363 9707
rect 24305 9667 24363 9673
rect 24964 9676 25268 9704
rect 12437 9639 12495 9645
rect 12437 9636 12449 9639
rect 12308 9608 12449 9636
rect 12308 9596 12314 9608
rect 12437 9605 12449 9608
rect 12483 9605 12495 9639
rect 14553 9639 14611 9645
rect 14553 9636 14565 9639
rect 12437 9599 12495 9605
rect 12728 9608 13400 9636
rect 14531 9608 14565 9636
rect 12728 9568 12756 9608
rect 12176 9540 12756 9568
rect 11977 9531 12035 9537
rect 10778 9460 10784 9512
rect 10836 9460 10842 9512
rect 11992 9500 12020 9531
rect 12802 9528 12808 9580
rect 12860 9568 12866 9580
rect 13265 9571 13323 9577
rect 13265 9568 13277 9571
rect 12860 9540 13277 9568
rect 12860 9528 12866 9540
rect 13265 9537 13277 9540
rect 13311 9537 13323 9571
rect 13265 9531 13323 9537
rect 11348 9472 12020 9500
rect 12345 9503 12403 9509
rect 11348 9441 11376 9472
rect 12345 9469 12357 9503
rect 12391 9469 12403 9503
rect 12710 9500 12716 9512
rect 12345 9463 12403 9469
rect 12452 9472 12716 9500
rect 8536 9404 9904 9432
rect 11333 9435 11391 9441
rect 8536 9392 8542 9404
rect 11333 9401 11345 9435
rect 11379 9401 11391 9435
rect 11333 9395 11391 9401
rect 11422 9392 11428 9444
rect 11480 9432 11486 9444
rect 12250 9432 12256 9444
rect 11480 9404 12256 9432
rect 11480 9392 11486 9404
rect 12250 9392 12256 9404
rect 12308 9392 12314 9444
rect 12360 9432 12388 9463
rect 12452 9432 12480 9472
rect 12710 9460 12716 9472
rect 12768 9460 12774 9512
rect 13170 9460 13176 9512
rect 13228 9460 13234 9512
rect 13372 9509 13400 9608
rect 14553 9605 14565 9608
rect 14599 9605 14611 9639
rect 14753 9639 14811 9645
rect 14753 9636 14765 9639
rect 14553 9599 14611 9605
rect 14660 9608 14765 9636
rect 13446 9528 13452 9580
rect 13504 9528 13510 9580
rect 14277 9571 14335 9577
rect 14277 9537 14289 9571
rect 14323 9568 14335 9571
rect 14366 9568 14372 9580
rect 14323 9540 14372 9568
rect 14323 9537 14335 9540
rect 14277 9531 14335 9537
rect 13357 9503 13415 9509
rect 13357 9469 13369 9503
rect 13403 9500 13415 9503
rect 14292 9500 14320 9531
rect 14366 9528 14372 9540
rect 14424 9528 14430 9580
rect 14461 9571 14519 9577
rect 14461 9537 14473 9571
rect 14507 9568 14519 9571
rect 14507 9540 14596 9568
rect 14507 9537 14519 9540
rect 14461 9531 14519 9537
rect 14568 9512 14596 9540
rect 13403 9472 14320 9500
rect 13403 9469 13415 9472
rect 13357 9463 13415 9469
rect 14550 9460 14556 9512
rect 14608 9460 14614 9512
rect 12989 9435 13047 9441
rect 12989 9432 13001 9435
rect 12360 9404 12480 9432
rect 12728 9404 13001 9432
rect 7098 9324 7104 9376
rect 7156 9364 7162 9376
rect 7377 9367 7435 9373
rect 7377 9364 7389 9367
rect 7156 9336 7389 9364
rect 7156 9324 7162 9336
rect 7377 9333 7389 9336
rect 7423 9364 7435 9367
rect 7558 9364 7564 9376
rect 7423 9336 7564 9364
rect 7423 9333 7435 9336
rect 7377 9327 7435 9333
rect 7558 9324 7564 9336
rect 7616 9324 7622 9376
rect 8573 9367 8631 9373
rect 8573 9333 8585 9367
rect 8619 9364 8631 9367
rect 8938 9364 8944 9376
rect 8619 9336 8944 9364
rect 8619 9333 8631 9336
rect 8573 9327 8631 9333
rect 8938 9324 8944 9336
rect 8996 9324 9002 9376
rect 9030 9324 9036 9376
rect 9088 9364 9094 9376
rect 9585 9367 9643 9373
rect 9585 9364 9597 9367
rect 9088 9336 9597 9364
rect 9088 9324 9094 9336
rect 9585 9333 9597 9336
rect 9631 9333 9643 9367
rect 9585 9327 9643 9333
rect 10870 9324 10876 9376
rect 10928 9364 10934 9376
rect 11517 9367 11575 9373
rect 11517 9364 11529 9367
rect 10928 9336 11529 9364
rect 10928 9324 10934 9336
rect 11517 9333 11529 9336
rect 11563 9333 11575 9367
rect 11517 9327 11575 9333
rect 11606 9324 11612 9376
rect 11664 9364 11670 9376
rect 12728 9364 12756 9404
rect 12989 9401 13001 9404
rect 13035 9401 13047 9435
rect 14660 9432 14688 9608
rect 14753 9605 14765 9608
rect 14799 9605 14811 9639
rect 16209 9639 16267 9645
rect 16209 9636 16221 9639
rect 14753 9599 14811 9605
rect 15212 9608 16221 9636
rect 15212 9577 15240 9608
rect 16209 9605 16221 9608
rect 16255 9605 16267 9639
rect 16209 9599 16267 9605
rect 19058 9596 19064 9648
rect 19116 9636 19122 9648
rect 22554 9636 22560 9648
rect 19116 9608 21956 9636
rect 19116 9596 19122 9608
rect 15105 9571 15163 9577
rect 15105 9568 15117 9571
rect 14936 9540 15117 9568
rect 14936 9441 14964 9540
rect 15105 9537 15117 9540
rect 15151 9537 15163 9571
rect 15105 9531 15163 9537
rect 15197 9571 15255 9577
rect 15197 9537 15209 9571
rect 15243 9537 15255 9571
rect 15197 9531 15255 9537
rect 15378 9528 15384 9580
rect 15436 9528 15442 9580
rect 15473 9571 15531 9577
rect 15473 9537 15485 9571
rect 15519 9568 15531 9571
rect 15838 9568 15844 9580
rect 15519 9540 15844 9568
rect 15519 9537 15531 9540
rect 15473 9531 15531 9537
rect 15838 9528 15844 9540
rect 15896 9528 15902 9580
rect 15930 9528 15936 9580
rect 15988 9528 15994 9580
rect 16025 9571 16083 9577
rect 16025 9537 16037 9571
rect 16071 9568 16083 9571
rect 17034 9568 17040 9580
rect 16071 9540 17040 9568
rect 16071 9537 16083 9540
rect 16025 9531 16083 9537
rect 17034 9528 17040 9540
rect 17092 9528 17098 9580
rect 17770 9528 17776 9580
rect 17828 9568 17834 9580
rect 18141 9571 18199 9577
rect 18141 9568 18153 9571
rect 17828 9540 18153 9568
rect 17828 9528 17834 9540
rect 18141 9537 18153 9540
rect 18187 9537 18199 9571
rect 18141 9531 18199 9537
rect 18325 9571 18383 9577
rect 18325 9537 18337 9571
rect 18371 9568 18383 9571
rect 19242 9568 19248 9580
rect 18371 9540 19248 9568
rect 18371 9537 18383 9540
rect 18325 9531 18383 9537
rect 19242 9528 19248 9540
rect 19300 9528 19306 9580
rect 19334 9528 19340 9580
rect 19392 9568 19398 9580
rect 20530 9568 20536 9580
rect 19392 9540 20536 9568
rect 19392 9528 19398 9540
rect 20530 9528 20536 9540
rect 20588 9528 20594 9580
rect 20717 9571 20775 9577
rect 20717 9537 20729 9571
rect 20763 9568 20775 9571
rect 20806 9568 20812 9580
rect 20763 9540 20812 9568
rect 20763 9537 20775 9540
rect 20717 9531 20775 9537
rect 20806 9528 20812 9540
rect 20864 9528 20870 9580
rect 16209 9503 16267 9509
rect 16209 9469 16221 9503
rect 16255 9500 16267 9503
rect 17494 9500 17500 9512
rect 16255 9472 17500 9500
rect 16255 9469 16267 9472
rect 16209 9463 16267 9469
rect 17494 9460 17500 9472
rect 17552 9460 17558 9512
rect 18417 9503 18475 9509
rect 18417 9469 18429 9503
rect 18463 9469 18475 9503
rect 18417 9463 18475 9469
rect 12989 9395 13047 9401
rect 13832 9404 14688 9432
rect 14921 9435 14979 9441
rect 11664 9336 12756 9364
rect 12897 9367 12955 9373
rect 11664 9324 11670 9336
rect 12897 9333 12909 9367
rect 12943 9364 12955 9367
rect 13832 9364 13860 9404
rect 14921 9401 14933 9435
rect 14967 9401 14979 9435
rect 14921 9395 14979 9401
rect 15010 9392 15016 9444
rect 15068 9432 15074 9444
rect 15930 9432 15936 9444
rect 15068 9404 15936 9432
rect 15068 9392 15074 9404
rect 15930 9392 15936 9404
rect 15988 9392 15994 9444
rect 18432 9432 18460 9463
rect 18690 9460 18696 9512
rect 18748 9500 18754 9512
rect 21174 9500 21180 9512
rect 18748 9472 21180 9500
rect 18748 9460 18754 9472
rect 21174 9460 21180 9472
rect 21232 9460 21238 9512
rect 19334 9432 19340 9444
rect 18432 9404 19340 9432
rect 19334 9392 19340 9404
rect 19392 9392 19398 9444
rect 21928 9432 21956 9608
rect 22112 9608 22560 9636
rect 22112 9577 22140 9608
rect 22554 9596 22560 9608
rect 22612 9596 22618 9648
rect 23106 9596 23112 9648
rect 23164 9636 23170 9648
rect 24964 9645 24992 9676
rect 24949 9639 25007 9645
rect 23164 9608 24256 9636
rect 23164 9596 23170 9608
rect 22097 9571 22155 9577
rect 22097 9537 22109 9571
rect 22143 9537 22155 9571
rect 22097 9531 22155 9537
rect 22002 9460 22008 9512
rect 22060 9500 22066 9512
rect 22112 9500 22140 9531
rect 22278 9528 22284 9580
rect 22336 9568 22342 9580
rect 22373 9571 22431 9577
rect 22373 9568 22385 9571
rect 22336 9540 22385 9568
rect 22336 9528 22342 9540
rect 22373 9537 22385 9540
rect 22419 9568 22431 9571
rect 22833 9571 22891 9577
rect 22833 9568 22845 9571
rect 22419 9540 22845 9568
rect 22419 9537 22431 9540
rect 22373 9531 22431 9537
rect 22833 9537 22845 9540
rect 22879 9537 22891 9571
rect 22833 9531 22891 9537
rect 23017 9571 23075 9577
rect 23017 9537 23029 9571
rect 23063 9537 23075 9571
rect 23017 9531 23075 9537
rect 22060 9472 22140 9500
rect 22060 9460 22066 9472
rect 22186 9460 22192 9512
rect 22244 9460 22250 9512
rect 23032 9500 23060 9531
rect 23934 9528 23940 9580
rect 23992 9568 23998 9580
rect 24121 9571 24179 9577
rect 24121 9568 24133 9571
rect 23992 9540 24133 9568
rect 23992 9528 23998 9540
rect 24121 9537 24133 9540
rect 24167 9537 24179 9571
rect 24228 9568 24256 9608
rect 24949 9605 24961 9639
rect 24995 9605 25007 9639
rect 25149 9639 25207 9645
rect 25149 9636 25161 9639
rect 24949 9599 25007 9605
rect 25148 9605 25161 9636
rect 25195 9605 25207 9639
rect 25240 9636 25268 9676
rect 25314 9664 25320 9716
rect 25372 9664 25378 9716
rect 28626 9664 28632 9716
rect 28684 9664 28690 9716
rect 30742 9664 30748 9716
rect 30800 9704 30806 9716
rect 30837 9707 30895 9713
rect 30837 9704 30849 9707
rect 30800 9676 30849 9704
rect 30800 9664 30806 9676
rect 30837 9673 30849 9676
rect 30883 9673 30895 9707
rect 30837 9667 30895 9673
rect 34422 9664 34428 9716
rect 34480 9704 34486 9716
rect 34885 9707 34943 9713
rect 34480 9676 34744 9704
rect 34480 9664 34486 9676
rect 25590 9636 25596 9648
rect 25240 9608 25596 9636
rect 25148 9599 25207 9605
rect 25148 9568 25176 9599
rect 25590 9596 25596 9608
rect 25648 9596 25654 9648
rect 26786 9596 26792 9648
rect 26844 9636 26850 9648
rect 26973 9639 27031 9645
rect 26973 9636 26985 9639
rect 26844 9608 26985 9636
rect 26844 9596 26850 9608
rect 26973 9605 26985 9608
rect 27019 9605 27031 9639
rect 26973 9599 27031 9605
rect 27062 9596 27068 9648
rect 27120 9636 27126 9648
rect 27890 9636 27896 9648
rect 27120 9608 27896 9636
rect 27120 9596 27126 9608
rect 27890 9596 27896 9608
rect 27948 9596 27954 9648
rect 29086 9596 29092 9648
rect 29144 9636 29150 9648
rect 29181 9639 29239 9645
rect 29181 9636 29193 9639
rect 29144 9608 29193 9636
rect 29144 9596 29150 9608
rect 29181 9605 29193 9608
rect 29227 9605 29239 9639
rect 29181 9599 29239 9605
rect 29822 9596 29828 9648
rect 29880 9596 29886 9648
rect 30926 9636 30932 9648
rect 30300 9608 30932 9636
rect 24228 9540 25268 9568
rect 24121 9531 24179 9537
rect 25130 9500 25136 9512
rect 22296 9472 22968 9500
rect 23032 9472 25136 9500
rect 22296 9432 22324 9472
rect 22940 9432 22968 9472
rect 25130 9460 25136 9472
rect 25188 9460 25194 9512
rect 25240 9500 25268 9540
rect 26878 9528 26884 9580
rect 26936 9568 26942 9580
rect 27430 9568 27436 9580
rect 26936 9540 27436 9568
rect 26936 9528 26942 9540
rect 27430 9528 27436 9540
rect 27488 9568 27494 9580
rect 27801 9571 27859 9577
rect 27801 9568 27813 9571
rect 27488 9540 27813 9568
rect 27488 9528 27494 9540
rect 27801 9537 27813 9540
rect 27847 9568 27859 9571
rect 28442 9568 28448 9580
rect 27847 9540 28448 9568
rect 27847 9537 27859 9540
rect 27801 9531 27859 9537
rect 28442 9528 28448 9540
rect 28500 9528 28506 9580
rect 28813 9571 28871 9577
rect 28813 9537 28825 9571
rect 28859 9537 28871 9571
rect 28813 9531 28871 9537
rect 25682 9500 25688 9512
rect 25240 9472 25688 9500
rect 25682 9460 25688 9472
rect 25740 9460 25746 9512
rect 26418 9460 26424 9512
rect 26476 9500 26482 9512
rect 27062 9500 27068 9512
rect 26476 9472 27068 9500
rect 26476 9460 26482 9472
rect 27062 9460 27068 9472
rect 27120 9460 27126 9512
rect 27338 9460 27344 9512
rect 27396 9460 27402 9512
rect 27890 9460 27896 9512
rect 27948 9460 27954 9512
rect 28828 9500 28856 9531
rect 29822 9500 29828 9512
rect 28828 9472 29828 9500
rect 29822 9460 29828 9472
rect 29880 9460 29886 9512
rect 30193 9503 30251 9509
rect 30193 9469 30205 9503
rect 30239 9500 30251 9503
rect 30300 9500 30328 9608
rect 30926 9596 30932 9608
rect 30984 9636 30990 9648
rect 31386 9636 31392 9648
rect 30984 9608 31392 9636
rect 30984 9596 30990 9608
rect 31386 9596 31392 9608
rect 31444 9596 31450 9648
rect 34609 9639 34667 9645
rect 34609 9636 34621 9639
rect 31726 9608 34621 9636
rect 30374 9528 30380 9580
rect 30432 9568 30438 9580
rect 31018 9568 31024 9580
rect 30432 9540 31024 9568
rect 30432 9528 30438 9540
rect 31018 9528 31024 9540
rect 31076 9528 31082 9580
rect 31113 9571 31171 9577
rect 31113 9537 31125 9571
rect 31159 9537 31171 9571
rect 31113 9531 31171 9537
rect 31205 9571 31263 9577
rect 31205 9537 31217 9571
rect 31251 9537 31263 9571
rect 31205 9531 31263 9537
rect 31128 9500 31156 9531
rect 30239 9472 30328 9500
rect 30668 9472 31156 9500
rect 30239 9469 30251 9472
rect 30193 9463 30251 9469
rect 30098 9432 30104 9444
rect 20640 9404 21036 9432
rect 21928 9404 22324 9432
rect 22388 9404 22876 9432
rect 22940 9404 30104 9432
rect 12943 9336 13860 9364
rect 12943 9333 12955 9336
rect 12897 9327 12955 9333
rect 14458 9324 14464 9376
rect 14516 9364 14522 9376
rect 14737 9367 14795 9373
rect 14737 9364 14749 9367
rect 14516 9336 14749 9364
rect 14516 9324 14522 9336
rect 14737 9333 14749 9336
rect 14783 9333 14795 9367
rect 14737 9327 14795 9333
rect 15838 9324 15844 9376
rect 15896 9364 15902 9376
rect 17586 9364 17592 9376
rect 15896 9336 17592 9364
rect 15896 9324 15902 9336
rect 17586 9324 17592 9336
rect 17644 9364 17650 9376
rect 17957 9367 18015 9373
rect 17957 9364 17969 9367
rect 17644 9336 17969 9364
rect 17644 9324 17650 9336
rect 17957 9333 17969 9336
rect 18003 9333 18015 9367
rect 17957 9327 18015 9333
rect 20346 9324 20352 9376
rect 20404 9364 20410 9376
rect 20640 9373 20668 9404
rect 20625 9367 20683 9373
rect 20625 9364 20637 9367
rect 20404 9336 20637 9364
rect 20404 9324 20410 9336
rect 20625 9333 20637 9336
rect 20671 9333 20683 9367
rect 20625 9327 20683 9333
rect 20898 9324 20904 9376
rect 20956 9324 20962 9376
rect 21008 9364 21036 9404
rect 22388 9373 22416 9404
rect 22373 9367 22431 9373
rect 22373 9364 22385 9367
rect 21008 9336 22385 9364
rect 22373 9333 22385 9336
rect 22419 9333 22431 9367
rect 22373 9327 22431 9333
rect 22554 9324 22560 9376
rect 22612 9324 22618 9376
rect 22848 9373 22876 9404
rect 30098 9392 30104 9404
rect 30156 9392 30162 9444
rect 30282 9392 30288 9444
rect 30340 9432 30346 9444
rect 30668 9432 30696 9472
rect 30340 9404 30696 9432
rect 30340 9392 30346 9404
rect 30742 9392 30748 9444
rect 30800 9432 30806 9444
rect 31220 9432 31248 9531
rect 30800 9404 31248 9432
rect 30800 9392 30806 9404
rect 22833 9367 22891 9373
rect 22833 9333 22845 9367
rect 22879 9333 22891 9367
rect 22833 9327 22891 9333
rect 25133 9367 25191 9373
rect 25133 9333 25145 9367
rect 25179 9364 25191 9367
rect 25222 9364 25228 9376
rect 25179 9336 25228 9364
rect 25179 9333 25191 9336
rect 25133 9327 25191 9333
rect 25222 9324 25228 9336
rect 25280 9324 25286 9376
rect 25406 9324 25412 9376
rect 25464 9364 25470 9376
rect 25958 9364 25964 9376
rect 25464 9336 25964 9364
rect 25464 9324 25470 9336
rect 25958 9324 25964 9336
rect 26016 9364 26022 9376
rect 26234 9364 26240 9376
rect 26016 9336 26240 9364
rect 26016 9324 26022 9336
rect 26234 9324 26240 9336
rect 26292 9324 26298 9376
rect 27433 9367 27491 9373
rect 27433 9333 27445 9367
rect 27479 9364 27491 9367
rect 27614 9364 27620 9376
rect 27479 9336 27620 9364
rect 27479 9333 27491 9336
rect 27433 9327 27491 9333
rect 27614 9324 27620 9336
rect 27672 9364 27678 9376
rect 27798 9364 27804 9376
rect 27672 9336 27804 9364
rect 27672 9324 27678 9336
rect 27798 9324 27804 9336
rect 27856 9364 27862 9376
rect 28626 9364 28632 9376
rect 27856 9336 28632 9364
rect 27856 9324 27862 9336
rect 28626 9324 28632 9336
rect 28684 9324 28690 9376
rect 28994 9324 29000 9376
rect 29052 9364 29058 9376
rect 29089 9367 29147 9373
rect 29089 9364 29101 9367
rect 29052 9336 29101 9364
rect 29052 9324 29058 9336
rect 29089 9333 29101 9336
rect 29135 9333 29147 9367
rect 29089 9327 29147 9333
rect 30374 9324 30380 9376
rect 30432 9324 30438 9376
rect 30466 9324 30472 9376
rect 30524 9364 30530 9376
rect 31726 9364 31754 9608
rect 34609 9605 34621 9608
rect 34655 9605 34667 9639
rect 34716 9636 34744 9676
rect 34885 9673 34897 9707
rect 34931 9704 34943 9707
rect 35342 9704 35348 9716
rect 34931 9676 35348 9704
rect 34931 9673 34943 9676
rect 34885 9667 34943 9673
rect 35342 9664 35348 9676
rect 35400 9664 35406 9716
rect 36262 9704 36268 9716
rect 35820 9676 36268 9704
rect 35207 9639 35265 9645
rect 35207 9636 35219 9639
rect 34716 9608 35219 9636
rect 34609 9599 34667 9605
rect 35207 9605 35219 9608
rect 35253 9605 35265 9639
rect 35207 9599 35265 9605
rect 35437 9639 35495 9645
rect 35437 9605 35449 9639
rect 35483 9636 35495 9639
rect 35618 9636 35624 9648
rect 35483 9608 35624 9636
rect 35483 9605 35495 9608
rect 35437 9599 35495 9605
rect 35618 9596 35624 9608
rect 35676 9596 35682 9648
rect 35713 9639 35771 9645
rect 35713 9605 35725 9639
rect 35759 9636 35771 9639
rect 35820 9636 35848 9676
rect 36262 9664 36268 9676
rect 36320 9664 36326 9716
rect 36630 9664 36636 9716
rect 36688 9704 36694 9716
rect 36725 9707 36783 9713
rect 36725 9704 36737 9707
rect 36688 9676 36737 9704
rect 36688 9664 36694 9676
rect 36725 9673 36737 9676
rect 36771 9673 36783 9707
rect 36725 9667 36783 9673
rect 35759 9608 35848 9636
rect 35759 9605 35771 9608
rect 35713 9599 35771 9605
rect 36078 9596 36084 9648
rect 36136 9596 36142 9648
rect 36173 9639 36231 9645
rect 36173 9605 36185 9639
rect 36219 9605 36231 9639
rect 36173 9599 36231 9605
rect 32122 9528 32128 9580
rect 32180 9528 32186 9580
rect 32309 9571 32367 9577
rect 32309 9537 32321 9571
rect 32355 9537 32367 9571
rect 32309 9531 32367 9537
rect 32493 9571 32551 9577
rect 32493 9537 32505 9571
rect 32539 9568 32551 9571
rect 32582 9568 32588 9580
rect 32539 9540 32588 9568
rect 32539 9537 32551 9540
rect 32493 9531 32551 9537
rect 32324 9500 32352 9531
rect 32582 9528 32588 9540
rect 32640 9528 32646 9580
rect 32674 9528 32680 9580
rect 32732 9528 32738 9580
rect 32858 9528 32864 9580
rect 32916 9528 32922 9580
rect 33318 9528 33324 9580
rect 33376 9568 33382 9580
rect 33870 9568 33876 9580
rect 33376 9540 33876 9568
rect 33376 9528 33382 9540
rect 33870 9528 33876 9540
rect 33928 9528 33934 9580
rect 34146 9528 34152 9580
rect 34204 9568 34210 9580
rect 34241 9571 34299 9577
rect 34241 9568 34253 9571
rect 34204 9540 34253 9568
rect 34204 9528 34210 9540
rect 34241 9537 34253 9540
rect 34287 9537 34299 9571
rect 34241 9531 34299 9537
rect 34389 9571 34447 9577
rect 34389 9537 34401 9571
rect 34435 9568 34447 9571
rect 34435 9537 34468 9568
rect 34389 9531 34468 9537
rect 33594 9500 33600 9512
rect 32324 9472 33600 9500
rect 33594 9460 33600 9472
rect 33652 9460 33658 9512
rect 34440 9432 34468 9531
rect 34514 9528 34520 9580
rect 34572 9528 34578 9580
rect 34698 9528 34704 9580
rect 34756 9577 34762 9580
rect 34756 9568 34764 9577
rect 34756 9540 34801 9568
rect 34756 9531 34764 9540
rect 34756 9528 34762 9531
rect 34882 9528 34888 9580
rect 34940 9568 34946 9580
rect 35069 9571 35127 9577
rect 35069 9568 35081 9571
rect 34940 9540 35081 9568
rect 34940 9528 34946 9540
rect 35069 9537 35081 9540
rect 35115 9537 35127 9571
rect 35069 9531 35127 9537
rect 35084 9500 35112 9531
rect 35342 9528 35348 9580
rect 35400 9528 35406 9580
rect 35526 9528 35532 9580
rect 35584 9528 35590 9580
rect 35986 9577 35992 9580
rect 35963 9571 35992 9577
rect 35963 9537 35975 9571
rect 35963 9531 35992 9537
rect 35986 9528 35992 9531
rect 36044 9528 36050 9580
rect 36188 9568 36216 9599
rect 36446 9596 36452 9648
rect 36504 9636 36510 9648
rect 37734 9636 37740 9648
rect 36504 9608 37740 9636
rect 36504 9596 36510 9608
rect 37734 9596 37740 9608
rect 37792 9596 37798 9648
rect 38010 9596 38016 9648
rect 38068 9596 38074 9648
rect 38289 9639 38347 9645
rect 38289 9605 38301 9639
rect 38335 9636 38347 9639
rect 39942 9636 39948 9648
rect 38335 9608 39948 9636
rect 38335 9605 38347 9608
rect 38289 9599 38347 9605
rect 39942 9596 39948 9608
rect 40000 9596 40006 9648
rect 36096 9540 36216 9568
rect 35805 9503 35863 9509
rect 35805 9500 35817 9503
rect 35084 9472 35817 9500
rect 35805 9469 35817 9472
rect 35851 9469 35863 9503
rect 36096 9500 36124 9540
rect 36262 9528 36268 9580
rect 36320 9528 36326 9580
rect 36538 9528 36544 9580
rect 36596 9568 36602 9580
rect 36633 9571 36691 9577
rect 36633 9568 36645 9571
rect 36596 9540 36645 9568
rect 36596 9528 36602 9540
rect 36633 9537 36645 9540
rect 36679 9537 36691 9571
rect 36633 9531 36691 9537
rect 37642 9528 37648 9580
rect 37700 9528 37706 9580
rect 37829 9571 37887 9577
rect 37829 9537 37841 9571
rect 37875 9537 37887 9571
rect 37829 9531 37887 9537
rect 38657 9571 38715 9577
rect 38657 9537 38669 9571
rect 38703 9537 38715 9571
rect 38657 9531 38715 9537
rect 36354 9500 36360 9512
rect 36096 9472 36360 9500
rect 35805 9463 35863 9469
rect 36354 9460 36360 9472
rect 36412 9460 36418 9512
rect 36449 9503 36507 9509
rect 36449 9469 36461 9503
rect 36495 9500 36507 9503
rect 37182 9500 37188 9512
rect 36495 9472 37188 9500
rect 36495 9469 36507 9472
rect 36449 9463 36507 9469
rect 37182 9460 37188 9472
rect 37240 9460 37246 9512
rect 37844 9500 37872 9531
rect 37292 9472 37872 9500
rect 36170 9432 36176 9444
rect 34440 9404 36176 9432
rect 36170 9392 36176 9404
rect 36228 9392 36234 9444
rect 36262 9392 36268 9444
rect 36320 9432 36326 9444
rect 37292 9432 37320 9472
rect 36320 9404 37320 9432
rect 36320 9392 36326 9404
rect 30524 9336 31754 9364
rect 30524 9324 30530 9336
rect 34606 9324 34612 9376
rect 34664 9364 34670 9376
rect 35526 9364 35532 9376
rect 34664 9336 35532 9364
rect 34664 9324 34670 9336
rect 35526 9324 35532 9336
rect 35584 9364 35590 9376
rect 36372 9364 36400 9404
rect 37458 9392 37464 9444
rect 37516 9392 37522 9444
rect 37550 9392 37556 9444
rect 37608 9432 37614 9444
rect 38473 9435 38531 9441
rect 38473 9432 38485 9435
rect 37608 9404 38485 9432
rect 37608 9392 37614 9404
rect 38473 9401 38485 9404
rect 38519 9401 38531 9435
rect 38473 9395 38531 9401
rect 35584 9336 36400 9364
rect 35584 9324 35590 9336
rect 36814 9324 36820 9376
rect 36872 9364 36878 9376
rect 38197 9367 38255 9373
rect 38197 9364 38209 9367
rect 36872 9336 38209 9364
rect 36872 9324 36878 9336
rect 38197 9333 38209 9336
rect 38243 9364 38255 9367
rect 38672 9364 38700 9531
rect 38243 9336 38700 9364
rect 38243 9333 38255 9336
rect 38197 9327 38255 9333
rect 1104 9274 40572 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 40572 9274
rect 1104 9200 40572 9222
rect 9122 9160 9128 9172
rect 7668 9132 9128 9160
rect 7668 9092 7696 9132
rect 9122 9120 9128 9132
rect 9180 9160 9186 9172
rect 9858 9160 9864 9172
rect 9180 9132 9864 9160
rect 9180 9120 9186 9132
rect 9858 9120 9864 9132
rect 9916 9160 9922 9172
rect 10318 9160 10324 9172
rect 9916 9132 10324 9160
rect 9916 9120 9922 9132
rect 10318 9120 10324 9132
rect 10376 9120 10382 9172
rect 10686 9120 10692 9172
rect 10744 9160 10750 9172
rect 12805 9163 12863 9169
rect 10744 9132 11652 9160
rect 10744 9120 10750 9132
rect 7484 9064 7696 9092
rect 5258 8984 5264 9036
rect 5316 9024 5322 9036
rect 6822 9024 6828 9036
rect 5316 8996 6828 9024
rect 5316 8984 5322 8996
rect 6822 8984 6828 8996
rect 6880 9024 6886 9036
rect 7484 9024 7512 9064
rect 7742 9052 7748 9104
rect 7800 9092 7806 9104
rect 7929 9095 7987 9101
rect 7929 9092 7941 9095
rect 7800 9064 7941 9092
rect 7800 9052 7806 9064
rect 7929 9061 7941 9064
rect 7975 9061 7987 9095
rect 7929 9055 7987 9061
rect 8018 9052 8024 9104
rect 8076 9092 8082 9104
rect 8076 9064 9812 9092
rect 8076 9052 8082 9064
rect 8110 9024 8116 9036
rect 6880 8996 7512 9024
rect 6880 8984 6886 8996
rect 6917 8959 6975 8965
rect 6917 8925 6929 8959
rect 6963 8956 6975 8959
rect 7098 8956 7104 8968
rect 6963 8928 7104 8956
rect 6963 8925 6975 8928
rect 6917 8919 6975 8925
rect 7098 8916 7104 8928
rect 7156 8916 7162 8968
rect 7282 8916 7288 8968
rect 7340 8916 7346 8968
rect 7484 8965 7512 8996
rect 7760 8996 8116 9024
rect 7760 8965 7788 8996
rect 8110 8984 8116 8996
rect 8168 8984 8174 9036
rect 8938 9024 8944 9036
rect 8220 8996 8944 9024
rect 7469 8959 7527 8965
rect 7469 8925 7481 8959
rect 7515 8925 7527 8959
rect 7469 8919 7527 8925
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8925 7711 8959
rect 7653 8919 7711 8925
rect 7745 8959 7803 8965
rect 7745 8925 7757 8959
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 7006 8848 7012 8900
rect 7064 8848 7070 8900
rect 7193 8891 7251 8897
rect 7193 8857 7205 8891
rect 7239 8888 7251 8891
rect 7668 8888 7696 8919
rect 7834 8916 7840 8968
rect 7892 8956 7898 8968
rect 8220 8965 8248 8996
rect 8938 8984 8944 8996
rect 8996 8984 9002 9036
rect 8205 8959 8263 8965
rect 8205 8956 8217 8959
rect 7892 8928 8217 8956
rect 7892 8916 7898 8928
rect 8205 8925 8217 8928
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8956 8447 8959
rect 9030 8956 9036 8968
rect 8435 8928 9036 8956
rect 8435 8925 8447 8928
rect 8389 8919 8447 8925
rect 9030 8916 9036 8928
rect 9088 8916 9094 8968
rect 7929 8891 7987 8897
rect 7239 8860 7880 8888
rect 7239 8857 7251 8860
rect 7193 8851 7251 8857
rect 7484 8832 7512 8860
rect 6638 8780 6644 8832
rect 6696 8820 6702 8832
rect 6917 8823 6975 8829
rect 6917 8820 6929 8823
rect 6696 8792 6929 8820
rect 6696 8780 6702 8792
rect 6917 8789 6929 8792
rect 6963 8789 6975 8823
rect 6917 8783 6975 8789
rect 7098 8780 7104 8832
rect 7156 8820 7162 8832
rect 7377 8823 7435 8829
rect 7377 8820 7389 8823
rect 7156 8792 7389 8820
rect 7156 8780 7162 8792
rect 7377 8789 7389 8792
rect 7423 8789 7435 8823
rect 7377 8783 7435 8789
rect 7466 8780 7472 8832
rect 7524 8780 7530 8832
rect 7852 8820 7880 8860
rect 7929 8857 7941 8891
rect 7975 8888 7987 8891
rect 8297 8891 8355 8897
rect 8297 8888 8309 8891
rect 7975 8860 8309 8888
rect 7975 8857 7987 8860
rect 7929 8851 7987 8857
rect 8297 8857 8309 8860
rect 8343 8857 8355 8891
rect 9784 8888 9812 9064
rect 10778 9052 10784 9104
rect 10836 9092 10842 9104
rect 11624 9092 11652 9132
rect 12805 9129 12817 9163
rect 12851 9160 12863 9163
rect 13170 9160 13176 9172
rect 12851 9132 13176 9160
rect 12851 9129 12863 9132
rect 12805 9123 12863 9129
rect 13170 9120 13176 9132
rect 13228 9120 13234 9172
rect 20346 9120 20352 9172
rect 20404 9120 20410 9172
rect 20533 9163 20591 9169
rect 20533 9129 20545 9163
rect 20579 9160 20591 9163
rect 20990 9160 20996 9172
rect 20579 9132 20996 9160
rect 20579 9129 20591 9132
rect 20533 9123 20591 9129
rect 20990 9120 20996 9132
rect 21048 9120 21054 9172
rect 22186 9120 22192 9172
rect 22244 9160 22250 9172
rect 22281 9163 22339 9169
rect 22281 9160 22293 9163
rect 22244 9132 22293 9160
rect 22244 9120 22250 9132
rect 22281 9129 22293 9132
rect 22327 9129 22339 9163
rect 22281 9123 22339 9129
rect 22465 9163 22523 9169
rect 22465 9129 22477 9163
rect 22511 9129 22523 9163
rect 22465 9123 22523 9129
rect 12526 9092 12532 9104
rect 10836 9064 11560 9092
rect 11624 9064 11744 9092
rect 10836 9052 10842 9064
rect 11330 9024 11336 9036
rect 10704 8996 11336 9024
rect 10410 8916 10416 8968
rect 10468 8916 10474 8968
rect 10502 8916 10508 8968
rect 10560 8916 10566 8968
rect 10594 8916 10600 8968
rect 10652 8916 10658 8968
rect 10704 8965 10732 8996
rect 11330 8984 11336 8996
rect 11388 8984 11394 9036
rect 10689 8959 10747 8965
rect 10689 8925 10701 8959
rect 10735 8925 10747 8959
rect 10689 8919 10747 8925
rect 10873 8959 10931 8965
rect 10873 8925 10885 8959
rect 10919 8925 10931 8959
rect 10873 8919 10931 8925
rect 10428 8888 10456 8916
rect 10888 8888 10916 8919
rect 11146 8916 11152 8968
rect 11204 8916 11210 8968
rect 11422 8916 11428 8968
rect 11480 8916 11486 8968
rect 11532 8956 11560 9064
rect 11716 8965 11744 9064
rect 11808 9064 12532 9092
rect 11701 8959 11759 8965
rect 11532 8928 11652 8956
rect 9784 8860 10916 8888
rect 8297 8851 8355 8857
rect 11054 8848 11060 8900
rect 11112 8888 11118 8900
rect 11333 8891 11391 8897
rect 11333 8888 11345 8891
rect 11112 8860 11345 8888
rect 11112 8848 11118 8860
rect 11333 8857 11345 8860
rect 11379 8857 11391 8891
rect 11333 8851 11391 8857
rect 11517 8891 11575 8897
rect 11517 8857 11529 8891
rect 11563 8857 11575 8891
rect 11624 8888 11652 8928
rect 11701 8925 11713 8959
rect 11747 8925 11759 8959
rect 11701 8919 11759 8925
rect 11808 8888 11836 9064
rect 12526 9052 12532 9064
rect 12584 9052 12590 9104
rect 20806 9052 20812 9104
rect 20864 9092 20870 9104
rect 22480 9092 22508 9123
rect 23474 9120 23480 9172
rect 23532 9160 23538 9172
rect 24029 9163 24087 9169
rect 24029 9160 24041 9163
rect 23532 9132 24041 9160
rect 23532 9120 23538 9132
rect 24029 9129 24041 9132
rect 24075 9129 24087 9163
rect 24029 9123 24087 9129
rect 24578 9120 24584 9172
rect 24636 9120 24642 9172
rect 25038 9120 25044 9172
rect 25096 9160 25102 9172
rect 25096 9132 25268 9160
rect 25096 9120 25102 9132
rect 22554 9092 22560 9104
rect 20864 9064 22560 9092
rect 20864 9052 20870 9064
rect 22554 9052 22560 9064
rect 22612 9092 22618 9104
rect 24118 9092 24124 9104
rect 22612 9064 24124 9092
rect 22612 9052 22618 9064
rect 24118 9052 24124 9064
rect 24176 9052 24182 9104
rect 24596 9092 24624 9120
rect 25130 9092 25136 9104
rect 24596 9064 25136 9092
rect 25130 9052 25136 9064
rect 25188 9052 25194 9104
rect 25240 9092 25268 9132
rect 25314 9120 25320 9172
rect 25372 9160 25378 9172
rect 25501 9163 25559 9169
rect 25501 9160 25513 9163
rect 25372 9132 25513 9160
rect 25372 9120 25378 9132
rect 25501 9129 25513 9132
rect 25547 9160 25559 9163
rect 26142 9160 26148 9172
rect 25547 9132 26148 9160
rect 25547 9129 25559 9132
rect 25501 9123 25559 9129
rect 26142 9120 26148 9132
rect 26200 9120 26206 9172
rect 26234 9120 26240 9172
rect 26292 9160 26298 9172
rect 26513 9163 26571 9169
rect 26513 9160 26525 9163
rect 26292 9132 26525 9160
rect 26292 9120 26298 9132
rect 26513 9129 26525 9132
rect 26559 9129 26571 9163
rect 26513 9123 26571 9129
rect 26878 9120 26884 9172
rect 26936 9120 26942 9172
rect 26973 9163 27031 9169
rect 26973 9129 26985 9163
rect 27019 9160 27031 9163
rect 27614 9160 27620 9172
rect 27019 9132 27620 9160
rect 27019 9129 27031 9132
rect 26973 9123 27031 9129
rect 27614 9120 27620 9132
rect 27672 9120 27678 9172
rect 27706 9120 27712 9172
rect 27764 9120 27770 9172
rect 28350 9120 28356 9172
rect 28408 9160 28414 9172
rect 31110 9160 31116 9172
rect 28408 9132 31116 9160
rect 28408 9120 28414 9132
rect 31110 9120 31116 9132
rect 31168 9120 31174 9172
rect 31478 9120 31484 9172
rect 31536 9120 31542 9172
rect 33686 9160 33692 9172
rect 31726 9132 33692 9160
rect 28534 9092 28540 9104
rect 25240 9064 28540 9092
rect 28534 9052 28540 9064
rect 28592 9052 28598 9104
rect 28902 9052 28908 9104
rect 28960 9052 28966 9104
rect 30466 9092 30472 9104
rect 29012 9064 30472 9092
rect 11885 9027 11943 9033
rect 11885 8993 11897 9027
rect 11931 9024 11943 9027
rect 12710 9024 12716 9036
rect 11931 8996 12716 9024
rect 11931 8993 11943 8996
rect 11885 8987 11943 8993
rect 12161 8959 12219 8965
rect 12161 8925 12173 8959
rect 12207 8956 12219 8959
rect 12250 8956 12256 8968
rect 12207 8928 12256 8956
rect 12207 8925 12219 8928
rect 12161 8919 12219 8925
rect 12250 8916 12256 8928
rect 12308 8916 12314 8968
rect 12342 8916 12348 8968
rect 12400 8916 12406 8968
rect 12452 8965 12480 8996
rect 12710 8984 12716 8996
rect 12768 8984 12774 9036
rect 15470 9024 15476 9036
rect 14568 8996 15476 9024
rect 14568 8965 14596 8996
rect 15470 8984 15476 8996
rect 15528 8984 15534 9036
rect 17402 8984 17408 9036
rect 17460 9024 17466 9036
rect 18230 9024 18236 9036
rect 17460 8996 18236 9024
rect 17460 8984 17466 8996
rect 12437 8959 12495 8965
rect 12437 8925 12449 8959
rect 12483 8956 12495 8959
rect 14553 8959 14611 8965
rect 12483 8928 12517 8956
rect 12483 8925 12495 8928
rect 12437 8919 12495 8925
rect 14553 8925 14565 8959
rect 14599 8925 14611 8959
rect 14553 8919 14611 8925
rect 14642 8916 14648 8968
rect 14700 8956 14706 8968
rect 14737 8959 14795 8965
rect 14737 8956 14749 8959
rect 14700 8928 14749 8956
rect 14700 8916 14706 8928
rect 14737 8925 14749 8928
rect 14783 8956 14795 8959
rect 16482 8956 16488 8968
rect 14783 8928 16488 8956
rect 14783 8925 14795 8928
rect 14737 8919 14795 8925
rect 16482 8916 16488 8928
rect 16540 8916 16546 8968
rect 17880 8965 17908 8996
rect 18230 8984 18236 8996
rect 18288 9024 18294 9036
rect 26234 9024 26240 9036
rect 18288 8996 21220 9024
rect 18288 8984 18294 8996
rect 17681 8959 17739 8965
rect 17681 8925 17693 8959
rect 17727 8925 17739 8959
rect 17681 8919 17739 8925
rect 17865 8959 17923 8965
rect 17865 8925 17877 8959
rect 17911 8925 17923 8959
rect 17865 8919 17923 8925
rect 17957 8959 18015 8965
rect 17957 8925 17969 8959
rect 18003 8956 18015 8959
rect 18322 8956 18328 8968
rect 18003 8928 18328 8956
rect 18003 8925 18015 8928
rect 17957 8919 18015 8925
rect 11977 8891 12035 8897
rect 11977 8888 11989 8891
rect 11624 8860 11989 8888
rect 11517 8851 11575 8857
rect 11977 8857 11989 8860
rect 12023 8857 12035 8891
rect 11977 8851 12035 8857
rect 8386 8820 8392 8832
rect 7852 8792 8392 8820
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 10318 8780 10324 8832
rect 10376 8780 10382 8832
rect 10410 8780 10416 8832
rect 10468 8820 10474 8832
rect 10965 8823 11023 8829
rect 10965 8820 10977 8823
rect 10468 8792 10977 8820
rect 10468 8780 10474 8792
rect 10965 8789 10977 8792
rect 11011 8789 11023 8823
rect 10965 8783 11023 8789
rect 11146 8780 11152 8832
rect 11204 8820 11210 8832
rect 11532 8820 11560 8851
rect 12526 8848 12532 8900
rect 12584 8888 12590 8900
rect 12621 8891 12679 8897
rect 12621 8888 12633 8891
rect 12584 8860 12633 8888
rect 12584 8848 12590 8860
rect 12621 8857 12633 8860
rect 12667 8857 12679 8891
rect 17696 8888 17724 8919
rect 18322 8916 18328 8928
rect 18380 8916 18386 8968
rect 20640 8928 20852 8956
rect 17770 8888 17776 8900
rect 17696 8860 17776 8888
rect 12621 8851 12679 8857
rect 17770 8848 17776 8860
rect 17828 8888 17834 8900
rect 19610 8888 19616 8900
rect 17828 8860 19616 8888
rect 17828 8848 17834 8860
rect 19610 8848 19616 8860
rect 19668 8888 19674 8900
rect 20162 8888 20168 8900
rect 19668 8860 20168 8888
rect 19668 8848 19674 8860
rect 20162 8848 20168 8860
rect 20220 8848 20226 8900
rect 20254 8848 20260 8900
rect 20312 8888 20318 8900
rect 20501 8891 20559 8897
rect 20501 8888 20513 8891
rect 20312 8860 20513 8888
rect 20312 8848 20318 8860
rect 20501 8857 20513 8860
rect 20547 8888 20559 8891
rect 20640 8888 20668 8928
rect 20547 8860 20668 8888
rect 20547 8857 20559 8860
rect 20501 8851 20559 8857
rect 20714 8848 20720 8900
rect 20772 8848 20778 8900
rect 20824 8888 20852 8928
rect 21192 8897 21220 8996
rect 25056 8996 26240 9024
rect 25056 8968 25084 8996
rect 26234 8984 26240 8996
rect 26292 8984 26298 9036
rect 26418 8984 26424 9036
rect 26476 9024 26482 9036
rect 26789 9027 26847 9033
rect 26789 9024 26801 9027
rect 26476 8996 26801 9024
rect 26476 8984 26482 8996
rect 26789 8993 26801 8996
rect 26835 9024 26847 9027
rect 27522 9024 27528 9036
rect 26835 8996 27528 9024
rect 26835 8993 26847 8996
rect 26789 8987 26847 8993
rect 27522 8984 27528 8996
rect 27580 9024 27586 9036
rect 29012 9024 29040 9064
rect 30466 9052 30472 9064
rect 30524 9052 30530 9104
rect 30558 9052 30564 9104
rect 30616 9092 30622 9104
rect 31726 9092 31754 9132
rect 33686 9120 33692 9132
rect 33744 9120 33750 9172
rect 35342 9120 35348 9172
rect 35400 9160 35406 9172
rect 35529 9163 35587 9169
rect 35529 9160 35541 9163
rect 35400 9132 35541 9160
rect 35400 9120 35406 9132
rect 35529 9129 35541 9132
rect 35575 9129 35587 9163
rect 35529 9123 35587 9129
rect 37369 9163 37427 9169
rect 37369 9129 37381 9163
rect 37415 9160 37427 9163
rect 37642 9160 37648 9172
rect 37415 9132 37648 9160
rect 37415 9129 37427 9132
rect 37369 9123 37427 9129
rect 37642 9120 37648 9132
rect 37700 9120 37706 9172
rect 37829 9163 37887 9169
rect 37829 9129 37841 9163
rect 37875 9160 37887 9163
rect 38010 9160 38016 9172
rect 37875 9132 38016 9160
rect 37875 9129 37887 9132
rect 37829 9123 37887 9129
rect 38010 9120 38016 9132
rect 38068 9120 38074 9172
rect 30616 9064 31754 9092
rect 30616 9052 30622 9064
rect 27580 8996 27660 9024
rect 27580 8984 27586 8996
rect 23106 8956 23112 8968
rect 22066 8928 23112 8956
rect 20961 8891 21019 8897
rect 20961 8888 20973 8891
rect 20824 8860 20973 8888
rect 20961 8857 20973 8860
rect 21007 8888 21019 8891
rect 21177 8891 21235 8897
rect 21007 8860 21128 8888
rect 21007 8857 21019 8860
rect 20961 8851 21019 8857
rect 11204 8792 11560 8820
rect 11204 8780 11210 8792
rect 11882 8780 11888 8832
rect 11940 8820 11946 8832
rect 12250 8820 12256 8832
rect 11940 8792 12256 8820
rect 11940 8780 11946 8792
rect 12250 8780 12256 8792
rect 12308 8820 12314 8832
rect 15378 8820 15384 8832
rect 12308 8792 15384 8820
rect 12308 8780 12314 8792
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 19978 8780 19984 8832
rect 20036 8820 20042 8832
rect 20622 8820 20628 8832
rect 20036 8792 20628 8820
rect 20036 8780 20042 8792
rect 20622 8780 20628 8792
rect 20680 8820 20686 8832
rect 20809 8823 20867 8829
rect 20809 8820 20821 8823
rect 20680 8792 20821 8820
rect 20680 8780 20686 8792
rect 20809 8789 20821 8792
rect 20855 8789 20867 8823
rect 21100 8820 21128 8860
rect 21177 8857 21189 8891
rect 21223 8857 21235 8891
rect 21177 8851 21235 8857
rect 22066 8820 22094 8928
rect 23106 8916 23112 8928
rect 23164 8916 23170 8968
rect 24210 8916 24216 8968
rect 24268 8916 24274 8968
rect 24762 8916 24768 8968
rect 24820 8916 24826 8968
rect 25038 8916 25044 8968
rect 25096 8916 25102 8968
rect 25406 8956 25412 8968
rect 25240 8928 25412 8956
rect 22649 8891 22707 8897
rect 22649 8857 22661 8891
rect 22695 8888 22707 8891
rect 22738 8888 22744 8900
rect 22695 8860 22744 8888
rect 22695 8857 22707 8860
rect 22649 8851 22707 8857
rect 22738 8848 22744 8860
rect 22796 8888 22802 8900
rect 23014 8888 23020 8900
rect 22796 8860 23020 8888
rect 22796 8848 22802 8860
rect 23014 8848 23020 8860
rect 23072 8848 23078 8900
rect 24394 8848 24400 8900
rect 24452 8848 24458 8900
rect 24613 8891 24671 8897
rect 24613 8888 24625 8891
rect 24504 8860 24625 8888
rect 21100 8792 22094 8820
rect 22449 8823 22507 8829
rect 20809 8783 20867 8789
rect 22449 8789 22461 8823
rect 22495 8820 22507 8823
rect 22922 8820 22928 8832
rect 22495 8792 22928 8820
rect 22495 8789 22507 8792
rect 22449 8783 22507 8789
rect 22922 8780 22928 8792
rect 22980 8780 22986 8832
rect 24026 8780 24032 8832
rect 24084 8820 24090 8832
rect 24504 8820 24532 8860
rect 24613 8857 24625 8860
rect 24659 8888 24671 8891
rect 24780 8888 24808 8916
rect 24659 8860 24808 8888
rect 24857 8891 24915 8897
rect 24659 8857 24671 8860
rect 24613 8851 24671 8857
rect 24857 8857 24869 8891
rect 24903 8888 24915 8891
rect 25056 8888 25084 8916
rect 25240 8888 25268 8928
rect 25406 8916 25412 8928
rect 25464 8916 25470 8968
rect 26050 8916 26056 8968
rect 26108 8956 26114 8968
rect 26145 8959 26203 8965
rect 26145 8956 26157 8959
rect 26108 8928 26157 8956
rect 26108 8916 26114 8928
rect 26145 8925 26157 8928
rect 26191 8925 26203 8959
rect 26145 8919 26203 8925
rect 26326 8916 26332 8968
rect 26384 8956 26390 8968
rect 27062 8956 27068 8968
rect 26384 8928 27068 8956
rect 26384 8916 26390 8928
rect 27062 8916 27068 8928
rect 27120 8916 27126 8968
rect 27338 8916 27344 8968
rect 27396 8916 27402 8968
rect 27632 8965 27660 8996
rect 28092 8996 29040 9024
rect 29089 9027 29147 9033
rect 27617 8959 27675 8965
rect 27617 8925 27629 8959
rect 27663 8925 27675 8959
rect 27617 8919 27675 8925
rect 24903 8860 25084 8888
rect 25148 8860 25268 8888
rect 24903 8857 24915 8860
rect 24857 8851 24915 8857
rect 24084 8792 24532 8820
rect 24084 8780 24090 8792
rect 24762 8780 24768 8832
rect 24820 8780 24826 8832
rect 25062 8823 25120 8829
rect 25062 8789 25074 8823
rect 25108 8820 25120 8823
rect 25148 8820 25176 8860
rect 25314 8848 25320 8900
rect 25372 8848 25378 8900
rect 25533 8891 25591 8897
rect 25533 8857 25545 8891
rect 25579 8888 25591 8891
rect 26237 8891 26295 8897
rect 25579 8860 26188 8888
rect 25579 8857 25591 8860
rect 25533 8851 25591 8857
rect 25108 8792 25176 8820
rect 25108 8789 25120 8792
rect 25062 8783 25120 8789
rect 25222 8780 25228 8832
rect 25280 8780 25286 8832
rect 25682 8780 25688 8832
rect 25740 8780 25746 8832
rect 26160 8820 26188 8860
rect 26237 8857 26249 8891
rect 26283 8888 26295 8891
rect 26694 8888 26700 8900
rect 26283 8860 26700 8888
rect 26283 8857 26295 8860
rect 26237 8851 26295 8857
rect 26694 8848 26700 8860
rect 26752 8888 26758 8900
rect 28092 8888 28120 8996
rect 29089 8993 29101 9027
rect 29135 9024 29147 9027
rect 29178 9024 29184 9036
rect 29135 8996 29184 9024
rect 29135 8993 29147 8996
rect 29089 8987 29147 8993
rect 29178 8984 29184 8996
rect 29236 8984 29242 9036
rect 29288 8996 32352 9024
rect 28258 8916 28264 8968
rect 28316 8916 28322 8968
rect 28718 8916 28724 8968
rect 28776 8916 28782 8968
rect 29288 8965 29316 8996
rect 28997 8959 29055 8965
rect 28997 8925 29009 8959
rect 29043 8925 29055 8959
rect 28997 8919 29055 8925
rect 29273 8959 29331 8965
rect 29273 8925 29285 8959
rect 29319 8925 29331 8959
rect 29273 8919 29331 8925
rect 26752 8860 28120 8888
rect 26752 8848 26758 8860
rect 28626 8848 28632 8900
rect 28684 8888 28690 8900
rect 29012 8888 29040 8919
rect 29730 8916 29736 8968
rect 29788 8916 29794 8968
rect 30098 8916 30104 8968
rect 30156 8916 30162 8968
rect 30650 8916 30656 8968
rect 30708 8916 30714 8968
rect 30837 8959 30895 8965
rect 30837 8925 30849 8959
rect 30883 8925 30895 8959
rect 30837 8919 30895 8925
rect 28684 8860 29040 8888
rect 28684 8848 28690 8860
rect 29086 8848 29092 8900
rect 29144 8888 29150 8900
rect 29549 8891 29607 8897
rect 29549 8888 29561 8891
rect 29144 8860 29561 8888
rect 29144 8848 29150 8860
rect 29549 8857 29561 8860
rect 29595 8857 29607 8891
rect 29549 8851 29607 8857
rect 30374 8848 30380 8900
rect 30432 8848 30438 8900
rect 30852 8888 30880 8919
rect 31110 8916 31116 8968
rect 31168 8916 31174 8968
rect 31202 8916 31208 8968
rect 31260 8956 31266 8968
rect 31297 8959 31355 8965
rect 31297 8956 31309 8959
rect 31260 8928 31309 8956
rect 31260 8916 31266 8928
rect 31297 8925 31309 8928
rect 31343 8925 31355 8959
rect 32324 8956 32352 8996
rect 32398 8984 32404 9036
rect 32456 9024 32462 9036
rect 32953 9027 33011 9033
rect 32953 9024 32965 9027
rect 32456 8996 32965 9024
rect 32456 8984 32462 8996
rect 32953 8993 32965 8996
rect 32999 8993 33011 9027
rect 33410 9024 33416 9036
rect 32953 8987 33011 8993
rect 33244 8996 33416 9024
rect 32582 8956 32588 8968
rect 32324 8928 32588 8956
rect 31297 8919 31355 8925
rect 32582 8916 32588 8928
rect 32640 8916 32646 8968
rect 32769 8959 32827 8965
rect 32769 8925 32781 8959
rect 32815 8956 32827 8959
rect 32858 8956 32864 8968
rect 32815 8928 32864 8956
rect 32815 8925 32827 8928
rect 32769 8919 32827 8925
rect 32858 8916 32864 8928
rect 32916 8956 32922 8968
rect 33244 8956 33272 8996
rect 33410 8984 33416 8996
rect 33468 8984 33474 9036
rect 38289 9027 38347 9033
rect 38289 9024 38301 9027
rect 37292 8996 38301 9024
rect 35158 8956 35164 8968
rect 32916 8928 33272 8956
rect 33336 8928 35164 8956
rect 32916 8916 32922 8928
rect 33336 8900 33364 8928
rect 35158 8916 35164 8928
rect 35216 8916 35222 8968
rect 35434 8916 35440 8968
rect 35492 8956 35498 8968
rect 35713 8959 35771 8965
rect 35713 8956 35725 8959
rect 35492 8928 35725 8956
rect 35492 8916 35498 8928
rect 35713 8925 35725 8928
rect 35759 8925 35771 8959
rect 35713 8919 35771 8925
rect 36078 8916 36084 8968
rect 36136 8956 36142 8968
rect 37185 8959 37243 8965
rect 37185 8956 37197 8959
rect 36136 8928 37197 8956
rect 36136 8916 36142 8928
rect 37185 8925 37197 8928
rect 37231 8956 37243 8959
rect 37292 8956 37320 8996
rect 38289 8993 38301 8996
rect 38335 8993 38347 9027
rect 38289 8987 38347 8993
rect 37231 8928 37320 8956
rect 37369 8959 37427 8965
rect 37231 8925 37243 8928
rect 37185 8919 37243 8925
rect 37369 8925 37381 8959
rect 37415 8956 37427 8959
rect 37550 8956 37556 8968
rect 37415 8928 37556 8956
rect 37415 8925 37427 8928
rect 37369 8919 37427 8925
rect 37550 8916 37556 8928
rect 37608 8916 37614 8968
rect 37734 8956 37740 8968
rect 37676 8925 37740 8956
rect 31478 8888 31484 8900
rect 30852 8860 31484 8888
rect 31478 8848 31484 8860
rect 31536 8848 31542 8900
rect 33318 8848 33324 8900
rect 33376 8848 33382 8900
rect 33505 8891 33563 8897
rect 33505 8857 33517 8891
rect 33551 8888 33563 8891
rect 33594 8888 33600 8900
rect 33551 8860 33600 8888
rect 33551 8857 33563 8860
rect 33505 8851 33563 8857
rect 33594 8848 33600 8860
rect 33652 8888 33658 8900
rect 34422 8888 34428 8900
rect 33652 8860 34428 8888
rect 33652 8848 33658 8860
rect 34422 8848 34428 8860
rect 34480 8848 34486 8900
rect 36170 8848 36176 8900
rect 36228 8888 36234 8900
rect 37461 8891 37519 8897
rect 37676 8894 37703 8925
rect 37461 8888 37473 8891
rect 36228 8860 37473 8888
rect 36228 8848 36234 8860
rect 37461 8857 37473 8860
rect 37507 8857 37519 8891
rect 37691 8891 37703 8894
rect 37737 8916 37740 8925
rect 37792 8916 37798 8968
rect 37918 8916 37924 8968
rect 37976 8916 37982 8968
rect 37737 8891 37749 8916
rect 37691 8885 37749 8891
rect 38473 8891 38531 8897
rect 37461 8851 37519 8857
rect 38473 8857 38485 8891
rect 38519 8857 38531 8891
rect 38473 8851 38531 8857
rect 26326 8820 26332 8832
rect 26160 8792 26332 8820
rect 26326 8780 26332 8792
rect 26384 8780 26390 8832
rect 28534 8780 28540 8832
rect 28592 8820 28598 8832
rect 28902 8820 28908 8832
rect 28592 8792 28908 8820
rect 28592 8780 28598 8792
rect 28902 8780 28908 8792
rect 28960 8820 28966 8832
rect 30926 8820 30932 8832
rect 28960 8792 30932 8820
rect 28960 8780 28966 8792
rect 30926 8780 30932 8792
rect 30984 8780 30990 8832
rect 32674 8780 32680 8832
rect 32732 8820 32738 8832
rect 33413 8823 33471 8829
rect 33413 8820 33425 8823
rect 32732 8792 33425 8820
rect 32732 8780 32738 8792
rect 33413 8789 33425 8792
rect 33459 8820 33471 8823
rect 34514 8820 34520 8832
rect 33459 8792 34520 8820
rect 33459 8789 33471 8792
rect 33413 8783 33471 8789
rect 34514 8780 34520 8792
rect 34572 8820 34578 8832
rect 34974 8820 34980 8832
rect 34572 8792 34980 8820
rect 34572 8780 34578 8792
rect 34974 8780 34980 8792
rect 35032 8780 35038 8832
rect 35250 8780 35256 8832
rect 35308 8820 35314 8832
rect 38105 8823 38163 8829
rect 38105 8820 38117 8823
rect 35308 8792 38117 8820
rect 35308 8780 35314 8792
rect 38105 8789 38117 8792
rect 38151 8820 38163 8823
rect 38488 8820 38516 8851
rect 38151 8792 38516 8820
rect 38151 8789 38163 8792
rect 38105 8783 38163 8789
rect 1104 8730 40572 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 40572 8730
rect 1104 8656 40572 8678
rect 4249 8619 4307 8625
rect 4249 8585 4261 8619
rect 4295 8616 4307 8619
rect 5626 8616 5632 8628
rect 4295 8588 5632 8616
rect 4295 8585 4307 8588
rect 4249 8579 4307 8585
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 6914 8576 6920 8628
rect 6972 8616 6978 8628
rect 7193 8619 7251 8625
rect 7193 8616 7205 8619
rect 6972 8588 7205 8616
rect 6972 8576 6978 8588
rect 7193 8585 7205 8588
rect 7239 8585 7251 8619
rect 7193 8579 7251 8585
rect 7558 8576 7564 8628
rect 7616 8616 7622 8628
rect 8478 8616 8484 8628
rect 7616 8588 8484 8616
rect 7616 8576 7622 8588
rect 8478 8576 8484 8588
rect 8536 8616 8542 8628
rect 8536 8588 8800 8616
rect 8536 8576 8542 8588
rect 4706 8508 4712 8560
rect 4764 8508 4770 8560
rect 8294 8548 8300 8560
rect 6012 8520 8300 8548
rect 6012 8489 6040 8520
rect 8294 8508 8300 8520
rect 8352 8508 8358 8560
rect 5997 8483 6055 8489
rect 5997 8449 6009 8483
rect 6043 8449 6055 8483
rect 5997 8443 6055 8449
rect 6638 8440 6644 8492
rect 6696 8440 6702 8492
rect 6822 8440 6828 8492
rect 6880 8440 6886 8492
rect 6917 8483 6975 8489
rect 6917 8449 6929 8483
rect 6963 8480 6975 8483
rect 7098 8480 7104 8492
rect 6963 8452 7104 8480
rect 6963 8449 6975 8452
rect 6917 8443 6975 8449
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 7190 8440 7196 8492
rect 7248 8480 7254 8492
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 7248 8452 7389 8480
rect 7248 8440 7254 8452
rect 7377 8449 7389 8452
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 7466 8440 7472 8492
rect 7524 8440 7530 8492
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 5718 8372 5724 8424
rect 5776 8372 5782 8424
rect 6733 8415 6791 8421
rect 6733 8381 6745 8415
rect 6779 8412 6791 8415
rect 7006 8412 7012 8424
rect 6779 8384 7012 8412
rect 6779 8381 6791 8384
rect 6733 8375 6791 8381
rect 7006 8372 7012 8384
rect 7064 8372 7070 8424
rect 7282 8372 7288 8424
rect 7340 8412 7346 8424
rect 7576 8412 7604 8443
rect 7742 8440 7748 8492
rect 7800 8440 7806 8492
rect 7837 8483 7895 8489
rect 7837 8449 7849 8483
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 7340 8384 7604 8412
rect 7340 8372 7346 8384
rect 6454 8236 6460 8288
rect 6512 8236 6518 8288
rect 7852 8276 7880 8443
rect 8202 8440 8208 8492
rect 8260 8440 8266 8492
rect 8389 8483 8447 8489
rect 8389 8449 8401 8483
rect 8435 8480 8447 8483
rect 8478 8480 8484 8492
rect 8435 8452 8484 8480
rect 8435 8449 8447 8452
rect 8389 8443 8447 8449
rect 8478 8440 8484 8452
rect 8536 8440 8542 8492
rect 8772 8489 8800 8588
rect 8938 8576 8944 8628
rect 8996 8616 9002 8628
rect 11422 8616 11428 8628
rect 8996 8588 11428 8616
rect 8996 8576 9002 8588
rect 11422 8576 11428 8588
rect 11480 8576 11486 8628
rect 15562 8616 15568 8628
rect 13280 8588 15568 8616
rect 9858 8508 9864 8560
rect 9916 8548 9922 8560
rect 9916 8520 10548 8548
rect 9916 8508 9922 8520
rect 8757 8483 8815 8489
rect 8757 8449 8769 8483
rect 8803 8449 8815 8483
rect 8757 8443 8815 8449
rect 9030 8440 9036 8492
rect 9088 8440 9094 8492
rect 9122 8440 9128 8492
rect 9180 8480 9186 8492
rect 10321 8483 10379 8489
rect 10321 8480 10333 8483
rect 9180 8452 10333 8480
rect 9180 8440 9186 8452
rect 10321 8449 10333 8452
rect 10367 8480 10379 8483
rect 10410 8480 10416 8492
rect 10367 8452 10416 8480
rect 10367 8449 10379 8452
rect 10321 8443 10379 8449
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 10520 8489 10548 8520
rect 10505 8483 10563 8489
rect 10505 8449 10517 8483
rect 10551 8449 10563 8483
rect 10505 8443 10563 8449
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8449 10655 8483
rect 10597 8443 10655 8449
rect 7926 8372 7932 8424
rect 7984 8372 7990 8424
rect 8294 8421 8300 8424
rect 8113 8415 8171 8421
rect 8113 8381 8125 8415
rect 8159 8381 8171 8415
rect 8288 8412 8300 8421
rect 8255 8384 8300 8412
rect 8113 8375 8171 8381
rect 8288 8375 8300 8384
rect 8128 8344 8156 8375
rect 8294 8372 8300 8375
rect 8352 8372 8358 8424
rect 8662 8372 8668 8424
rect 8720 8412 8726 8424
rect 10612 8412 10640 8443
rect 10870 8440 10876 8492
rect 10928 8440 10934 8492
rect 11882 8440 11888 8492
rect 11940 8440 11946 8492
rect 12345 8483 12403 8489
rect 12345 8449 12357 8483
rect 12391 8480 12403 8483
rect 12526 8480 12532 8492
rect 12391 8452 12532 8480
rect 12391 8449 12403 8452
rect 12345 8443 12403 8449
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 8720 8384 10640 8412
rect 8720 8372 8726 8384
rect 10962 8372 10968 8424
rect 11020 8412 11026 8424
rect 11517 8415 11575 8421
rect 11517 8412 11529 8415
rect 11020 8384 11529 8412
rect 11020 8372 11026 8384
rect 11517 8381 11529 8384
rect 11563 8381 11575 8415
rect 13280 8412 13308 8588
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 15841 8619 15899 8625
rect 15841 8585 15853 8619
rect 15887 8585 15899 8619
rect 15841 8579 15899 8585
rect 14366 8508 14372 8560
rect 14424 8548 14430 8560
rect 14734 8548 14740 8560
rect 14424 8520 14740 8548
rect 14424 8508 14430 8520
rect 14734 8508 14740 8520
rect 14792 8508 14798 8560
rect 14829 8551 14887 8557
rect 14829 8517 14841 8551
rect 14875 8548 14887 8551
rect 15856 8548 15884 8579
rect 17862 8576 17868 8628
rect 17920 8616 17926 8628
rect 18782 8616 18788 8628
rect 17920 8588 18788 8616
rect 17920 8576 17926 8588
rect 18782 8576 18788 8588
rect 18840 8576 18846 8628
rect 20070 8576 20076 8628
rect 20128 8616 20134 8628
rect 20128 8588 20668 8616
rect 20128 8576 20134 8588
rect 19426 8548 19432 8560
rect 14875 8520 15884 8548
rect 18616 8520 19432 8548
rect 14875 8517 14887 8520
rect 14829 8511 14887 8517
rect 15194 8440 15200 8492
rect 15252 8440 15258 8492
rect 15286 8440 15292 8492
rect 15344 8440 15350 8492
rect 15473 8483 15531 8489
rect 15473 8449 15485 8483
rect 15519 8449 15531 8483
rect 15473 8443 15531 8449
rect 15565 8483 15623 8489
rect 15565 8449 15577 8483
rect 15611 8449 15623 8483
rect 15565 8443 15623 8449
rect 11517 8375 11575 8381
rect 12406 8384 13308 8412
rect 13357 8415 13415 8421
rect 8128 8316 8248 8344
rect 8110 8276 8116 8288
rect 7852 8248 8116 8276
rect 8110 8236 8116 8248
rect 8168 8236 8174 8288
rect 8220 8276 8248 8316
rect 8478 8304 8484 8356
rect 8536 8344 8542 8356
rect 8573 8347 8631 8353
rect 8573 8344 8585 8347
rect 8536 8316 8585 8344
rect 8536 8304 8542 8316
rect 8573 8313 8585 8316
rect 8619 8313 8631 8347
rect 8573 8307 8631 8313
rect 10413 8347 10471 8353
rect 10413 8313 10425 8347
rect 10459 8344 10471 8347
rect 10689 8347 10747 8353
rect 10689 8344 10701 8347
rect 10459 8316 10701 8344
rect 10459 8313 10471 8316
rect 10413 8307 10471 8313
rect 10689 8313 10701 8316
rect 10735 8313 10747 8347
rect 10689 8307 10747 8313
rect 11057 8347 11115 8353
rect 11057 8313 11069 8347
rect 11103 8344 11115 8347
rect 12406 8344 12434 8384
rect 13357 8381 13369 8415
rect 13403 8412 13415 8415
rect 14734 8412 14740 8424
rect 13403 8384 14740 8412
rect 13403 8381 13415 8384
rect 13357 8375 13415 8381
rect 14734 8372 14740 8384
rect 14792 8412 14798 8424
rect 15105 8415 15163 8421
rect 14792 8384 15056 8412
rect 14792 8372 14798 8384
rect 11103 8316 12434 8344
rect 15028 8344 15056 8384
rect 15105 8381 15117 8415
rect 15151 8412 15163 8415
rect 15378 8412 15384 8424
rect 15151 8384 15384 8412
rect 15151 8381 15163 8384
rect 15105 8375 15163 8381
rect 15378 8372 15384 8384
rect 15436 8372 15442 8424
rect 15488 8344 15516 8443
rect 15580 8412 15608 8443
rect 15654 8440 15660 8492
rect 15712 8440 15718 8492
rect 17586 8440 17592 8492
rect 17644 8440 17650 8492
rect 18616 8489 18644 8520
rect 19426 8508 19432 8520
rect 19484 8508 19490 8560
rect 20165 8551 20223 8557
rect 20165 8548 20177 8551
rect 19812 8520 20177 8548
rect 18601 8483 18659 8489
rect 18601 8449 18613 8483
rect 18647 8449 18659 8483
rect 18601 8443 18659 8449
rect 18690 8440 18696 8492
rect 18748 8440 18754 8492
rect 18782 8440 18788 8492
rect 18840 8480 18846 8492
rect 18877 8483 18935 8489
rect 18877 8480 18889 8483
rect 18840 8452 18889 8480
rect 18840 8440 18846 8452
rect 18877 8449 18889 8452
rect 18923 8449 18935 8483
rect 18877 8443 18935 8449
rect 19061 8483 19119 8489
rect 19061 8449 19073 8483
rect 19107 8480 19119 8483
rect 19150 8480 19156 8492
rect 19107 8452 19156 8480
rect 19107 8449 19119 8452
rect 19061 8443 19119 8449
rect 19150 8440 19156 8452
rect 19208 8440 19214 8492
rect 19610 8440 19616 8492
rect 19668 8440 19674 8492
rect 17310 8412 17316 8424
rect 15580 8384 17316 8412
rect 17310 8372 17316 8384
rect 17368 8372 17374 8424
rect 17678 8372 17684 8424
rect 17736 8372 17742 8424
rect 17865 8415 17923 8421
rect 17865 8381 17877 8415
rect 17911 8412 17923 8415
rect 17954 8412 17960 8424
rect 17911 8384 17960 8412
rect 17911 8381 17923 8384
rect 17865 8375 17923 8381
rect 17954 8372 17960 8384
rect 18012 8372 18018 8424
rect 19242 8372 19248 8424
rect 19300 8412 19306 8424
rect 19812 8421 19840 8520
rect 20165 8517 20177 8520
rect 20211 8517 20223 8551
rect 20165 8511 20223 8517
rect 20254 8508 20260 8560
rect 20312 8548 20318 8560
rect 20312 8520 20576 8548
rect 20312 8508 20318 8520
rect 19889 8483 19947 8489
rect 19889 8449 19901 8483
rect 19935 8480 19947 8483
rect 19978 8480 19984 8492
rect 19935 8452 19984 8480
rect 19935 8449 19947 8452
rect 19889 8443 19947 8449
rect 19978 8440 19984 8452
rect 20036 8440 20042 8492
rect 20070 8440 20076 8492
rect 20128 8440 20134 8492
rect 20548 8489 20576 8520
rect 20640 8492 20668 8588
rect 20990 8576 20996 8628
rect 21048 8616 21054 8628
rect 21048 8588 23060 8616
rect 21048 8576 21054 8588
rect 20714 8508 20720 8560
rect 20772 8548 20778 8560
rect 21821 8551 21879 8557
rect 21821 8548 21833 8551
rect 20772 8520 21833 8548
rect 20772 8508 20778 8520
rect 21821 8517 21833 8520
rect 21867 8548 21879 8551
rect 22031 8551 22089 8557
rect 21867 8520 21956 8548
rect 21867 8517 21879 8520
rect 21821 8511 21879 8517
rect 20441 8483 20499 8489
rect 20441 8449 20453 8483
rect 20487 8449 20499 8483
rect 20441 8443 20499 8449
rect 20533 8483 20591 8489
rect 20533 8449 20545 8483
rect 20579 8449 20591 8483
rect 20533 8443 20591 8449
rect 19797 8415 19855 8421
rect 19797 8412 19809 8415
rect 19300 8384 19809 8412
rect 19300 8372 19306 8384
rect 19797 8381 19809 8384
rect 19843 8381 19855 8415
rect 20456 8412 20484 8443
rect 20622 8440 20628 8492
rect 20680 8440 20686 8492
rect 20806 8440 20812 8492
rect 20864 8440 20870 8492
rect 21174 8440 21180 8492
rect 21232 8480 21238 8492
rect 21361 8483 21419 8489
rect 21361 8480 21373 8483
rect 21232 8452 21373 8480
rect 21232 8440 21238 8452
rect 21361 8449 21373 8452
rect 21407 8449 21419 8483
rect 21928 8480 21956 8520
rect 22031 8517 22043 8551
rect 22077 8548 22089 8551
rect 22278 8548 22284 8560
rect 22077 8520 22284 8548
rect 22077 8517 22089 8520
rect 22031 8511 22089 8517
rect 22278 8508 22284 8520
rect 22336 8508 22342 8560
rect 22738 8480 22744 8492
rect 21928 8452 22744 8480
rect 21361 8443 21419 8449
rect 22738 8440 22744 8452
rect 22796 8440 22802 8492
rect 21726 8412 21732 8424
rect 20456 8384 21732 8412
rect 19797 8375 19855 8381
rect 21726 8372 21732 8384
rect 21784 8412 21790 8424
rect 22646 8412 22652 8424
rect 21784 8384 22652 8412
rect 21784 8372 21790 8384
rect 22646 8372 22652 8384
rect 22704 8372 22710 8424
rect 23032 8412 23060 8588
rect 23106 8576 23112 8628
rect 23164 8576 23170 8628
rect 23290 8576 23296 8628
rect 23348 8616 23354 8628
rect 23385 8619 23443 8625
rect 23385 8616 23397 8619
rect 23348 8588 23397 8616
rect 23348 8576 23354 8588
rect 23385 8585 23397 8588
rect 23431 8585 23443 8619
rect 23842 8616 23848 8628
rect 23385 8579 23443 8585
rect 23492 8588 23848 8616
rect 23293 8483 23351 8489
rect 23293 8449 23305 8483
rect 23339 8480 23351 8483
rect 23492 8480 23520 8588
rect 23842 8576 23848 8588
rect 23900 8576 23906 8628
rect 24946 8616 24952 8628
rect 24780 8588 24952 8616
rect 23553 8551 23611 8557
rect 23553 8517 23565 8551
rect 23599 8548 23611 8551
rect 23599 8517 23612 8548
rect 23553 8511 23612 8517
rect 23339 8452 23520 8480
rect 23339 8449 23351 8452
rect 23293 8443 23351 8449
rect 23584 8412 23612 8511
rect 23750 8508 23756 8560
rect 23808 8508 23814 8560
rect 24118 8508 24124 8560
rect 24176 8508 24182 8560
rect 24210 8508 24216 8560
rect 24268 8508 24274 8560
rect 24780 8557 24808 8588
rect 24946 8576 24952 8588
rect 25004 8576 25010 8628
rect 27062 8576 27068 8628
rect 27120 8576 27126 8628
rect 28169 8619 28227 8625
rect 28169 8616 28181 8619
rect 27172 8588 28181 8616
rect 24765 8551 24823 8557
rect 24765 8517 24777 8551
rect 24811 8517 24823 8551
rect 24765 8511 24823 8517
rect 26142 8508 26148 8560
rect 26200 8548 26206 8560
rect 27172 8548 27200 8588
rect 28169 8585 28181 8588
rect 28215 8616 28227 8619
rect 28215 8588 28580 8616
rect 28215 8585 28227 8588
rect 28169 8579 28227 8585
rect 26200 8520 27200 8548
rect 26200 8508 26206 8520
rect 27430 8508 27436 8560
rect 27488 8548 27494 8560
rect 27488 8520 27660 8548
rect 27488 8508 27494 8520
rect 24026 8440 24032 8492
rect 24084 8440 24090 8492
rect 24397 8483 24455 8489
rect 24397 8449 24409 8483
rect 24443 8480 24455 8483
rect 24578 8480 24584 8492
rect 24443 8452 24584 8480
rect 24443 8449 24455 8452
rect 24397 8443 24455 8449
rect 24412 8412 24440 8443
rect 24578 8440 24584 8452
rect 24636 8440 24642 8492
rect 24857 8483 24915 8489
rect 24857 8449 24869 8483
rect 24903 8449 24915 8483
rect 24857 8443 24915 8449
rect 23032 8384 24440 8412
rect 24762 8372 24768 8424
rect 24820 8412 24826 8424
rect 24872 8412 24900 8443
rect 25222 8440 25228 8492
rect 25280 8440 25286 8492
rect 25682 8440 25688 8492
rect 25740 8440 25746 8492
rect 25774 8440 25780 8492
rect 25832 8480 25838 8492
rect 25961 8483 26019 8489
rect 25961 8480 25973 8483
rect 25832 8452 25973 8480
rect 25832 8440 25838 8452
rect 25961 8449 25973 8452
rect 26007 8449 26019 8483
rect 25961 8443 26019 8449
rect 26694 8440 26700 8492
rect 26752 8440 26758 8492
rect 27249 8483 27307 8489
rect 27249 8449 27261 8483
rect 27295 8480 27307 8483
rect 27522 8480 27528 8492
rect 27295 8452 27528 8480
rect 27295 8449 27307 8452
rect 27249 8443 27307 8449
rect 27522 8440 27528 8452
rect 27580 8440 27586 8492
rect 27632 8489 27660 8520
rect 27706 8508 27712 8560
rect 27764 8548 27770 8560
rect 28552 8548 28580 8588
rect 28626 8576 28632 8628
rect 28684 8576 28690 8628
rect 28718 8576 28724 8628
rect 28776 8576 28782 8628
rect 28810 8576 28816 8628
rect 28868 8616 28874 8628
rect 31202 8616 31208 8628
rect 28868 8588 31208 8616
rect 28868 8576 28874 8588
rect 31202 8576 31208 8588
rect 31260 8576 31266 8628
rect 33778 8576 33784 8628
rect 33836 8576 33842 8628
rect 33962 8576 33968 8628
rect 34020 8616 34026 8628
rect 34020 8588 34192 8616
rect 34020 8576 34026 8588
rect 28994 8548 29000 8560
rect 27764 8520 28396 8548
rect 28552 8520 29000 8548
rect 27764 8508 27770 8520
rect 28368 8489 28396 8520
rect 28994 8508 29000 8520
rect 29052 8548 29058 8560
rect 29052 8520 29224 8548
rect 29052 8508 29058 8520
rect 27617 8483 27675 8489
rect 27617 8449 27629 8483
rect 27663 8480 27675 8483
rect 27893 8483 27951 8489
rect 27893 8480 27905 8483
rect 27663 8452 27905 8480
rect 27663 8449 27675 8452
rect 27617 8443 27675 8449
rect 27893 8449 27905 8452
rect 27939 8449 27951 8483
rect 27893 8443 27951 8449
rect 28261 8483 28319 8489
rect 28261 8449 28273 8483
rect 28307 8449 28319 8483
rect 28261 8443 28319 8449
rect 28353 8483 28411 8489
rect 28353 8449 28365 8483
rect 28399 8449 28411 8483
rect 28353 8443 28411 8449
rect 24820 8384 24900 8412
rect 24820 8372 24826 8384
rect 27062 8372 27068 8424
rect 27120 8412 27126 8424
rect 27338 8412 27344 8424
rect 27120 8384 27344 8412
rect 27120 8372 27126 8384
rect 27338 8372 27344 8384
rect 27396 8412 27402 8424
rect 27709 8415 27767 8421
rect 27709 8412 27721 8415
rect 27396 8384 27721 8412
rect 27396 8372 27402 8384
rect 27709 8381 27721 8384
rect 27755 8412 27767 8415
rect 28276 8412 28304 8443
rect 28902 8440 28908 8492
rect 28960 8440 28966 8492
rect 29086 8440 29092 8492
rect 29144 8440 29150 8492
rect 29196 8489 29224 8520
rect 29822 8508 29828 8560
rect 29880 8548 29886 8560
rect 34054 8548 34060 8560
rect 29880 8520 34060 8548
rect 29880 8508 29886 8520
rect 29181 8483 29239 8489
rect 29181 8449 29193 8483
rect 29227 8449 29239 8483
rect 29181 8443 29239 8449
rect 29641 8483 29699 8489
rect 29641 8449 29653 8483
rect 29687 8449 29699 8483
rect 29641 8443 29699 8449
rect 29104 8412 29132 8440
rect 27755 8384 29132 8412
rect 29656 8412 29684 8443
rect 29730 8440 29736 8492
rect 29788 8440 29794 8492
rect 29840 8452 30604 8480
rect 29840 8412 29868 8452
rect 29656 8384 29868 8412
rect 27755 8381 27767 8384
rect 27709 8375 27767 8381
rect 30006 8372 30012 8424
rect 30064 8372 30070 8424
rect 30576 8412 30604 8452
rect 30650 8440 30656 8492
rect 30708 8440 30714 8492
rect 31570 8440 31576 8492
rect 31628 8480 31634 8492
rect 31754 8480 31760 8492
rect 31628 8452 31760 8480
rect 31628 8440 31634 8452
rect 31754 8440 31760 8452
rect 31812 8440 31818 8492
rect 32324 8489 32352 8520
rect 34054 8508 34060 8520
rect 34112 8508 34118 8560
rect 34164 8548 34192 8588
rect 34238 8576 34244 8628
rect 34296 8576 34302 8628
rect 34514 8576 34520 8628
rect 34572 8576 34578 8628
rect 36078 8576 36084 8628
rect 36136 8576 36142 8628
rect 36170 8576 36176 8628
rect 36228 8576 36234 8628
rect 37734 8576 37740 8628
rect 37792 8616 37798 8628
rect 37921 8619 37979 8625
rect 37921 8616 37933 8619
rect 37792 8588 37933 8616
rect 37792 8576 37798 8588
rect 37921 8585 37933 8588
rect 37967 8585 37979 8619
rect 37921 8579 37979 8585
rect 38562 8576 38568 8628
rect 38620 8576 38626 8628
rect 34609 8551 34667 8557
rect 34609 8548 34621 8551
rect 34164 8520 34621 8548
rect 34609 8517 34621 8520
rect 34655 8548 34667 8551
rect 35434 8548 35440 8560
rect 34655 8520 35440 8548
rect 34655 8517 34667 8520
rect 34609 8511 34667 8517
rect 35434 8508 35440 8520
rect 35492 8548 35498 8560
rect 36633 8551 36691 8557
rect 36633 8548 36645 8551
rect 35492 8520 36645 8548
rect 35492 8508 35498 8520
rect 36633 8517 36645 8520
rect 36679 8548 36691 8551
rect 37458 8548 37464 8560
rect 36679 8520 37464 8548
rect 36679 8517 36691 8520
rect 36633 8511 36691 8517
rect 37458 8508 37464 8520
rect 37516 8508 37522 8560
rect 38580 8548 38608 8576
rect 38749 8551 38807 8557
rect 38749 8548 38761 8551
rect 38580 8520 38761 8548
rect 38749 8517 38761 8520
rect 38795 8517 38807 8551
rect 38749 8511 38807 8517
rect 39022 8508 39028 8560
rect 39080 8548 39086 8560
rect 39080 8520 39238 8548
rect 39080 8508 39086 8520
rect 32309 8483 32367 8489
rect 32309 8449 32321 8483
rect 32355 8449 32367 8483
rect 32309 8443 32367 8449
rect 32582 8440 32588 8492
rect 32640 8480 32646 8492
rect 33962 8480 33968 8492
rect 32640 8452 33968 8480
rect 32640 8440 32646 8452
rect 33962 8440 33968 8452
rect 34020 8440 34026 8492
rect 35897 8483 35955 8489
rect 34440 8480 34560 8483
rect 35897 8480 35909 8483
rect 34164 8455 35909 8480
rect 34164 8452 34468 8455
rect 34532 8452 35909 8455
rect 30742 8412 30748 8424
rect 30576 8384 30748 8412
rect 30742 8372 30748 8384
rect 30800 8372 30806 8424
rect 30926 8372 30932 8424
rect 30984 8412 30990 8424
rect 33042 8412 33048 8424
rect 30984 8384 33048 8412
rect 30984 8372 30990 8384
rect 33042 8372 33048 8384
rect 33100 8372 33106 8424
rect 33321 8415 33379 8421
rect 33321 8381 33333 8415
rect 33367 8412 33379 8415
rect 33870 8412 33876 8424
rect 33367 8384 33876 8412
rect 33367 8381 33379 8384
rect 33321 8375 33379 8381
rect 33870 8372 33876 8384
rect 33928 8372 33934 8424
rect 34164 8412 34192 8452
rect 35897 8449 35909 8452
rect 35943 8480 35955 8483
rect 36538 8480 36544 8492
rect 35943 8452 36544 8480
rect 35943 8449 35955 8452
rect 35897 8443 35955 8449
rect 36538 8440 36544 8452
rect 36596 8440 36602 8492
rect 37734 8440 37740 8492
rect 37792 8440 37798 8492
rect 33980 8384 34192 8412
rect 34400 8415 34458 8421
rect 17696 8344 17724 8372
rect 15028 8316 15516 8344
rect 15764 8316 17724 8344
rect 11103 8313 11115 8316
rect 11057 8307 11115 8313
rect 8386 8276 8392 8288
rect 8220 8248 8392 8276
rect 8386 8236 8392 8248
rect 8444 8276 8450 8288
rect 9122 8276 9128 8288
rect 8444 8248 9128 8276
rect 8444 8236 8450 8248
rect 9122 8236 9128 8248
rect 9180 8236 9186 8288
rect 15102 8236 15108 8288
rect 15160 8276 15166 8288
rect 15764 8276 15792 8316
rect 18322 8304 18328 8356
rect 18380 8344 18386 8356
rect 18785 8347 18843 8353
rect 18785 8344 18797 8347
rect 18380 8316 18797 8344
rect 18380 8304 18386 8316
rect 18785 8313 18797 8316
rect 18831 8313 18843 8347
rect 18785 8307 18843 8313
rect 18874 8304 18880 8356
rect 18932 8344 18938 8356
rect 19337 8347 19395 8353
rect 19337 8344 19349 8347
rect 18932 8316 19349 8344
rect 18932 8304 18938 8316
rect 19337 8313 19349 8316
rect 19383 8313 19395 8347
rect 19337 8307 19395 8313
rect 22186 8304 22192 8356
rect 22244 8304 22250 8356
rect 23934 8304 23940 8356
rect 23992 8344 23998 8356
rect 28258 8344 28264 8356
rect 23992 8316 28264 8344
rect 23992 8304 23998 8316
rect 28258 8304 28264 8316
rect 28316 8304 28322 8356
rect 28442 8304 28448 8356
rect 28500 8344 28506 8356
rect 28500 8316 28764 8344
rect 28500 8304 28506 8316
rect 15160 8248 15792 8276
rect 15160 8236 15166 8248
rect 15838 8236 15844 8288
rect 15896 8276 15902 8288
rect 17221 8279 17279 8285
rect 17221 8276 17233 8279
rect 15896 8248 17233 8276
rect 15896 8236 15902 8248
rect 17221 8245 17233 8248
rect 17267 8245 17279 8279
rect 17221 8239 17279 8245
rect 18414 8236 18420 8288
rect 18472 8236 18478 8288
rect 19705 8279 19763 8285
rect 19705 8245 19717 8279
rect 19751 8276 19763 8279
rect 20438 8276 20444 8288
rect 19751 8248 20444 8276
rect 19751 8245 19763 8248
rect 19705 8239 19763 8245
rect 20438 8236 20444 8248
rect 20496 8236 20502 8288
rect 20898 8236 20904 8288
rect 20956 8276 20962 8288
rect 21269 8279 21327 8285
rect 21269 8276 21281 8279
rect 20956 8248 21281 8276
rect 20956 8236 20962 8248
rect 21269 8245 21281 8248
rect 21315 8276 21327 8279
rect 21634 8276 21640 8288
rect 21315 8248 21640 8276
rect 21315 8245 21327 8248
rect 21269 8239 21327 8245
rect 21634 8236 21640 8248
rect 21692 8236 21698 8288
rect 21818 8236 21824 8288
rect 21876 8276 21882 8288
rect 22005 8279 22063 8285
rect 22005 8276 22017 8279
rect 21876 8248 22017 8276
rect 21876 8236 21882 8248
rect 22005 8245 22017 8248
rect 22051 8245 22063 8279
rect 22005 8239 22063 8245
rect 23474 8236 23480 8288
rect 23532 8276 23538 8288
rect 23569 8279 23627 8285
rect 23569 8276 23581 8279
rect 23532 8248 23581 8276
rect 23532 8236 23538 8248
rect 23569 8245 23581 8248
rect 23615 8245 23627 8279
rect 23569 8239 23627 8245
rect 23842 8236 23848 8288
rect 23900 8236 23906 8288
rect 26418 8236 26424 8288
rect 26476 8276 26482 8288
rect 26970 8276 26976 8288
rect 26476 8248 26976 8276
rect 26476 8236 26482 8248
rect 26970 8236 26976 8248
rect 27028 8236 27034 8288
rect 27249 8279 27307 8285
rect 27249 8245 27261 8279
rect 27295 8276 27307 8279
rect 27798 8276 27804 8288
rect 27295 8248 27804 8276
rect 27295 8245 27307 8248
rect 27249 8239 27307 8245
rect 27798 8236 27804 8248
rect 27856 8236 27862 8288
rect 27985 8279 28043 8285
rect 27985 8245 27997 8279
rect 28031 8276 28043 8279
rect 28626 8276 28632 8288
rect 28031 8248 28632 8276
rect 28031 8245 28043 8248
rect 27985 8239 28043 8245
rect 28626 8236 28632 8248
rect 28684 8236 28690 8288
rect 28736 8276 28764 8316
rect 28994 8304 29000 8356
rect 29052 8304 29058 8356
rect 29089 8347 29147 8353
rect 29089 8313 29101 8347
rect 29135 8344 29147 8347
rect 29135 8316 33640 8344
rect 29135 8313 29147 8316
rect 29089 8307 29147 8313
rect 29457 8279 29515 8285
rect 29457 8276 29469 8279
rect 28736 8248 29469 8276
rect 29457 8245 29469 8248
rect 29503 8276 29515 8279
rect 29822 8276 29828 8288
rect 29503 8248 29828 8276
rect 29503 8245 29515 8248
rect 29457 8239 29515 8245
rect 29822 8236 29828 8248
rect 29880 8236 29886 8288
rect 30190 8236 30196 8288
rect 30248 8276 30254 8288
rect 30374 8276 30380 8288
rect 30248 8248 30380 8276
rect 30248 8236 30254 8248
rect 30374 8236 30380 8248
rect 30432 8236 30438 8288
rect 31018 8236 31024 8288
rect 31076 8276 31082 8288
rect 32125 8279 32183 8285
rect 32125 8276 32137 8279
rect 31076 8248 32137 8276
rect 31076 8236 31082 8248
rect 32125 8245 32137 8248
rect 32171 8245 32183 8279
rect 32125 8239 32183 8245
rect 32306 8236 32312 8288
rect 32364 8276 32370 8288
rect 32401 8279 32459 8285
rect 32401 8276 32413 8279
rect 32364 8248 32413 8276
rect 32364 8236 32370 8248
rect 32401 8245 32413 8248
rect 32447 8245 32459 8279
rect 33612 8276 33640 8316
rect 33686 8304 33692 8356
rect 33744 8304 33750 8356
rect 33980 8344 34008 8384
rect 34400 8381 34412 8415
rect 34446 8381 34458 8415
rect 34400 8375 34458 8381
rect 33888 8316 34008 8344
rect 34415 8344 34443 8375
rect 34514 8372 34520 8424
rect 34572 8412 34578 8424
rect 34885 8415 34943 8421
rect 34885 8412 34897 8415
rect 34572 8384 34897 8412
rect 34572 8372 34578 8384
rect 34885 8381 34897 8384
rect 34931 8381 34943 8415
rect 34885 8375 34943 8381
rect 34698 8344 34704 8356
rect 34415 8316 34704 8344
rect 33888 8276 33916 8316
rect 34698 8304 34704 8316
rect 34756 8304 34762 8356
rect 34900 8344 34928 8375
rect 34974 8372 34980 8424
rect 35032 8412 35038 8424
rect 35032 8384 36676 8412
rect 35032 8372 35038 8384
rect 36170 8344 36176 8356
rect 34900 8316 36176 8344
rect 36170 8304 36176 8316
rect 36228 8304 36234 8356
rect 36648 8353 36676 8384
rect 38470 8372 38476 8424
rect 38528 8372 38534 8424
rect 40221 8415 40279 8421
rect 40221 8412 40233 8415
rect 38580 8384 40233 8412
rect 36633 8347 36691 8353
rect 36633 8313 36645 8347
rect 36679 8344 36691 8347
rect 37550 8344 37556 8356
rect 36679 8316 37556 8344
rect 36679 8313 36691 8316
rect 36633 8307 36691 8313
rect 37550 8304 37556 8316
rect 37608 8304 37614 8356
rect 33612 8248 33916 8276
rect 32401 8239 32459 8245
rect 35158 8236 35164 8288
rect 35216 8276 35222 8288
rect 37826 8276 37832 8288
rect 35216 8248 37832 8276
rect 35216 8236 35222 8248
rect 37826 8236 37832 8248
rect 37884 8276 37890 8288
rect 38580 8276 38608 8384
rect 40221 8381 40233 8384
rect 40267 8381 40279 8415
rect 40221 8375 40279 8381
rect 37884 8248 38608 8276
rect 37884 8236 37890 8248
rect 1104 8186 40572 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 40572 8186
rect 1104 8112 40572 8134
rect 5169 8075 5227 8081
rect 5169 8041 5181 8075
rect 5215 8072 5227 8075
rect 5718 8072 5724 8084
rect 5215 8044 5724 8072
rect 5215 8041 5227 8044
rect 5169 8035 5227 8041
rect 5718 8032 5724 8044
rect 5776 8032 5782 8084
rect 6730 8032 6736 8084
rect 6788 8072 6794 8084
rect 7926 8072 7932 8084
rect 6788 8044 7932 8072
rect 6788 8032 6794 8044
rect 7926 8032 7932 8044
rect 7984 8032 7990 8084
rect 8202 8032 8208 8084
rect 8260 8072 8266 8084
rect 11241 8075 11299 8081
rect 8260 8044 9812 8072
rect 8260 8032 8266 8044
rect 7101 8007 7159 8013
rect 7101 7973 7113 8007
rect 7147 8004 7159 8007
rect 7190 8004 7196 8016
rect 7147 7976 7196 8004
rect 7147 7973 7159 7976
rect 7101 7967 7159 7973
rect 7190 7964 7196 7976
rect 7248 7964 7254 8016
rect 7837 8007 7895 8013
rect 7837 7973 7849 8007
rect 7883 8004 7895 8007
rect 8021 8007 8079 8013
rect 8021 8004 8033 8007
rect 7883 7976 8033 8004
rect 7883 7973 7895 7976
rect 7837 7967 7895 7973
rect 8021 7973 8033 7976
rect 8067 7973 8079 8007
rect 9030 8004 9036 8016
rect 8021 7967 8079 7973
rect 8128 7976 9036 8004
rect 5626 7896 5632 7948
rect 5684 7896 5690 7948
rect 5813 7939 5871 7945
rect 5813 7905 5825 7939
rect 5859 7936 5871 7939
rect 6546 7936 6552 7948
rect 5859 7908 6552 7936
rect 5859 7905 5871 7908
rect 5813 7899 5871 7905
rect 6546 7896 6552 7908
rect 6604 7896 6610 7948
rect 6825 7939 6883 7945
rect 6825 7905 6837 7939
rect 6871 7936 6883 7939
rect 7377 7939 7435 7945
rect 7377 7936 7389 7939
rect 6871 7908 7389 7936
rect 6871 7905 6883 7908
rect 6825 7899 6883 7905
rect 7377 7905 7389 7908
rect 7423 7905 7435 7939
rect 7852 7936 7880 7967
rect 7377 7899 7435 7905
rect 7484 7908 7880 7936
rect 5537 7871 5595 7877
rect 5537 7837 5549 7871
rect 5583 7868 5595 7871
rect 6454 7868 6460 7880
rect 5583 7840 6460 7868
rect 5583 7837 5595 7840
rect 5537 7831 5595 7837
rect 6454 7828 6460 7840
rect 6512 7828 6518 7880
rect 6730 7828 6736 7880
rect 6788 7828 6794 7880
rect 7484 7877 7512 7908
rect 7926 7896 7932 7948
rect 7984 7896 7990 7948
rect 7285 7871 7343 7877
rect 7285 7837 7297 7871
rect 7331 7837 7343 7871
rect 7285 7831 7343 7837
rect 7469 7871 7527 7877
rect 7469 7837 7481 7871
rect 7515 7837 7527 7871
rect 7469 7831 7527 7837
rect 7300 7732 7328 7831
rect 7558 7828 7564 7880
rect 7616 7828 7622 7880
rect 7834 7828 7840 7880
rect 7892 7828 7898 7880
rect 7745 7803 7803 7809
rect 7745 7769 7757 7803
rect 7791 7800 7803 7803
rect 8128 7800 8156 7976
rect 9030 7964 9036 7976
rect 9088 7964 9094 8016
rect 9784 8004 9812 8044
rect 11241 8041 11253 8075
rect 11287 8072 11299 8075
rect 11882 8072 11888 8084
rect 11287 8044 11888 8072
rect 11287 8041 11299 8044
rect 11241 8035 11299 8041
rect 11882 8032 11888 8044
rect 11940 8032 11946 8084
rect 11974 8032 11980 8084
rect 12032 8072 12038 8084
rect 12710 8072 12716 8084
rect 12032 8044 12716 8072
rect 12032 8032 12038 8044
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 14553 8075 14611 8081
rect 14553 8041 14565 8075
rect 14599 8072 14611 8075
rect 15194 8072 15200 8084
rect 14599 8044 15200 8072
rect 14599 8041 14611 8044
rect 14553 8035 14611 8041
rect 15194 8032 15200 8044
rect 15252 8032 15258 8084
rect 15286 8032 15292 8084
rect 15344 8032 15350 8084
rect 16666 8072 16672 8084
rect 15672 8044 16672 8072
rect 10962 8004 10968 8016
rect 9784 7976 10968 8004
rect 8205 7939 8263 7945
rect 8205 7905 8217 7939
rect 8251 7936 8263 7939
rect 8294 7936 8300 7948
rect 8251 7908 8300 7936
rect 8251 7905 8263 7908
rect 8205 7899 8263 7905
rect 7791 7772 8156 7800
rect 7791 7769 7803 7772
rect 7745 7763 7803 7769
rect 8220 7732 8248 7899
rect 8294 7896 8300 7908
rect 8352 7896 8358 7948
rect 8386 7896 8392 7948
rect 8444 7896 8450 7948
rect 9784 7945 9812 7976
rect 10962 7964 10968 7976
rect 11020 7964 11026 8016
rect 11149 8007 11207 8013
rect 11149 7973 11161 8007
rect 11195 8004 11207 8007
rect 11422 8004 11428 8016
rect 11195 7976 11428 8004
rect 11195 7973 11207 7976
rect 11149 7967 11207 7973
rect 11422 7964 11428 7976
rect 11480 7964 11486 8016
rect 15102 7964 15108 8016
rect 15160 7964 15166 8016
rect 15562 7964 15568 8016
rect 15620 7964 15626 8016
rect 9769 7939 9827 7945
rect 9769 7905 9781 7939
rect 9815 7905 9827 7939
rect 9769 7899 9827 7905
rect 8481 7871 8539 7877
rect 8481 7837 8493 7871
rect 8527 7868 8539 7871
rect 9677 7871 9735 7877
rect 9677 7868 9689 7871
rect 8527 7840 9689 7868
rect 8527 7837 8539 7840
rect 8481 7831 8539 7837
rect 9677 7837 9689 7840
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 8297 7803 8355 7809
rect 8297 7769 8309 7803
rect 8343 7800 8355 7803
rect 9784 7800 9812 7899
rect 9858 7896 9864 7948
rect 9916 7896 9922 7948
rect 9953 7939 10011 7945
rect 9953 7905 9965 7939
rect 9999 7936 10011 7939
rect 10318 7936 10324 7948
rect 9999 7908 10324 7936
rect 9999 7905 10011 7908
rect 9953 7899 10011 7905
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 10686 7896 10692 7948
rect 10744 7936 10750 7948
rect 10781 7939 10839 7945
rect 10781 7936 10793 7939
rect 10744 7908 10793 7936
rect 10744 7896 10750 7908
rect 10781 7905 10793 7908
rect 10827 7905 10839 7939
rect 10781 7899 10839 7905
rect 13909 7871 13967 7877
rect 13909 7837 13921 7871
rect 13955 7868 13967 7871
rect 13998 7868 14004 7880
rect 13955 7840 14004 7868
rect 13955 7837 13967 7840
rect 13909 7831 13967 7837
rect 13998 7828 14004 7840
rect 14056 7828 14062 7880
rect 14090 7828 14096 7880
rect 14148 7828 14154 7880
rect 14369 7871 14427 7877
rect 14369 7837 14381 7871
rect 14415 7837 14427 7871
rect 14369 7831 14427 7837
rect 14553 7871 14611 7877
rect 14553 7837 14565 7871
rect 14599 7868 14611 7871
rect 14734 7868 14740 7880
rect 14599 7840 14740 7868
rect 14599 7837 14611 7840
rect 14553 7831 14611 7837
rect 8343 7772 9812 7800
rect 8343 7769 8355 7772
rect 8297 7763 8355 7769
rect 11606 7760 11612 7812
rect 11664 7800 11670 7812
rect 11790 7800 11796 7812
rect 11664 7772 11796 7800
rect 11664 7760 11670 7772
rect 11790 7760 11796 7772
rect 11848 7800 11854 7812
rect 14384 7800 14412 7831
rect 14734 7828 14740 7840
rect 14792 7828 14798 7880
rect 14829 7871 14887 7877
rect 14829 7837 14841 7871
rect 14875 7868 14887 7871
rect 15286 7868 15292 7880
rect 14875 7840 15292 7868
rect 14875 7837 14887 7840
rect 14829 7831 14887 7837
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 15580 7877 15608 7964
rect 15672 7877 15700 8044
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 17310 8032 17316 8084
rect 17368 8072 17374 8084
rect 18782 8072 18788 8084
rect 17368 8044 18788 8072
rect 17368 8032 17374 8044
rect 18782 8032 18788 8044
rect 18840 8032 18846 8084
rect 19426 8032 19432 8084
rect 19484 8032 19490 8084
rect 19536 8044 23336 8072
rect 19536 8004 19564 8044
rect 17420 7976 19564 8004
rect 20257 8007 20315 8013
rect 15746 7896 15752 7948
rect 15804 7936 15810 7948
rect 16025 7939 16083 7945
rect 16025 7936 16037 7939
rect 15804 7908 16037 7936
rect 15804 7896 15810 7908
rect 16025 7905 16037 7908
rect 16071 7905 16083 7939
rect 16025 7899 16083 7905
rect 16298 7896 16304 7948
rect 16356 7936 16362 7948
rect 17420 7936 17448 7976
rect 20257 7973 20269 8007
rect 20303 8004 20315 8007
rect 20346 8004 20352 8016
rect 20303 7976 20352 8004
rect 20303 7973 20315 7976
rect 20257 7967 20315 7973
rect 20346 7964 20352 7976
rect 20404 7964 20410 8016
rect 20622 7964 20628 8016
rect 20680 8004 20686 8016
rect 22370 8004 22376 8016
rect 20680 7976 22376 8004
rect 20680 7964 20686 7976
rect 22370 7964 22376 7976
rect 22428 7964 22434 8016
rect 22830 7964 22836 8016
rect 22888 8004 22894 8016
rect 22888 7976 23244 8004
rect 22888 7964 22894 7976
rect 19334 7936 19340 7948
rect 16356 7908 17448 7936
rect 18708 7908 19340 7936
rect 16356 7896 16362 7908
rect 15565 7871 15623 7877
rect 15565 7837 15577 7871
rect 15611 7837 15623 7871
rect 15565 7831 15623 7837
rect 15657 7871 15715 7877
rect 15657 7837 15669 7871
rect 15703 7837 15715 7871
rect 15657 7831 15715 7837
rect 15838 7828 15844 7880
rect 15896 7828 15902 7880
rect 15930 7828 15936 7880
rect 15988 7828 15994 7880
rect 18138 7828 18144 7880
rect 18196 7868 18202 7880
rect 18708 7877 18736 7908
rect 19334 7896 19340 7908
rect 19392 7896 19398 7948
rect 20714 7936 20720 7948
rect 19444 7908 20720 7936
rect 18693 7871 18751 7877
rect 18693 7868 18705 7871
rect 18196 7840 18705 7868
rect 18196 7828 18202 7840
rect 18693 7837 18705 7840
rect 18739 7837 18751 7871
rect 18693 7831 18751 7837
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7868 18935 7871
rect 19150 7868 19156 7880
rect 18923 7840 19156 7868
rect 18923 7837 18935 7840
rect 18877 7831 18935 7837
rect 19150 7828 19156 7840
rect 19208 7828 19214 7880
rect 19444 7877 19472 7908
rect 20714 7896 20720 7908
rect 20772 7896 20778 7948
rect 20898 7896 20904 7948
rect 20956 7896 20962 7948
rect 21818 7896 21824 7948
rect 21876 7936 21882 7948
rect 21876 7908 22968 7936
rect 21876 7896 21882 7908
rect 19245 7871 19303 7877
rect 19245 7837 19257 7871
rect 19291 7837 19303 7871
rect 19245 7831 19303 7837
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7837 19487 7871
rect 19429 7831 19487 7837
rect 11848 7772 14412 7800
rect 15381 7803 15439 7809
rect 11848 7760 11854 7772
rect 15381 7769 15393 7803
rect 15427 7800 15439 7803
rect 16301 7803 16359 7809
rect 16301 7800 16313 7803
rect 15427 7772 16313 7800
rect 15427 7769 15439 7772
rect 15381 7763 15439 7769
rect 16301 7769 16313 7772
rect 16347 7769 16359 7803
rect 16301 7763 16359 7769
rect 16758 7760 16764 7812
rect 16816 7760 16822 7812
rect 17770 7760 17776 7812
rect 17828 7800 17834 7812
rect 18049 7803 18107 7809
rect 18049 7800 18061 7803
rect 17828 7772 18061 7800
rect 17828 7760 17834 7772
rect 18049 7769 18061 7772
rect 18095 7800 18107 7803
rect 18966 7800 18972 7812
rect 18095 7772 18972 7800
rect 18095 7769 18107 7772
rect 18049 7763 18107 7769
rect 18966 7760 18972 7772
rect 19024 7760 19030 7812
rect 19260 7800 19288 7831
rect 20070 7828 20076 7880
rect 20128 7868 20134 7880
rect 20165 7871 20223 7877
rect 20165 7868 20177 7871
rect 20128 7840 20177 7868
rect 20128 7828 20134 7840
rect 20165 7837 20177 7840
rect 20211 7837 20223 7871
rect 20165 7831 20223 7837
rect 20346 7828 20352 7880
rect 20404 7828 20410 7880
rect 20441 7871 20499 7877
rect 20441 7837 20453 7871
rect 20487 7868 20499 7871
rect 20530 7868 20536 7880
rect 20487 7840 20536 7868
rect 20487 7837 20499 7840
rect 20441 7831 20499 7837
rect 20530 7828 20536 7840
rect 20588 7868 20594 7880
rect 21177 7871 21235 7877
rect 21177 7868 21189 7871
rect 20588 7840 21189 7868
rect 20588 7828 20594 7840
rect 21177 7837 21189 7840
rect 21223 7837 21235 7871
rect 21177 7831 21235 7837
rect 22094 7828 22100 7880
rect 22152 7828 22158 7880
rect 22189 7871 22247 7877
rect 22189 7837 22201 7871
rect 22235 7837 22247 7871
rect 22189 7831 22247 7837
rect 20622 7800 20628 7812
rect 19260 7772 20628 7800
rect 20622 7760 20628 7772
rect 20680 7760 20686 7812
rect 22204 7800 22232 7831
rect 22278 7828 22284 7880
rect 22336 7828 22342 7880
rect 22388 7877 22416 7908
rect 22373 7871 22431 7877
rect 22373 7837 22385 7871
rect 22419 7837 22431 7871
rect 22373 7831 22431 7837
rect 22462 7828 22468 7880
rect 22520 7868 22526 7880
rect 22557 7871 22615 7877
rect 22557 7868 22569 7871
rect 22520 7840 22569 7868
rect 22520 7828 22526 7840
rect 22557 7837 22569 7840
rect 22603 7837 22615 7871
rect 22557 7831 22615 7837
rect 22738 7828 22744 7880
rect 22796 7828 22802 7880
rect 22940 7877 22968 7908
rect 23014 7896 23020 7948
rect 23072 7896 23078 7948
rect 23216 7877 23244 7976
rect 23308 7936 23336 8044
rect 23382 8032 23388 8084
rect 23440 8032 23446 8084
rect 24670 8032 24676 8084
rect 24728 8032 24734 8084
rect 25498 8032 25504 8084
rect 25556 8072 25562 8084
rect 26050 8072 26056 8084
rect 25556 8044 26056 8072
rect 25556 8032 25562 8044
rect 26050 8032 26056 8044
rect 26108 8072 26114 8084
rect 26329 8075 26387 8081
rect 26108 8044 26188 8072
rect 26108 8032 26114 8044
rect 25225 8007 25283 8013
rect 25225 7973 25237 8007
rect 25271 8004 25283 8007
rect 25961 8007 26019 8013
rect 25961 8004 25973 8007
rect 25271 7976 25973 8004
rect 25271 7973 25283 7976
rect 25225 7967 25283 7973
rect 25961 7973 25973 7976
rect 26007 7973 26019 8007
rect 25961 7967 26019 7973
rect 25593 7939 25651 7945
rect 25593 7936 25605 7939
rect 23308 7908 25605 7936
rect 25593 7905 25605 7908
rect 25639 7936 25651 7939
rect 25774 7936 25780 7948
rect 25639 7908 25780 7936
rect 25639 7905 25651 7908
rect 25593 7899 25651 7905
rect 25774 7896 25780 7908
rect 25832 7896 25838 7948
rect 22925 7871 22983 7877
rect 22925 7837 22937 7871
rect 22971 7837 22983 7871
rect 22925 7831 22983 7837
rect 23109 7871 23167 7877
rect 23109 7837 23121 7871
rect 23155 7837 23167 7871
rect 23109 7831 23167 7837
rect 23201 7871 23259 7877
rect 23201 7837 23213 7871
rect 23247 7837 23259 7871
rect 23201 7831 23259 7837
rect 22204 7772 22508 7800
rect 7300 7704 8248 7732
rect 9490 7692 9496 7744
rect 9548 7692 9554 7744
rect 13814 7692 13820 7744
rect 13872 7692 13878 7744
rect 14185 7735 14243 7741
rect 14185 7701 14197 7735
rect 14231 7732 14243 7735
rect 14550 7732 14556 7744
rect 14231 7704 14556 7732
rect 14231 7701 14243 7704
rect 14185 7695 14243 7701
rect 14550 7692 14556 7704
rect 14608 7692 14614 7744
rect 15286 7692 15292 7744
rect 15344 7732 15350 7744
rect 19981 7735 20039 7741
rect 19981 7732 19993 7735
rect 15344 7704 19993 7732
rect 15344 7692 15350 7704
rect 19981 7701 19993 7704
rect 20027 7701 20039 7735
rect 19981 7695 20039 7701
rect 20070 7692 20076 7744
rect 20128 7732 20134 7744
rect 21913 7735 21971 7741
rect 21913 7732 21925 7735
rect 20128 7704 21925 7732
rect 20128 7692 20134 7704
rect 21913 7701 21925 7704
rect 21959 7701 21971 7735
rect 22480 7732 22508 7772
rect 22646 7760 22652 7812
rect 22704 7800 22710 7812
rect 23124 7800 23152 7831
rect 24118 7828 24124 7880
rect 24176 7828 24182 7880
rect 25869 7871 25927 7877
rect 25869 7837 25881 7871
rect 25915 7868 25927 7871
rect 26160 7868 26188 8044
rect 26329 8041 26341 8075
rect 26375 8072 26387 8075
rect 26418 8072 26424 8084
rect 26375 8044 26424 8072
rect 26375 8041 26387 8044
rect 26329 8035 26387 8041
rect 26418 8032 26424 8044
rect 26476 8032 26482 8084
rect 26510 8032 26516 8084
rect 26568 8072 26574 8084
rect 27249 8075 27307 8081
rect 27249 8072 27261 8075
rect 26568 8044 27261 8072
rect 26568 8032 26574 8044
rect 27249 8041 27261 8044
rect 27295 8072 27307 8075
rect 27430 8072 27436 8084
rect 27295 8044 27436 8072
rect 27295 8041 27307 8044
rect 27249 8035 27307 8041
rect 27430 8032 27436 8044
rect 27488 8032 27494 8084
rect 28258 8032 28264 8084
rect 28316 8032 28322 8084
rect 28626 8032 28632 8084
rect 28684 8032 28690 8084
rect 30193 8075 30251 8081
rect 30193 8041 30205 8075
rect 30239 8072 30251 8075
rect 30282 8072 30288 8084
rect 30239 8044 30288 8072
rect 30239 8041 30251 8044
rect 30193 8035 30251 8041
rect 30282 8032 30288 8044
rect 30340 8032 30346 8084
rect 30374 8032 30380 8084
rect 30432 8032 30438 8084
rect 30742 8032 30748 8084
rect 30800 8072 30806 8084
rect 30837 8075 30895 8081
rect 30837 8072 30849 8075
rect 30800 8044 30849 8072
rect 30800 8032 30806 8044
rect 30837 8041 30849 8044
rect 30883 8072 30895 8075
rect 31570 8072 31576 8084
rect 30883 8044 31576 8072
rect 30883 8041 30895 8044
rect 30837 8035 30895 8041
rect 31570 8032 31576 8044
rect 31628 8072 31634 8084
rect 31628 8044 35296 8072
rect 31628 8032 31634 8044
rect 26786 7964 26792 8016
rect 26844 7964 26850 8016
rect 27522 8004 27528 8016
rect 26995 7976 27528 8004
rect 26234 7896 26240 7948
rect 26292 7896 26298 7948
rect 26602 7896 26608 7948
rect 26660 7936 26666 7948
rect 26995 7936 27023 7976
rect 27522 7964 27528 7976
rect 27580 7964 27586 8016
rect 28166 7964 28172 8016
rect 28224 8004 28230 8016
rect 28445 8007 28503 8013
rect 28445 8004 28457 8007
rect 28224 7976 28457 8004
rect 28224 7964 28230 7976
rect 28445 7973 28457 7976
rect 28491 7973 28503 8007
rect 30300 8004 30328 8032
rect 35268 8004 35296 8044
rect 36170 8032 36176 8084
rect 36228 8072 36234 8084
rect 36541 8075 36599 8081
rect 36541 8072 36553 8075
rect 36228 8044 36553 8072
rect 36228 8032 36234 8044
rect 36541 8041 36553 8044
rect 36587 8041 36599 8075
rect 36541 8035 36599 8041
rect 36814 8032 36820 8084
rect 36872 8032 36878 8084
rect 35986 8004 35992 8016
rect 30300 7976 31892 8004
rect 28445 7967 28503 7973
rect 26660 7908 27023 7936
rect 26660 7896 26666 7908
rect 26988 7877 27016 7908
rect 27062 7896 27068 7948
rect 27120 7896 27126 7948
rect 27154 7896 27160 7948
rect 27212 7936 27218 7948
rect 28994 7936 29000 7948
rect 27212 7908 29000 7936
rect 27212 7896 27218 7908
rect 28994 7896 29000 7908
rect 29052 7896 29058 7948
rect 31386 7936 31392 7948
rect 30208 7908 31392 7936
rect 26329 7871 26387 7877
rect 26329 7868 26341 7871
rect 25915 7840 26096 7868
rect 26160 7840 26341 7868
rect 25915 7837 25927 7840
rect 25869 7831 25927 7837
rect 24949 7803 25007 7809
rect 22704 7772 24072 7800
rect 22704 7760 22710 7772
rect 22922 7732 22928 7744
rect 22480 7704 22928 7732
rect 21913 7695 21971 7701
rect 22922 7692 22928 7704
rect 22980 7692 22986 7744
rect 24044 7741 24072 7772
rect 24949 7769 24961 7803
rect 24995 7800 25007 7803
rect 24995 7772 25176 7800
rect 24995 7769 25007 7772
rect 24949 7763 25007 7769
rect 24029 7735 24087 7741
rect 24029 7701 24041 7735
rect 24075 7732 24087 7735
rect 24486 7732 24492 7744
rect 24075 7704 24492 7732
rect 24075 7701 24087 7704
rect 24029 7695 24087 7701
rect 24486 7692 24492 7704
rect 24544 7692 24550 7744
rect 24762 7692 24768 7744
rect 24820 7732 24826 7744
rect 24857 7735 24915 7741
rect 24857 7732 24869 7735
rect 24820 7704 24869 7732
rect 24820 7692 24826 7704
rect 24857 7701 24869 7704
rect 24903 7701 24915 7735
rect 24857 7695 24915 7701
rect 25038 7692 25044 7744
rect 25096 7692 25102 7744
rect 25148 7732 25176 7772
rect 25317 7735 25375 7741
rect 25317 7732 25329 7735
rect 25148 7704 25329 7732
rect 25317 7701 25329 7704
rect 25363 7701 25375 7735
rect 26068 7732 26096 7840
rect 26329 7837 26341 7840
rect 26375 7837 26387 7871
rect 26329 7831 26387 7837
rect 26973 7871 27031 7877
rect 26973 7837 26985 7871
rect 27019 7837 27031 7871
rect 26973 7831 27031 7837
rect 27249 7871 27307 7877
rect 27249 7837 27261 7871
rect 27295 7868 27307 7871
rect 27798 7868 27804 7880
rect 27295 7840 27804 7868
rect 27295 7837 27307 7840
rect 27249 7831 27307 7837
rect 27798 7828 27804 7840
rect 27856 7868 27862 7880
rect 28721 7871 28779 7877
rect 28721 7868 28733 7871
rect 27856 7840 28733 7868
rect 27856 7828 27862 7840
rect 28721 7837 28733 7840
rect 28767 7837 28779 7871
rect 28721 7831 28779 7837
rect 28810 7828 28816 7880
rect 28868 7828 28874 7880
rect 29178 7828 29184 7880
rect 29236 7828 29242 7880
rect 29365 7871 29423 7877
rect 29365 7837 29377 7871
rect 29411 7868 29423 7871
rect 29638 7868 29644 7880
rect 29411 7840 29644 7868
rect 29411 7837 29423 7840
rect 29365 7831 29423 7837
rect 29638 7828 29644 7840
rect 29696 7828 29702 7880
rect 29733 7871 29791 7877
rect 29733 7837 29745 7871
rect 29779 7837 29791 7871
rect 29733 7831 29791 7837
rect 28074 7760 28080 7812
rect 28132 7760 28138 7812
rect 29748 7800 29776 7831
rect 29822 7828 29828 7880
rect 29880 7828 29886 7880
rect 30208 7877 30236 7908
rect 30193 7871 30251 7877
rect 30193 7837 30205 7871
rect 30239 7837 30251 7871
rect 30193 7831 30251 7837
rect 30282 7828 30288 7880
rect 30340 7868 30346 7880
rect 30852 7877 30880 7908
rect 31386 7896 31392 7908
rect 31444 7896 31450 7948
rect 31478 7896 31484 7948
rect 31536 7896 31542 7948
rect 31864 7936 31892 7976
rect 32416 7976 33364 8004
rect 32306 7936 32312 7948
rect 31864 7908 32312 7936
rect 30561 7871 30619 7877
rect 30561 7868 30573 7871
rect 30340 7840 30573 7868
rect 30340 7828 30346 7840
rect 30561 7837 30573 7840
rect 30607 7837 30619 7871
rect 30561 7831 30619 7837
rect 30837 7871 30895 7877
rect 30837 7837 30849 7871
rect 30883 7837 30895 7871
rect 30837 7831 30895 7837
rect 31018 7828 31024 7880
rect 31076 7868 31082 7880
rect 31956 7877 31984 7908
rect 32306 7896 32312 7908
rect 32364 7896 32370 7948
rect 32416 7945 32444 7976
rect 32401 7939 32459 7945
rect 32401 7905 32413 7939
rect 32447 7905 32459 7939
rect 32401 7899 32459 7905
rect 32585 7939 32643 7945
rect 32585 7905 32597 7939
rect 32631 7936 32643 7939
rect 33042 7936 33048 7948
rect 32631 7908 33048 7936
rect 32631 7905 32643 7908
rect 32585 7899 32643 7905
rect 33042 7896 33048 7908
rect 33100 7896 33106 7948
rect 33336 7945 33364 7976
rect 35268 7976 35992 8004
rect 33321 7939 33379 7945
rect 33321 7905 33333 7939
rect 33367 7936 33379 7939
rect 33410 7936 33416 7948
rect 33367 7908 33416 7936
rect 33367 7905 33379 7908
rect 33321 7899 33379 7905
rect 33410 7896 33416 7908
rect 33468 7896 33474 7948
rect 33502 7896 33508 7948
rect 33560 7896 33566 7948
rect 34790 7896 34796 7948
rect 34848 7936 34854 7948
rect 34885 7939 34943 7945
rect 34885 7936 34897 7939
rect 34848 7908 34897 7936
rect 34848 7896 34854 7908
rect 34885 7905 34897 7908
rect 34931 7905 34943 7939
rect 34885 7899 34943 7905
rect 31205 7871 31263 7877
rect 31205 7868 31217 7871
rect 31076 7840 31217 7868
rect 31076 7828 31082 7840
rect 31205 7837 31217 7840
rect 31251 7868 31263 7871
rect 31849 7871 31907 7877
rect 31849 7868 31861 7871
rect 31251 7840 31861 7868
rect 31251 7837 31263 7840
rect 31205 7831 31263 7837
rect 31849 7837 31861 7840
rect 31895 7837 31907 7871
rect 31849 7831 31907 7837
rect 31941 7871 31999 7877
rect 31941 7837 31953 7871
rect 31987 7837 31999 7871
rect 31941 7831 31999 7837
rect 32953 7871 33011 7877
rect 32953 7837 32965 7871
rect 32999 7868 33011 7871
rect 33778 7868 33784 7880
rect 32999 7840 33784 7868
rect 32999 7837 33011 7840
rect 32953 7831 33011 7837
rect 33778 7828 33784 7840
rect 33836 7868 33842 7880
rect 33965 7871 34023 7877
rect 33965 7868 33977 7871
rect 33836 7840 33977 7868
rect 33836 7828 33842 7840
rect 33965 7837 33977 7840
rect 34011 7868 34023 7871
rect 34011 7840 34560 7868
rect 34011 7837 34023 7840
rect 33965 7831 34023 7837
rect 31036 7800 31064 7828
rect 34532 7812 34560 7840
rect 34698 7828 34704 7880
rect 34756 7868 34762 7880
rect 35268 7877 35296 7976
rect 35986 7964 35992 7976
rect 36044 8004 36050 8016
rect 36832 8004 36860 8032
rect 36044 7976 36860 8004
rect 36044 7964 36050 7976
rect 35434 7896 35440 7948
rect 35492 7936 35498 7948
rect 35805 7939 35863 7945
rect 35805 7936 35817 7939
rect 35492 7908 35817 7936
rect 35492 7896 35498 7908
rect 35805 7905 35817 7908
rect 35851 7905 35863 7939
rect 35805 7899 35863 7905
rect 36725 7939 36783 7945
rect 36725 7905 36737 7939
rect 36771 7936 36783 7939
rect 38194 7936 38200 7948
rect 36771 7908 38200 7936
rect 36771 7905 36783 7908
rect 36725 7899 36783 7905
rect 38194 7896 38200 7908
rect 38252 7896 38258 7948
rect 35253 7871 35311 7877
rect 34756 7840 34928 7868
rect 34756 7828 34762 7840
rect 28184 7772 28994 7800
rect 29748 7772 31064 7800
rect 32033 7803 32091 7809
rect 28184 7732 28212 7772
rect 26068 7704 28212 7732
rect 25317 7695 25375 7701
rect 28258 7692 28264 7744
rect 28316 7741 28322 7744
rect 28316 7735 28335 7741
rect 28323 7701 28335 7735
rect 28966 7732 28994 7772
rect 32033 7769 32045 7803
rect 32079 7769 32091 7803
rect 32033 7763 32091 7769
rect 33137 7803 33195 7809
rect 33137 7769 33149 7803
rect 33183 7800 33195 7803
rect 33318 7800 33324 7812
rect 33183 7772 33324 7800
rect 33183 7769 33195 7772
rect 33137 7763 33195 7769
rect 30834 7732 30840 7744
rect 28966 7704 30840 7732
rect 28316 7695 28335 7701
rect 28316 7692 28322 7695
rect 30834 7692 30840 7704
rect 30892 7692 30898 7744
rect 31021 7735 31079 7741
rect 31021 7701 31033 7735
rect 31067 7732 31079 7735
rect 31294 7732 31300 7744
rect 31067 7704 31300 7732
rect 31067 7701 31079 7704
rect 31021 7695 31079 7701
rect 31294 7692 31300 7704
rect 31352 7692 31358 7744
rect 32048 7732 32076 7763
rect 33318 7760 33324 7772
rect 33376 7760 33382 7812
rect 34057 7803 34115 7809
rect 34057 7800 34069 7803
rect 33796 7772 34069 7800
rect 32306 7732 32312 7744
rect 32048 7704 32312 7732
rect 32306 7692 32312 7704
rect 32364 7732 32370 7744
rect 33045 7735 33103 7741
rect 33045 7732 33057 7735
rect 32364 7704 33057 7732
rect 32364 7692 32370 7704
rect 33045 7701 33057 7704
rect 33091 7732 33103 7735
rect 33796 7732 33824 7772
rect 34057 7769 34069 7772
rect 34103 7769 34115 7803
rect 34057 7763 34115 7769
rect 33091 7704 33824 7732
rect 33873 7735 33931 7741
rect 33091 7701 33103 7704
rect 33045 7695 33103 7701
rect 33873 7701 33885 7735
rect 33919 7732 33931 7735
rect 33962 7732 33968 7744
rect 33919 7704 33968 7732
rect 33919 7701 33931 7704
rect 33873 7695 33931 7701
rect 33962 7692 33968 7704
rect 34020 7692 34026 7744
rect 34072 7732 34100 7763
rect 34514 7760 34520 7812
rect 34572 7800 34578 7812
rect 34793 7803 34851 7809
rect 34793 7800 34805 7803
rect 34572 7772 34805 7800
rect 34572 7760 34578 7772
rect 34793 7769 34805 7772
rect 34839 7769 34851 7803
rect 34900 7800 34928 7840
rect 35253 7837 35265 7871
rect 35299 7837 35311 7871
rect 35253 7831 35311 7837
rect 35345 7871 35403 7877
rect 35345 7837 35357 7871
rect 35391 7868 35403 7871
rect 36078 7868 36084 7880
rect 35391 7840 36084 7868
rect 35391 7837 35403 7840
rect 35345 7831 35403 7837
rect 35360 7800 35388 7831
rect 36078 7828 36084 7840
rect 36136 7828 36142 7880
rect 40034 7828 40040 7880
rect 40092 7868 40098 7880
rect 40129 7871 40187 7877
rect 40129 7868 40141 7871
rect 40092 7840 40141 7868
rect 40092 7828 40098 7840
rect 40129 7837 40141 7840
rect 40175 7837 40187 7871
rect 40129 7831 40187 7837
rect 34900 7772 35388 7800
rect 36449 7803 36507 7809
rect 34793 7763 34851 7769
rect 36449 7769 36461 7803
rect 36495 7769 36507 7803
rect 36449 7763 36507 7769
rect 34606 7732 34612 7744
rect 34072 7704 34612 7732
rect 34606 7692 34612 7704
rect 34664 7692 34670 7744
rect 35066 7692 35072 7744
rect 35124 7732 35130 7744
rect 36354 7732 36360 7744
rect 35124 7704 36360 7732
rect 35124 7692 35130 7704
rect 36354 7692 36360 7704
rect 36412 7732 36418 7744
rect 36464 7732 36492 7763
rect 36998 7760 37004 7812
rect 37056 7760 37062 7812
rect 37458 7760 37464 7812
rect 37516 7760 37522 7812
rect 38749 7803 38807 7809
rect 38749 7800 38761 7803
rect 38304 7772 38761 7800
rect 36412 7704 36492 7732
rect 36412 7692 36418 7704
rect 37274 7692 37280 7744
rect 37332 7732 37338 7744
rect 38304 7732 38332 7772
rect 38749 7769 38761 7772
rect 38795 7769 38807 7803
rect 38749 7763 38807 7769
rect 37332 7704 38332 7732
rect 37332 7692 37338 7704
rect 39022 7692 39028 7744
rect 39080 7732 39086 7744
rect 39945 7735 40003 7741
rect 39945 7732 39957 7735
rect 39080 7704 39957 7732
rect 39080 7692 39086 7704
rect 39945 7701 39957 7704
rect 39991 7701 40003 7735
rect 39945 7695 40003 7701
rect 1104 7642 40572 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 40572 7642
rect 1104 7568 40572 7590
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 8021 7531 8079 7537
rect 8021 7528 8033 7531
rect 7340 7500 8033 7528
rect 7340 7488 7346 7500
rect 8021 7497 8033 7500
rect 8067 7528 8079 7531
rect 8662 7528 8668 7540
rect 8067 7500 8668 7528
rect 8067 7497 8079 7500
rect 8021 7491 8079 7497
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 9232 7500 11008 7528
rect 8202 7352 8208 7404
rect 8260 7352 8266 7404
rect 8294 7352 8300 7404
rect 8352 7352 8358 7404
rect 9232 7401 9260 7500
rect 10980 7472 11008 7500
rect 12066 7488 12072 7540
rect 12124 7528 12130 7540
rect 12342 7528 12348 7540
rect 12124 7500 12348 7528
rect 12124 7488 12130 7500
rect 12342 7488 12348 7500
rect 12400 7488 12406 7540
rect 12434 7488 12440 7540
rect 12492 7488 12498 7540
rect 14274 7488 14280 7540
rect 14332 7528 14338 7540
rect 14461 7531 14519 7537
rect 14461 7528 14473 7531
rect 14332 7500 14473 7528
rect 14332 7488 14338 7500
rect 14461 7497 14473 7500
rect 14507 7497 14519 7531
rect 14461 7491 14519 7497
rect 14550 7488 14556 7540
rect 14608 7528 14614 7540
rect 14608 7500 15424 7528
rect 14608 7488 14614 7500
rect 9490 7420 9496 7472
rect 9548 7420 9554 7472
rect 10962 7420 10968 7472
rect 11020 7460 11026 7472
rect 12452 7460 12480 7488
rect 14366 7460 14372 7472
rect 11020 7432 12756 7460
rect 14214 7432 14372 7460
rect 11020 7420 11026 7432
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7361 9275 7395
rect 9217 7355 9275 7361
rect 10594 7352 10600 7404
rect 10652 7352 10658 7404
rect 11977 7395 12035 7401
rect 11977 7361 11989 7395
rect 12023 7361 12035 7395
rect 11977 7355 12035 7361
rect 12437 7395 12495 7401
rect 12437 7361 12449 7395
rect 12483 7392 12495 7395
rect 12618 7392 12624 7404
rect 12483 7364 12624 7392
rect 12483 7361 12495 7364
rect 12437 7355 12495 7361
rect 4706 7284 4712 7336
rect 4764 7324 4770 7336
rect 10612 7324 10640 7352
rect 4764 7296 10640 7324
rect 4764 7284 4770 7296
rect 10686 7284 10692 7336
rect 10744 7324 10750 7336
rect 10965 7327 11023 7333
rect 10965 7324 10977 7327
rect 10744 7296 10977 7324
rect 10744 7284 10750 7296
rect 10965 7293 10977 7296
rect 11011 7293 11023 7327
rect 11992 7324 12020 7355
rect 12618 7352 12624 7364
rect 12676 7352 12682 7404
rect 12728 7401 12756 7432
rect 14366 7420 14372 7432
rect 14424 7420 14430 7472
rect 15105 7463 15163 7469
rect 15105 7460 15117 7463
rect 14752 7432 15117 7460
rect 14752 7401 14780 7432
rect 15105 7429 15117 7432
rect 15151 7429 15163 7463
rect 15105 7423 15163 7429
rect 12713 7395 12771 7401
rect 12713 7361 12725 7395
rect 12759 7361 12771 7395
rect 12713 7355 12771 7361
rect 14737 7395 14795 7401
rect 14737 7361 14749 7395
rect 14783 7361 14795 7395
rect 14737 7355 14795 7361
rect 15286 7352 15292 7404
rect 15344 7352 15350 7404
rect 15396 7401 15424 7500
rect 15930 7488 15936 7540
rect 15988 7528 15994 7540
rect 16761 7531 16819 7537
rect 16761 7528 16773 7531
rect 15988 7500 16773 7528
rect 15988 7488 15994 7500
rect 16761 7497 16773 7500
rect 16807 7497 16819 7531
rect 16761 7491 16819 7497
rect 17497 7531 17555 7537
rect 17497 7497 17509 7531
rect 17543 7528 17555 7531
rect 17586 7528 17592 7540
rect 17543 7500 17592 7528
rect 17543 7497 17555 7500
rect 17497 7491 17555 7497
rect 17586 7488 17592 7500
rect 17644 7488 17650 7540
rect 17954 7488 17960 7540
rect 18012 7488 18018 7540
rect 18125 7531 18183 7537
rect 18125 7497 18137 7531
rect 18171 7528 18183 7531
rect 20438 7528 20444 7540
rect 18171 7500 20444 7528
rect 18171 7497 18183 7500
rect 18125 7491 18183 7497
rect 20438 7488 20444 7500
rect 20496 7488 20502 7540
rect 21266 7488 21272 7540
rect 21324 7528 21330 7540
rect 21324 7500 21680 7528
rect 21324 7488 21330 7500
rect 16482 7420 16488 7472
rect 16540 7420 16546 7472
rect 17313 7463 17371 7469
rect 17313 7429 17325 7463
rect 17359 7460 17371 7463
rect 17770 7460 17776 7472
rect 17359 7432 17776 7460
rect 17359 7429 17371 7432
rect 17313 7423 17371 7429
rect 17770 7420 17776 7432
rect 17828 7420 17834 7472
rect 18325 7463 18383 7469
rect 18325 7429 18337 7463
rect 18371 7429 18383 7463
rect 18325 7423 18383 7429
rect 15381 7395 15439 7401
rect 15381 7361 15393 7395
rect 15427 7392 15439 7395
rect 16298 7392 16304 7404
rect 15427 7364 16304 7392
rect 15427 7361 15439 7364
rect 15381 7355 15439 7361
rect 16298 7352 16304 7364
rect 16356 7352 16362 7404
rect 16669 7395 16727 7401
rect 16669 7361 16681 7395
rect 16715 7392 16727 7395
rect 16758 7392 16764 7404
rect 16715 7364 16764 7392
rect 16715 7361 16727 7364
rect 16669 7355 16727 7361
rect 16758 7352 16764 7364
rect 16816 7352 16822 7404
rect 16853 7395 16911 7401
rect 16853 7361 16865 7395
rect 16899 7392 16911 7395
rect 17218 7392 17224 7404
rect 16899 7364 17224 7392
rect 16899 7361 16911 7364
rect 16853 7355 16911 7361
rect 17218 7352 17224 7364
rect 17276 7352 17282 7404
rect 18230 7352 18236 7404
rect 18288 7392 18294 7404
rect 18340 7392 18368 7423
rect 18966 7420 18972 7472
rect 19024 7460 19030 7472
rect 20806 7460 20812 7472
rect 19024 7432 20812 7460
rect 19024 7420 19030 7432
rect 20806 7420 20812 7432
rect 20864 7420 20870 7472
rect 21652 7469 21680 7500
rect 22002 7488 22008 7540
rect 22060 7488 22066 7540
rect 22186 7537 22192 7540
rect 22173 7531 22192 7537
rect 22173 7497 22185 7531
rect 22244 7528 22250 7540
rect 22244 7500 23520 7528
rect 22173 7491 22192 7497
rect 22186 7488 22192 7491
rect 22244 7488 22250 7500
rect 21637 7463 21695 7469
rect 21407 7429 21465 7435
rect 18288 7364 18368 7392
rect 18417 7395 18475 7401
rect 18288 7352 18294 7364
rect 18417 7361 18429 7395
rect 18463 7392 18475 7395
rect 18782 7392 18788 7404
rect 18463 7364 18788 7392
rect 18463 7361 18475 7364
rect 18417 7355 18475 7361
rect 18782 7352 18788 7364
rect 18840 7352 18846 7404
rect 20714 7352 20720 7404
rect 20772 7392 20778 7404
rect 20993 7395 21051 7401
rect 20993 7392 21005 7395
rect 20772 7364 21005 7392
rect 20772 7352 20778 7364
rect 20993 7361 21005 7364
rect 21039 7361 21051 7395
rect 20993 7355 21051 7361
rect 12526 7324 12532 7336
rect 11992 7296 12532 7324
rect 10965 7287 11023 7293
rect 12526 7284 12532 7296
rect 12584 7284 12590 7336
rect 12986 7284 12992 7336
rect 13044 7284 13050 7336
rect 13998 7284 14004 7336
rect 14056 7324 14062 7336
rect 14642 7324 14648 7336
rect 14056 7296 14648 7324
rect 14056 7284 14062 7296
rect 14642 7284 14648 7296
rect 14700 7324 14706 7336
rect 15013 7327 15071 7333
rect 15013 7324 15025 7327
rect 14700 7296 15025 7324
rect 14700 7284 14706 7296
rect 15013 7293 15025 7296
rect 15059 7293 15071 7327
rect 15013 7287 15071 7293
rect 15105 7327 15163 7333
rect 15105 7293 15117 7327
rect 15151 7293 15163 7327
rect 15105 7287 15163 7293
rect 15749 7327 15807 7333
rect 15749 7293 15761 7327
rect 15795 7324 15807 7327
rect 15930 7324 15936 7336
rect 15795 7296 15936 7324
rect 15795 7293 15807 7296
rect 15749 7287 15807 7293
rect 12529 7191 12587 7197
rect 12529 7157 12541 7191
rect 12575 7188 12587 7191
rect 14182 7188 14188 7200
rect 12575 7160 14188 7188
rect 12575 7157 12587 7160
rect 12529 7151 12587 7157
rect 14182 7148 14188 7160
rect 14240 7148 14246 7200
rect 14550 7148 14556 7200
rect 14608 7148 14614 7200
rect 14734 7148 14740 7200
rect 14792 7188 14798 7200
rect 14921 7191 14979 7197
rect 14921 7188 14933 7191
rect 14792 7160 14933 7188
rect 14792 7148 14798 7160
rect 14921 7157 14933 7160
rect 14967 7188 14979 7191
rect 15120 7188 15148 7287
rect 15930 7284 15936 7296
rect 15988 7284 15994 7336
rect 16574 7284 16580 7336
rect 16632 7324 16638 7336
rect 18509 7327 18567 7333
rect 18509 7324 18521 7327
rect 16632 7296 18521 7324
rect 16632 7284 16638 7296
rect 18509 7293 18521 7296
rect 18555 7293 18567 7327
rect 18509 7287 18567 7293
rect 20809 7327 20867 7333
rect 20809 7293 20821 7327
rect 20855 7293 20867 7327
rect 20809 7287 20867 7293
rect 16666 7216 16672 7268
rect 16724 7256 16730 7268
rect 16945 7259 17003 7265
rect 16945 7256 16957 7259
rect 16724 7228 16957 7256
rect 16724 7216 16730 7228
rect 16945 7225 16957 7228
rect 16991 7225 17003 7259
rect 16945 7219 17003 7225
rect 17678 7216 17684 7268
rect 17736 7256 17742 7268
rect 20625 7259 20683 7265
rect 20625 7256 20637 7259
rect 17736 7228 20637 7256
rect 17736 7216 17742 7228
rect 20625 7225 20637 7228
rect 20671 7225 20683 7259
rect 20824 7256 20852 7287
rect 20898 7284 20904 7336
rect 20956 7284 20962 7336
rect 21008 7324 21036 7355
rect 21082 7352 21088 7404
rect 21140 7352 21146 7404
rect 21407 7395 21419 7429
rect 21453 7426 21465 7429
rect 21637 7429 21649 7463
rect 21683 7429 21695 7463
rect 21453 7395 21475 7426
rect 21637 7423 21695 7429
rect 22370 7420 22376 7472
rect 22428 7420 22434 7472
rect 23492 7460 23520 7500
rect 24762 7488 24768 7540
rect 24820 7528 24826 7540
rect 24949 7531 25007 7537
rect 24949 7528 24961 7531
rect 24820 7500 24961 7528
rect 24820 7488 24826 7500
rect 24949 7497 24961 7500
rect 24995 7497 25007 7531
rect 24949 7491 25007 7497
rect 25038 7488 25044 7540
rect 25096 7488 25102 7540
rect 26326 7488 26332 7540
rect 26384 7528 26390 7540
rect 27433 7531 27491 7537
rect 27433 7528 27445 7531
rect 26384 7500 27445 7528
rect 26384 7488 26390 7500
rect 27433 7497 27445 7500
rect 27479 7497 27491 7531
rect 27433 7491 27491 7497
rect 29362 7488 29368 7540
rect 29420 7528 29426 7540
rect 29641 7531 29699 7537
rect 29641 7528 29653 7531
rect 29420 7500 29653 7528
rect 29420 7488 29426 7500
rect 29641 7497 29653 7500
rect 29687 7528 29699 7531
rect 30190 7528 30196 7540
rect 29687 7500 30196 7528
rect 29687 7497 29699 7500
rect 29641 7491 29699 7497
rect 30190 7488 30196 7500
rect 30248 7488 30254 7540
rect 30282 7488 30288 7540
rect 30340 7528 30346 7540
rect 31297 7531 31355 7537
rect 31297 7528 31309 7531
rect 30340 7500 31309 7528
rect 30340 7488 30346 7500
rect 31297 7497 31309 7500
rect 31343 7497 31355 7531
rect 31297 7491 31355 7497
rect 32401 7531 32459 7537
rect 32401 7497 32413 7531
rect 32447 7528 32459 7531
rect 33410 7528 33416 7540
rect 32447 7500 33416 7528
rect 32447 7497 32459 7500
rect 32401 7491 32459 7497
rect 33410 7488 33416 7500
rect 33468 7528 33474 7540
rect 33873 7531 33931 7537
rect 33873 7528 33885 7531
rect 33468 7500 33885 7528
rect 33468 7488 33474 7500
rect 33873 7497 33885 7500
rect 33919 7528 33931 7531
rect 34698 7528 34704 7540
rect 33919 7500 34704 7528
rect 33919 7497 33931 7500
rect 33873 7491 33931 7497
rect 34698 7488 34704 7500
rect 34756 7488 34762 7540
rect 37369 7531 37427 7537
rect 37369 7497 37381 7531
rect 37415 7528 37427 7531
rect 37734 7528 37740 7540
rect 37415 7500 37740 7528
rect 37415 7497 37427 7500
rect 37369 7491 37427 7497
rect 37734 7488 37740 7500
rect 37792 7488 37798 7540
rect 39942 7488 39948 7540
rect 40000 7528 40006 7540
rect 40037 7531 40095 7537
rect 40037 7528 40049 7531
rect 40000 7500 40049 7528
rect 40000 7488 40006 7500
rect 40037 7497 40049 7500
rect 40083 7497 40095 7531
rect 40037 7491 40095 7497
rect 26237 7463 26295 7469
rect 26237 7460 26249 7463
rect 23492 7432 26249 7460
rect 26237 7429 26249 7432
rect 26283 7429 26295 7463
rect 26237 7423 26295 7429
rect 29546 7420 29552 7472
rect 29604 7420 29610 7472
rect 31113 7463 31171 7469
rect 31113 7429 31125 7463
rect 31159 7460 31171 7463
rect 31386 7460 31392 7472
rect 31159 7432 31392 7460
rect 31159 7429 31171 7432
rect 31113 7423 31171 7429
rect 31386 7420 31392 7432
rect 31444 7420 31450 7472
rect 38470 7460 38476 7472
rect 31726 7432 38476 7460
rect 21407 7392 21475 7395
rect 23290 7392 23296 7404
rect 21407 7389 23296 7392
rect 21447 7364 23296 7389
rect 21266 7324 21272 7336
rect 21008 7296 21272 7324
rect 21266 7284 21272 7296
rect 21324 7284 21330 7336
rect 21447 7256 21475 7364
rect 23290 7352 23296 7364
rect 23348 7352 23354 7404
rect 24302 7352 24308 7404
rect 24360 7392 24366 7404
rect 24397 7395 24455 7401
rect 24397 7392 24409 7395
rect 24360 7364 24409 7392
rect 24360 7352 24366 7364
rect 24397 7361 24409 7364
rect 24443 7361 24455 7395
rect 24397 7355 24455 7361
rect 24486 7352 24492 7404
rect 24544 7392 24550 7404
rect 25593 7395 25651 7401
rect 25593 7392 25605 7395
rect 24544 7364 25605 7392
rect 24544 7352 24550 7364
rect 25593 7361 25605 7364
rect 25639 7361 25651 7395
rect 25593 7355 25651 7361
rect 26510 7352 26516 7404
rect 26568 7352 26574 7404
rect 26602 7352 26608 7404
rect 26660 7352 26666 7404
rect 26973 7395 27031 7401
rect 26973 7361 26985 7395
rect 27019 7392 27031 7395
rect 27062 7392 27068 7404
rect 27019 7364 27068 7392
rect 27019 7361 27031 7364
rect 26973 7355 27031 7361
rect 27062 7352 27068 7364
rect 27120 7352 27126 7404
rect 27341 7395 27399 7401
rect 27341 7392 27353 7395
rect 27172 7364 27353 7392
rect 24673 7327 24731 7333
rect 24673 7293 24685 7327
rect 24719 7293 24731 7327
rect 24673 7287 24731 7293
rect 20824 7228 21475 7256
rect 20625 7219 20683 7225
rect 24394 7216 24400 7268
rect 24452 7256 24458 7268
rect 24688 7256 24716 7287
rect 25314 7284 25320 7336
rect 25372 7284 25378 7336
rect 26421 7327 26479 7333
rect 26421 7293 26433 7327
rect 26467 7293 26479 7327
rect 26421 7287 26479 7293
rect 26697 7327 26755 7333
rect 26697 7293 26709 7327
rect 26743 7324 26755 7327
rect 27172 7324 27200 7364
rect 27341 7361 27353 7364
rect 27387 7361 27399 7395
rect 27341 7355 27399 7361
rect 27430 7352 27436 7404
rect 27488 7392 27494 7404
rect 27525 7395 27583 7401
rect 27525 7392 27537 7395
rect 27488 7364 27537 7392
rect 27488 7352 27494 7364
rect 27525 7361 27537 7364
rect 27571 7361 27583 7395
rect 27525 7355 27583 7361
rect 27614 7352 27620 7404
rect 27672 7392 27678 7404
rect 27801 7395 27859 7401
rect 27801 7392 27813 7395
rect 27672 7364 27813 7392
rect 27672 7352 27678 7364
rect 27801 7361 27813 7364
rect 27847 7361 27859 7395
rect 27801 7355 27859 7361
rect 29178 7352 29184 7404
rect 29236 7392 29242 7404
rect 30650 7392 30656 7404
rect 29236 7364 30656 7392
rect 29236 7352 29242 7364
rect 30650 7352 30656 7364
rect 30708 7352 30714 7404
rect 31018 7352 31024 7404
rect 31076 7392 31082 7404
rect 31205 7395 31263 7401
rect 31205 7392 31217 7395
rect 31076 7364 31217 7392
rect 31076 7352 31082 7364
rect 31205 7361 31217 7364
rect 31251 7361 31263 7395
rect 31205 7355 31263 7361
rect 31726 7336 31754 7432
rect 32398 7352 32404 7404
rect 32456 7392 32462 7404
rect 32769 7395 32827 7401
rect 32769 7392 32781 7395
rect 32456 7364 32781 7392
rect 32456 7352 32462 7364
rect 32769 7361 32781 7364
rect 32815 7361 32827 7395
rect 32769 7355 32827 7361
rect 33778 7352 33784 7404
rect 33836 7352 33842 7404
rect 33962 7352 33968 7404
rect 34020 7352 34026 7404
rect 34330 7352 34336 7404
rect 34388 7352 34394 7404
rect 34517 7395 34575 7401
rect 34517 7361 34529 7395
rect 34563 7392 34575 7395
rect 34606 7392 34612 7404
rect 34563 7364 34612 7392
rect 34563 7361 34575 7364
rect 34517 7355 34575 7361
rect 34606 7352 34612 7364
rect 34664 7352 34670 7404
rect 35066 7392 35072 7404
rect 34716 7364 35072 7392
rect 26743 7296 27200 7324
rect 26743 7293 26755 7296
rect 26697 7287 26755 7293
rect 24452 7228 24716 7256
rect 26436 7256 26464 7287
rect 27062 7256 27068 7268
rect 26436 7228 27068 7256
rect 24452 7216 24458 7228
rect 27062 7216 27068 7228
rect 27120 7216 27126 7268
rect 27172 7256 27200 7296
rect 27246 7284 27252 7336
rect 27304 7324 27310 7336
rect 31294 7324 31300 7336
rect 27304 7296 31300 7324
rect 27304 7284 27310 7296
rect 31294 7284 31300 7296
rect 31352 7284 31358 7336
rect 31570 7284 31576 7336
rect 31628 7284 31634 7336
rect 31662 7284 31668 7336
rect 31720 7296 31754 7336
rect 32306 7333 32312 7336
rect 32284 7327 32312 7333
rect 31720 7284 31726 7296
rect 32284 7293 32296 7327
rect 32284 7287 32312 7293
rect 32306 7284 32312 7287
rect 32364 7284 32370 7336
rect 32493 7327 32551 7333
rect 32493 7293 32505 7327
rect 32539 7324 32551 7327
rect 33796 7324 33824 7352
rect 32539 7296 33824 7324
rect 32539 7293 32551 7296
rect 32493 7287 32551 7293
rect 34054 7284 34060 7336
rect 34112 7324 34118 7336
rect 34716 7324 34744 7364
rect 35066 7352 35072 7364
rect 35124 7392 35130 7404
rect 35253 7395 35311 7401
rect 35253 7392 35265 7395
rect 35124 7364 35265 7392
rect 35124 7352 35130 7364
rect 35253 7361 35265 7364
rect 35299 7361 35311 7395
rect 35253 7355 35311 7361
rect 35434 7352 35440 7404
rect 35492 7352 35498 7404
rect 35805 7395 35863 7401
rect 35805 7361 35817 7395
rect 35851 7392 35863 7395
rect 35986 7392 35992 7404
rect 35851 7364 35992 7392
rect 35851 7361 35863 7364
rect 35805 7355 35863 7361
rect 35986 7352 35992 7364
rect 36044 7352 36050 7404
rect 37274 7352 37280 7404
rect 37332 7352 37338 7404
rect 38304 7401 38332 7432
rect 38470 7420 38476 7432
rect 38528 7420 38534 7472
rect 38565 7463 38623 7469
rect 38565 7429 38577 7463
rect 38611 7460 38623 7463
rect 38654 7460 38660 7472
rect 38611 7432 38660 7460
rect 38611 7429 38623 7432
rect 38565 7423 38623 7429
rect 38654 7420 38660 7432
rect 38712 7420 38718 7472
rect 39022 7420 39028 7472
rect 39080 7420 39086 7472
rect 37461 7395 37519 7401
rect 37461 7361 37473 7395
rect 37507 7361 37519 7395
rect 37461 7355 37519 7361
rect 38289 7395 38347 7401
rect 38289 7361 38301 7395
rect 38335 7361 38347 7395
rect 38289 7355 38347 7361
rect 34112 7296 34744 7324
rect 35161 7327 35219 7333
rect 34112 7284 34118 7296
rect 35161 7293 35173 7327
rect 35207 7324 35219 7327
rect 35342 7324 35348 7336
rect 35207 7296 35348 7324
rect 35207 7293 35219 7296
rect 35161 7287 35219 7293
rect 27798 7256 27804 7268
rect 27172 7228 27804 7256
rect 27798 7216 27804 7228
rect 27856 7216 27862 7268
rect 28258 7216 28264 7268
rect 28316 7256 28322 7268
rect 34885 7259 34943 7265
rect 28316 7228 34432 7256
rect 28316 7216 28322 7228
rect 15562 7188 15568 7200
rect 14967 7160 15568 7188
rect 14967 7157 14979 7160
rect 14921 7151 14979 7157
rect 15562 7148 15568 7160
rect 15620 7188 15626 7200
rect 17310 7188 17316 7200
rect 15620 7160 17316 7188
rect 15620 7148 15626 7160
rect 17310 7148 17316 7160
rect 17368 7148 17374 7200
rect 18138 7148 18144 7200
rect 18196 7148 18202 7200
rect 18414 7148 18420 7200
rect 18472 7148 18478 7200
rect 18785 7191 18843 7197
rect 18785 7157 18797 7191
rect 18831 7188 18843 7191
rect 19334 7188 19340 7200
rect 18831 7160 19340 7188
rect 18831 7157 18843 7160
rect 18785 7151 18843 7157
rect 19334 7148 19340 7160
rect 19392 7148 19398 7200
rect 20714 7148 20720 7200
rect 20772 7188 20778 7200
rect 21269 7191 21327 7197
rect 21269 7188 21281 7191
rect 20772 7160 21281 7188
rect 20772 7148 20778 7160
rect 21269 7157 21281 7160
rect 21315 7157 21327 7191
rect 21269 7151 21327 7157
rect 21450 7148 21456 7200
rect 21508 7148 21514 7200
rect 22189 7191 22247 7197
rect 22189 7157 22201 7191
rect 22235 7188 22247 7191
rect 22554 7188 22560 7200
rect 22235 7160 22560 7188
rect 22235 7157 22247 7160
rect 22189 7151 22247 7157
rect 22554 7148 22560 7160
rect 22612 7148 22618 7200
rect 24765 7191 24823 7197
rect 24765 7157 24777 7191
rect 24811 7188 24823 7191
rect 25225 7191 25283 7197
rect 25225 7188 25237 7191
rect 24811 7160 25237 7188
rect 24811 7157 24823 7160
rect 24765 7151 24823 7157
rect 25225 7157 25237 7160
rect 25271 7188 25283 7191
rect 25498 7188 25504 7200
rect 25271 7160 25504 7188
rect 25271 7157 25283 7160
rect 25225 7151 25283 7157
rect 25498 7148 25504 7160
rect 25556 7188 25562 7200
rect 27982 7188 27988 7200
rect 25556 7160 27988 7188
rect 25556 7148 25562 7160
rect 27982 7148 27988 7160
rect 28040 7188 28046 7200
rect 28810 7188 28816 7200
rect 28040 7160 28816 7188
rect 28040 7148 28046 7160
rect 28810 7148 28816 7160
rect 28868 7148 28874 7200
rect 30929 7191 30987 7197
rect 30929 7157 30941 7191
rect 30975 7188 30987 7191
rect 31202 7188 31208 7200
rect 30975 7160 31208 7188
rect 30975 7157 30987 7160
rect 30929 7151 30987 7157
rect 31202 7148 31208 7160
rect 31260 7148 31266 7200
rect 31294 7148 31300 7200
rect 31352 7188 31358 7200
rect 32125 7191 32183 7197
rect 32125 7188 32137 7191
rect 31352 7160 32137 7188
rect 31352 7148 31358 7160
rect 32125 7157 32137 7160
rect 32171 7157 32183 7191
rect 34404 7188 34432 7228
rect 34885 7225 34897 7259
rect 34931 7256 34943 7259
rect 35066 7256 35072 7268
rect 34931 7228 35072 7256
rect 34931 7225 34943 7228
rect 34885 7219 34943 7225
rect 35066 7216 35072 7228
rect 35124 7216 35130 7268
rect 35176 7188 35204 7287
rect 35342 7284 35348 7296
rect 35400 7284 35406 7336
rect 35526 7284 35532 7336
rect 35584 7324 35590 7336
rect 37476 7324 37504 7355
rect 35584 7296 37504 7324
rect 35584 7284 35590 7296
rect 34404 7160 35204 7188
rect 32125 7151 32183 7157
rect 37458 7148 37464 7200
rect 37516 7188 37522 7200
rect 39022 7188 39028 7200
rect 37516 7160 39028 7188
rect 37516 7148 37522 7160
rect 39022 7148 39028 7160
rect 39080 7148 39086 7200
rect 1104 7098 40572 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 40572 7098
rect 1104 7024 40572 7046
rect 12345 6987 12403 6993
rect 12345 6953 12357 6987
rect 12391 6984 12403 6987
rect 12710 6984 12716 6996
rect 12391 6956 12716 6984
rect 12391 6953 12403 6956
rect 12345 6947 12403 6953
rect 12710 6944 12716 6956
rect 12768 6944 12774 6996
rect 12986 6944 12992 6996
rect 13044 6984 13050 6996
rect 13265 6987 13323 6993
rect 13265 6984 13277 6987
rect 13044 6956 13277 6984
rect 13044 6944 13050 6956
rect 13265 6953 13277 6956
rect 13311 6953 13323 6987
rect 13265 6947 13323 6953
rect 14200 6956 16712 6984
rect 14200 6928 14228 6956
rect 13464 6888 13952 6916
rect 11609 6851 11667 6857
rect 11609 6817 11621 6851
rect 11655 6848 11667 6851
rect 12161 6851 12219 6857
rect 12161 6848 12173 6851
rect 11655 6820 12173 6848
rect 11655 6817 11667 6820
rect 11609 6811 11667 6817
rect 12161 6817 12173 6820
rect 12207 6848 12219 6851
rect 12894 6848 12900 6860
rect 12207 6820 12900 6848
rect 12207 6817 12219 6820
rect 12161 6811 12219 6817
rect 12894 6808 12900 6820
rect 12952 6808 12958 6860
rect 13464 6857 13492 6888
rect 13449 6851 13507 6857
rect 13449 6817 13461 6851
rect 13495 6817 13507 6851
rect 13449 6811 13507 6817
rect 13541 6851 13599 6857
rect 13541 6817 13553 6851
rect 13587 6848 13599 6851
rect 13814 6848 13820 6860
rect 13587 6820 13820 6848
rect 13587 6817 13599 6820
rect 13541 6811 13599 6817
rect 13814 6808 13820 6820
rect 13872 6808 13878 6860
rect 13924 6848 13952 6888
rect 14182 6876 14188 6928
rect 14240 6876 14246 6928
rect 14366 6876 14372 6928
rect 14424 6916 14430 6928
rect 15378 6916 15384 6928
rect 14424 6888 15384 6916
rect 14424 6876 14430 6888
rect 15378 6876 15384 6888
rect 15436 6876 15442 6928
rect 15657 6919 15715 6925
rect 15657 6885 15669 6919
rect 15703 6916 15715 6919
rect 15703 6888 15792 6916
rect 15703 6885 15715 6888
rect 15657 6879 15715 6885
rect 14921 6851 14979 6857
rect 14921 6848 14933 6851
rect 13924 6820 14933 6848
rect 14921 6817 14933 6820
rect 14967 6817 14979 6851
rect 14921 6811 14979 6817
rect 15102 6808 15108 6860
rect 15160 6848 15166 6860
rect 15160 6820 15516 6848
rect 15160 6808 15166 6820
rect 11514 6740 11520 6792
rect 11572 6740 11578 6792
rect 11790 6740 11796 6792
rect 11848 6740 11854 6792
rect 11974 6740 11980 6792
rect 12032 6780 12038 6792
rect 12250 6780 12256 6792
rect 12032 6752 12256 6780
rect 12032 6740 12038 6752
rect 12250 6740 12256 6752
rect 12308 6780 12314 6792
rect 12345 6783 12403 6789
rect 12345 6780 12357 6783
rect 12308 6752 12357 6780
rect 12308 6740 12314 6752
rect 12345 6749 12357 6752
rect 12391 6749 12403 6783
rect 12345 6743 12403 6749
rect 12526 6740 12532 6792
rect 12584 6780 12590 6792
rect 13630 6780 13636 6792
rect 12584 6752 13636 6780
rect 12584 6740 12590 6752
rect 13630 6740 13636 6752
rect 13688 6740 13694 6792
rect 13725 6783 13783 6789
rect 13725 6749 13737 6783
rect 13771 6780 13783 6783
rect 14550 6780 14556 6792
rect 13771 6752 14556 6780
rect 13771 6749 13783 6752
rect 13725 6743 13783 6749
rect 14550 6740 14556 6752
rect 14608 6740 14614 6792
rect 14737 6783 14795 6789
rect 14737 6749 14749 6783
rect 14783 6780 14795 6783
rect 15286 6780 15292 6792
rect 14783 6752 15292 6780
rect 14783 6749 14795 6752
rect 14737 6743 14795 6749
rect 15286 6740 15292 6752
rect 15344 6740 15350 6792
rect 15488 6789 15516 6820
rect 15562 6808 15568 6860
rect 15620 6848 15626 6860
rect 15764 6848 15792 6888
rect 16574 6848 16580 6860
rect 15620 6820 15700 6848
rect 15764 6820 16580 6848
rect 15620 6808 15626 6820
rect 15672 6789 15700 6820
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 16684 6848 16712 6956
rect 17126 6944 17132 6996
rect 17184 6984 17190 6996
rect 20530 6984 20536 6996
rect 17184 6956 20536 6984
rect 17184 6944 17190 6956
rect 20530 6944 20536 6956
rect 20588 6944 20594 6996
rect 20622 6944 20628 6996
rect 20680 6984 20686 6996
rect 24210 6984 24216 6996
rect 20680 6956 24216 6984
rect 20680 6944 20686 6956
rect 24210 6944 24216 6956
rect 24268 6944 24274 6996
rect 33870 6944 33876 6996
rect 33928 6984 33934 6996
rect 35526 6984 35532 6996
rect 33928 6956 35532 6984
rect 33928 6944 33934 6956
rect 19610 6876 19616 6928
rect 19668 6916 19674 6928
rect 21177 6919 21235 6925
rect 21177 6916 21189 6919
rect 19668 6888 21189 6916
rect 19668 6876 19674 6888
rect 21177 6885 21189 6888
rect 21223 6916 21235 6919
rect 21450 6916 21456 6928
rect 21223 6888 21456 6916
rect 21223 6885 21235 6888
rect 21177 6879 21235 6885
rect 21450 6876 21456 6888
rect 21508 6876 21514 6928
rect 22278 6876 22284 6928
rect 22336 6916 22342 6928
rect 28258 6916 28264 6928
rect 22336 6888 28264 6916
rect 22336 6876 22342 6888
rect 28258 6876 28264 6888
rect 28316 6876 28322 6928
rect 33980 6925 34008 6956
rect 35526 6944 35532 6956
rect 35584 6944 35590 6996
rect 36354 6944 36360 6996
rect 36412 6944 36418 6996
rect 37274 6984 37280 6996
rect 36832 6956 37280 6984
rect 30377 6919 30435 6925
rect 30377 6885 30389 6919
rect 30423 6885 30435 6919
rect 30377 6879 30435 6885
rect 33965 6919 34023 6925
rect 33965 6885 33977 6919
rect 34011 6885 34023 6919
rect 36832 6916 36860 6956
rect 37274 6944 37280 6956
rect 37332 6944 37338 6996
rect 37366 6944 37372 6996
rect 37424 6984 37430 6996
rect 37841 6987 37899 6993
rect 37841 6984 37853 6987
rect 37424 6956 37853 6984
rect 37424 6944 37430 6956
rect 37841 6953 37853 6956
rect 37887 6953 37899 6987
rect 37841 6947 37899 6953
rect 33965 6879 34023 6885
rect 34256 6888 36860 6916
rect 17221 6851 17279 6857
rect 17221 6848 17233 6851
rect 16684 6820 17233 6848
rect 17221 6817 17233 6820
rect 17267 6817 17279 6851
rect 17221 6811 17279 6817
rect 17405 6851 17463 6857
rect 17405 6817 17417 6851
rect 17451 6848 17463 6851
rect 18874 6848 18880 6860
rect 17451 6820 18880 6848
rect 17451 6817 17463 6820
rect 17405 6811 17463 6817
rect 18874 6808 18880 6820
rect 18932 6808 18938 6860
rect 24946 6808 24952 6860
rect 25004 6848 25010 6860
rect 25958 6848 25964 6860
rect 25004 6820 25964 6848
rect 25004 6808 25010 6820
rect 25958 6808 25964 6820
rect 26016 6848 26022 6860
rect 28994 6848 29000 6860
rect 26016 6820 29000 6848
rect 26016 6808 26022 6820
rect 28994 6808 29000 6820
rect 29052 6848 29058 6860
rect 30392 6848 30420 6879
rect 29052 6820 29960 6848
rect 29052 6808 29058 6820
rect 29932 6792 29960 6820
rect 30024 6820 30420 6848
rect 15473 6783 15531 6789
rect 15473 6749 15485 6783
rect 15519 6749 15531 6783
rect 15473 6743 15531 6749
rect 15657 6783 15715 6789
rect 15657 6749 15669 6783
rect 15703 6749 15715 6783
rect 15657 6743 15715 6749
rect 20530 6740 20536 6792
rect 20588 6780 20594 6792
rect 20901 6783 20959 6789
rect 20901 6780 20913 6783
rect 20588 6752 20913 6780
rect 20588 6740 20594 6752
rect 20901 6749 20913 6752
rect 20947 6749 20959 6783
rect 20901 6743 20959 6749
rect 29270 6740 29276 6792
rect 29328 6780 29334 6792
rect 29549 6783 29607 6789
rect 29549 6780 29561 6783
rect 29328 6752 29561 6780
rect 29328 6740 29334 6752
rect 29549 6749 29561 6752
rect 29595 6749 29607 6783
rect 29549 6743 29607 6749
rect 29914 6740 29920 6792
rect 29972 6740 29978 6792
rect 11882 6672 11888 6724
rect 11940 6712 11946 6724
rect 12069 6715 12127 6721
rect 12069 6712 12081 6715
rect 11940 6684 12081 6712
rect 11940 6672 11946 6684
rect 12069 6681 12081 6684
rect 12115 6681 12127 6715
rect 12069 6675 12127 6681
rect 14185 6715 14243 6721
rect 14185 6681 14197 6715
rect 14231 6681 14243 6715
rect 14185 6675 14243 6681
rect 15766 6715 15824 6721
rect 15766 6681 15778 6715
rect 15812 6712 15824 6715
rect 15930 6712 15936 6724
rect 15812 6684 15936 6712
rect 15812 6681 15824 6684
rect 15766 6675 15824 6681
rect 12529 6647 12587 6653
rect 12529 6613 12541 6647
rect 12575 6644 12587 6647
rect 14200 6644 14228 6675
rect 15930 6672 15936 6684
rect 15988 6672 15994 6724
rect 18598 6672 18604 6724
rect 18656 6712 18662 6724
rect 21542 6712 21548 6724
rect 18656 6684 21548 6712
rect 18656 6672 18662 6684
rect 21542 6672 21548 6684
rect 21600 6672 21606 6724
rect 29454 6672 29460 6724
rect 29512 6712 29518 6724
rect 29733 6715 29791 6721
rect 29733 6712 29745 6715
rect 29512 6684 29745 6712
rect 29512 6672 29518 6684
rect 29733 6681 29745 6684
rect 29779 6681 29791 6715
rect 29733 6675 29791 6681
rect 29825 6715 29883 6721
rect 29825 6681 29837 6715
rect 29871 6712 29883 6715
rect 30024 6712 30052 6820
rect 33594 6808 33600 6860
rect 33652 6848 33658 6860
rect 33781 6851 33839 6857
rect 33781 6848 33793 6851
rect 33652 6820 33793 6848
rect 33652 6808 33658 6820
rect 33781 6817 33793 6820
rect 33827 6817 33839 6851
rect 33781 6811 33839 6817
rect 30190 6740 30196 6792
rect 30248 6740 30254 6792
rect 33686 6740 33692 6792
rect 33744 6780 33750 6792
rect 34256 6789 34284 6888
rect 37458 6848 37464 6860
rect 36648 6820 37464 6848
rect 34241 6783 34299 6789
rect 34241 6780 34253 6783
rect 33744 6752 34253 6780
rect 33744 6740 33750 6752
rect 34241 6749 34253 6752
rect 34287 6749 34299 6783
rect 34241 6743 34299 6749
rect 36648 6712 36676 6820
rect 37458 6808 37464 6820
rect 37516 6808 37522 6860
rect 38105 6851 38163 6857
rect 38105 6817 38117 6851
rect 38151 6848 38163 6851
rect 38194 6848 38200 6860
rect 38151 6820 38200 6848
rect 38151 6817 38163 6820
rect 38105 6811 38163 6817
rect 38194 6808 38200 6820
rect 38252 6808 38258 6860
rect 29871 6684 30052 6712
rect 30208 6698 36676 6712
rect 30208 6684 36662 6698
rect 29871 6681 29883 6684
rect 29825 6675 29883 6681
rect 12575 6616 14228 6644
rect 14645 6647 14703 6653
rect 12575 6613 12587 6616
rect 12529 6607 12587 6613
rect 14645 6613 14657 6647
rect 14691 6644 14703 6647
rect 15010 6644 15016 6656
rect 14691 6616 15016 6644
rect 14691 6613 14703 6616
rect 14645 6607 14703 6613
rect 15010 6604 15016 6616
rect 15068 6644 15074 6656
rect 16666 6644 16672 6656
rect 15068 6616 16672 6644
rect 15068 6604 15074 6616
rect 16666 6604 16672 6616
rect 16724 6604 16730 6656
rect 16758 6604 16764 6656
rect 16816 6604 16822 6656
rect 17126 6604 17132 6656
rect 17184 6644 17190 6656
rect 25314 6644 25320 6656
rect 17184 6616 25320 6644
rect 17184 6604 17190 6616
rect 25314 6604 25320 6616
rect 25372 6604 25378 6656
rect 28074 6604 28080 6656
rect 28132 6644 28138 6656
rect 29840 6644 29868 6675
rect 30208 6656 30236 6684
rect 28132 6616 29868 6644
rect 28132 6604 28138 6616
rect 30098 6604 30104 6656
rect 30156 6604 30162 6656
rect 30190 6604 30196 6656
rect 30248 6604 30254 6656
rect 1104 6554 40572 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 40572 6554
rect 1104 6480 40572 6502
rect 11882 6400 11888 6452
rect 11940 6400 11946 6452
rect 13630 6400 13636 6452
rect 13688 6440 13694 6452
rect 15102 6440 15108 6452
rect 13688 6412 15108 6440
rect 13688 6400 13694 6412
rect 15102 6400 15108 6412
rect 15160 6400 15166 6452
rect 16390 6400 16396 6452
rect 16448 6440 16454 6452
rect 17126 6440 17132 6452
rect 16448 6412 17132 6440
rect 16448 6400 16454 6412
rect 17126 6400 17132 6412
rect 17184 6400 17190 6452
rect 17865 6443 17923 6449
rect 17865 6409 17877 6443
rect 17911 6440 17923 6443
rect 19058 6440 19064 6452
rect 17911 6412 19064 6440
rect 17911 6409 17923 6412
rect 17865 6403 17923 6409
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 21266 6400 21272 6452
rect 21324 6440 21330 6452
rect 21453 6443 21511 6449
rect 21453 6440 21465 6443
rect 21324 6412 21465 6440
rect 21324 6400 21330 6412
rect 21453 6409 21465 6412
rect 21499 6409 21511 6443
rect 21453 6403 21511 6409
rect 24486 6400 24492 6452
rect 24544 6440 24550 6452
rect 26510 6440 26516 6452
rect 24544 6412 26516 6440
rect 24544 6400 24550 6412
rect 26510 6400 26516 6412
rect 26568 6440 26574 6452
rect 26605 6443 26663 6449
rect 26605 6440 26617 6443
rect 26568 6412 26617 6440
rect 26568 6400 26574 6412
rect 26605 6409 26617 6412
rect 26651 6409 26663 6443
rect 26605 6403 26663 6409
rect 26878 6400 26884 6452
rect 26936 6440 26942 6452
rect 29178 6440 29184 6452
rect 26936 6412 29184 6440
rect 26936 6400 26942 6412
rect 29178 6400 29184 6412
rect 29236 6400 29242 6452
rect 29457 6443 29515 6449
rect 29457 6409 29469 6443
rect 29503 6440 29515 6443
rect 29546 6440 29552 6452
rect 29503 6412 29552 6440
rect 29503 6409 29515 6412
rect 29457 6403 29515 6409
rect 29546 6400 29552 6412
rect 29604 6400 29610 6452
rect 30098 6400 30104 6452
rect 30156 6440 30162 6452
rect 30156 6412 30972 6440
rect 30156 6400 30162 6412
rect 15194 6372 15200 6384
rect 14660 6344 15200 6372
rect 14660 6313 14688 6344
rect 15194 6332 15200 6344
rect 15252 6332 15258 6384
rect 15378 6332 15384 6384
rect 15436 6332 15442 6384
rect 16850 6332 16856 6384
rect 16908 6372 16914 6384
rect 17678 6372 17684 6384
rect 16908 6344 17684 6372
rect 16908 6332 16914 6344
rect 17678 6332 17684 6344
rect 17736 6372 17742 6384
rect 17736 6344 18170 6372
rect 17736 6332 17742 6344
rect 19334 6332 19340 6384
rect 19392 6332 19398 6384
rect 20254 6332 20260 6384
rect 20312 6372 20318 6384
rect 20312 6344 20470 6372
rect 20312 6332 20318 6344
rect 22370 6332 22376 6384
rect 22428 6372 22434 6384
rect 26234 6372 26240 6384
rect 22428 6344 26240 6372
rect 22428 6332 22434 6344
rect 26234 6332 26240 6344
rect 26292 6332 26298 6384
rect 27617 6375 27675 6381
rect 27617 6372 27629 6375
rect 27264 6344 27629 6372
rect 11977 6307 12035 6313
rect 11977 6273 11989 6307
rect 12023 6304 12035 6307
rect 12345 6307 12403 6313
rect 12345 6304 12357 6307
rect 12023 6276 12357 6304
rect 12023 6273 12035 6276
rect 11977 6267 12035 6273
rect 12345 6273 12357 6276
rect 12391 6273 12403 6307
rect 12345 6267 12403 6273
rect 14645 6307 14703 6313
rect 14645 6273 14657 6307
rect 14691 6273 14703 6307
rect 14645 6267 14703 6273
rect 24946 6264 24952 6316
rect 25004 6264 25010 6316
rect 25406 6304 25412 6316
rect 25056 6276 25412 6304
rect 12161 6239 12219 6245
rect 12161 6205 12173 6239
rect 12207 6205 12219 6239
rect 12161 6199 12219 6205
rect 12176 6168 12204 6199
rect 12250 6196 12256 6248
rect 12308 6236 12314 6248
rect 12897 6239 12955 6245
rect 12897 6236 12909 6239
rect 12308 6208 12909 6236
rect 12308 6196 12314 6208
rect 12897 6205 12909 6208
rect 12943 6205 12955 6239
rect 12897 6199 12955 6205
rect 14921 6239 14979 6245
rect 14921 6205 14933 6239
rect 14967 6236 14979 6239
rect 16758 6236 16764 6248
rect 14967 6208 16764 6236
rect 14967 6205 14979 6208
rect 14921 6199 14979 6205
rect 16758 6196 16764 6208
rect 16816 6196 16822 6248
rect 17218 6196 17224 6248
rect 17276 6236 17282 6248
rect 19613 6239 19671 6245
rect 19613 6236 19625 6239
rect 17276 6208 19625 6236
rect 17276 6196 17282 6208
rect 19613 6205 19625 6208
rect 19659 6236 19671 6239
rect 19705 6239 19763 6245
rect 19705 6236 19717 6239
rect 19659 6208 19717 6236
rect 19659 6205 19671 6208
rect 19613 6199 19671 6205
rect 19705 6205 19717 6208
rect 19751 6205 19763 6239
rect 19705 6199 19763 6205
rect 19981 6239 20039 6245
rect 19981 6205 19993 6239
rect 20027 6236 20039 6239
rect 20438 6236 20444 6248
rect 20027 6208 20444 6236
rect 20027 6205 20039 6208
rect 19981 6199 20039 6205
rect 20438 6196 20444 6208
rect 20496 6196 20502 6248
rect 22833 6239 22891 6245
rect 22833 6205 22845 6239
rect 22879 6236 22891 6239
rect 23014 6236 23020 6248
rect 22879 6208 23020 6236
rect 22879 6205 22891 6208
rect 22833 6199 22891 6205
rect 23014 6196 23020 6208
rect 23072 6196 23078 6248
rect 23750 6196 23756 6248
rect 23808 6236 23814 6248
rect 25056 6236 25084 6276
rect 25406 6264 25412 6276
rect 25464 6264 25470 6316
rect 26786 6264 26792 6316
rect 26844 6264 26850 6316
rect 26878 6264 26884 6316
rect 26936 6304 26942 6316
rect 27264 6313 27292 6344
rect 27617 6341 27629 6344
rect 27663 6341 27675 6375
rect 29362 6372 29368 6384
rect 27617 6335 27675 6341
rect 27908 6344 29368 6372
rect 27157 6307 27215 6313
rect 27157 6304 27169 6307
rect 26936 6276 27169 6304
rect 26936 6264 26942 6276
rect 27157 6273 27169 6276
rect 27203 6273 27215 6307
rect 27157 6267 27215 6273
rect 27249 6307 27307 6313
rect 27249 6273 27261 6307
rect 27295 6273 27307 6307
rect 27249 6267 27307 6273
rect 23808 6208 25084 6236
rect 23808 6196 23814 6208
rect 26234 6196 26240 6248
rect 26292 6236 26298 6248
rect 27264 6236 27292 6267
rect 27338 6264 27344 6316
rect 27396 6264 27402 6316
rect 27525 6307 27583 6313
rect 27525 6304 27537 6307
rect 27448 6276 27537 6304
rect 26292 6208 27292 6236
rect 26292 6196 26298 6208
rect 12986 6168 12992 6180
rect 12176 6140 12992 6168
rect 12986 6128 12992 6140
rect 13044 6128 13050 6180
rect 15930 6128 15936 6180
rect 15988 6168 15994 6180
rect 17236 6168 17264 6196
rect 15988 6140 17264 6168
rect 15988 6128 15994 6140
rect 22278 6128 22284 6180
rect 22336 6168 22342 6180
rect 22465 6171 22523 6177
rect 22465 6168 22477 6171
rect 22336 6140 22477 6168
rect 22336 6128 22342 6140
rect 22465 6137 22477 6140
rect 22511 6137 22523 6171
rect 22465 6131 22523 6137
rect 25590 6128 25596 6180
rect 25648 6168 25654 6180
rect 27448 6168 27476 6276
rect 27525 6273 27537 6276
rect 27571 6304 27583 6307
rect 27908 6304 27936 6344
rect 29362 6332 29368 6344
rect 29420 6332 29426 6384
rect 30190 6332 30196 6384
rect 30248 6332 30254 6384
rect 30944 6381 30972 6412
rect 30929 6375 30987 6381
rect 30929 6341 30941 6375
rect 30975 6341 30987 6375
rect 30929 6335 30987 6341
rect 27571 6276 27936 6304
rect 27985 6307 28043 6313
rect 27571 6273 27583 6276
rect 27525 6267 27583 6273
rect 27985 6273 27997 6307
rect 28031 6304 28043 6307
rect 28718 6304 28724 6316
rect 28031 6276 28724 6304
rect 28031 6273 28043 6276
rect 27985 6267 28043 6273
rect 28718 6264 28724 6276
rect 28776 6264 28782 6316
rect 31205 6307 31263 6313
rect 31205 6273 31217 6307
rect 31251 6304 31263 6307
rect 31294 6304 31300 6316
rect 31251 6276 31300 6304
rect 31251 6273 31263 6276
rect 31205 6267 31263 6273
rect 31294 6264 31300 6276
rect 31352 6304 31358 6316
rect 31662 6304 31668 6316
rect 31352 6276 31668 6304
rect 31352 6264 31358 6276
rect 31662 6264 31668 6276
rect 31720 6264 31726 6316
rect 25648 6140 27476 6168
rect 25648 6128 25654 6140
rect 10686 6060 10692 6112
rect 10744 6100 10750 6112
rect 11517 6103 11575 6109
rect 11517 6100 11529 6103
rect 10744 6072 11529 6100
rect 10744 6060 10750 6072
rect 11517 6069 11529 6072
rect 11563 6069 11575 6103
rect 11517 6063 11575 6069
rect 16206 6060 16212 6112
rect 16264 6100 16270 6112
rect 17954 6100 17960 6112
rect 16264 6072 17960 6100
rect 16264 6060 16270 6072
rect 17954 6060 17960 6072
rect 18012 6060 18018 6112
rect 19518 6060 19524 6112
rect 19576 6100 19582 6112
rect 21266 6100 21272 6112
rect 19576 6072 21272 6100
rect 19576 6060 19582 6072
rect 21266 6060 21272 6072
rect 21324 6060 21330 6112
rect 22186 6060 22192 6112
rect 22244 6100 22250 6112
rect 22370 6100 22376 6112
rect 22244 6072 22376 6100
rect 22244 6060 22250 6072
rect 22370 6060 22376 6072
rect 22428 6060 22434 6112
rect 23566 6060 23572 6112
rect 23624 6100 23630 6112
rect 24762 6100 24768 6112
rect 23624 6072 24768 6100
rect 23624 6060 23630 6072
rect 24762 6060 24768 6072
rect 24820 6060 24826 6112
rect 25130 6060 25136 6112
rect 25188 6060 25194 6112
rect 26973 6103 27031 6109
rect 26973 6069 26985 6103
rect 27019 6100 27031 6103
rect 27246 6100 27252 6112
rect 27019 6072 27252 6100
rect 27019 6069 27031 6072
rect 26973 6063 27031 6069
rect 27246 6060 27252 6072
rect 27304 6060 27310 6112
rect 27338 6060 27344 6112
rect 27396 6100 27402 6112
rect 29454 6100 29460 6112
rect 27396 6072 29460 6100
rect 27396 6060 27402 6072
rect 29454 6060 29460 6072
rect 29512 6060 29518 6112
rect 1104 6010 40572 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 40572 6010
rect 1104 5936 40572 5958
rect 18782 5856 18788 5908
rect 18840 5896 18846 5908
rect 18840 5868 19472 5896
rect 18840 5856 18846 5868
rect 19061 5831 19119 5837
rect 19061 5797 19073 5831
rect 19107 5828 19119 5831
rect 19334 5828 19340 5840
rect 19107 5800 19340 5828
rect 19107 5797 19119 5800
rect 19061 5791 19119 5797
rect 19334 5788 19340 5800
rect 19392 5788 19398 5840
rect 19444 5828 19472 5868
rect 19978 5856 19984 5908
rect 20036 5856 20042 5908
rect 20438 5856 20444 5908
rect 20496 5856 20502 5908
rect 21542 5856 21548 5908
rect 21600 5896 21606 5908
rect 25498 5896 25504 5908
rect 21600 5868 24808 5896
rect 21600 5856 21606 5868
rect 20714 5828 20720 5840
rect 19444 5800 20720 5828
rect 10413 5763 10471 5769
rect 10413 5729 10425 5763
rect 10459 5760 10471 5763
rect 10778 5760 10784 5772
rect 10459 5732 10784 5760
rect 10459 5729 10471 5732
rect 10413 5723 10471 5729
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 17681 5763 17739 5769
rect 17681 5729 17693 5763
rect 17727 5760 17739 5763
rect 18598 5760 18604 5772
rect 17727 5732 18604 5760
rect 17727 5729 17739 5732
rect 17681 5723 17739 5729
rect 18598 5720 18604 5732
rect 18656 5720 18662 5772
rect 18690 5720 18696 5772
rect 18748 5760 18754 5772
rect 19705 5763 19763 5769
rect 19705 5760 19717 5763
rect 18748 5732 19717 5760
rect 18748 5720 18754 5732
rect 19705 5729 19717 5732
rect 19751 5729 19763 5763
rect 19705 5723 19763 5729
rect 18506 5652 18512 5704
rect 18564 5652 18570 5704
rect 18782 5652 18788 5704
rect 18840 5652 18846 5704
rect 19150 5652 19156 5704
rect 19208 5692 19214 5704
rect 19337 5695 19395 5701
rect 19337 5692 19349 5695
rect 19208 5664 19349 5692
rect 19208 5652 19214 5664
rect 19337 5661 19349 5664
rect 19383 5661 19395 5695
rect 19337 5655 19395 5661
rect 19426 5652 19432 5704
rect 19484 5652 19490 5704
rect 19518 5652 19524 5704
rect 19576 5652 19582 5704
rect 19613 5695 19671 5701
rect 19613 5661 19625 5695
rect 19659 5661 19671 5695
rect 19613 5655 19671 5661
rect 19797 5695 19855 5701
rect 19797 5661 19809 5695
rect 19843 5692 19855 5695
rect 19886 5692 19892 5704
rect 19843 5664 19892 5692
rect 19843 5661 19855 5664
rect 19797 5655 19855 5661
rect 10686 5584 10692 5636
rect 10744 5584 10750 5636
rect 17405 5627 17463 5633
rect 10796 5596 11178 5624
rect 10594 5516 10600 5568
rect 10652 5556 10658 5568
rect 10796 5556 10824 5596
rect 17405 5593 17417 5627
rect 17451 5624 17463 5627
rect 18138 5624 18144 5636
rect 17451 5596 18144 5624
rect 17451 5593 17463 5596
rect 17405 5587 17463 5593
rect 18138 5584 18144 5596
rect 18196 5584 18202 5636
rect 19061 5627 19119 5633
rect 19061 5593 19073 5627
rect 19107 5624 19119 5627
rect 19444 5624 19472 5652
rect 19107 5596 19472 5624
rect 19107 5593 19119 5596
rect 19061 5587 19119 5593
rect 10652 5528 10824 5556
rect 10652 5516 10658 5528
rect 11330 5516 11336 5568
rect 11388 5556 11394 5568
rect 12161 5559 12219 5565
rect 12161 5556 12173 5559
rect 11388 5528 12173 5556
rect 11388 5516 11394 5528
rect 12161 5525 12173 5528
rect 12207 5556 12219 5559
rect 12250 5556 12256 5568
rect 12207 5528 12256 5556
rect 12207 5525 12219 5528
rect 12161 5519 12219 5525
rect 12250 5516 12256 5528
rect 12308 5516 12314 5568
rect 17034 5516 17040 5568
rect 17092 5516 17098 5568
rect 17497 5559 17555 5565
rect 17497 5525 17509 5559
rect 17543 5556 17555 5559
rect 17957 5559 18015 5565
rect 17957 5556 17969 5559
rect 17543 5528 17969 5556
rect 17543 5525 17555 5528
rect 17497 5519 17555 5525
rect 17957 5525 17969 5528
rect 18003 5525 18015 5559
rect 17957 5519 18015 5525
rect 18877 5559 18935 5565
rect 18877 5525 18889 5559
rect 18923 5556 18935 5559
rect 19242 5556 19248 5568
rect 18923 5528 19248 5556
rect 18923 5525 18935 5528
rect 18877 5519 18935 5525
rect 19242 5516 19248 5528
rect 19300 5516 19306 5568
rect 19429 5559 19487 5565
rect 19429 5525 19441 5559
rect 19475 5556 19487 5559
rect 19628 5556 19656 5655
rect 19886 5652 19892 5664
rect 19944 5692 19950 5704
rect 19944 5664 20024 5692
rect 19944 5652 19950 5664
rect 19996 5624 20024 5664
rect 20070 5652 20076 5704
rect 20128 5652 20134 5704
rect 20257 5695 20315 5701
rect 20257 5661 20269 5695
rect 20303 5692 20315 5695
rect 20364 5692 20392 5800
rect 20714 5788 20720 5800
rect 20772 5788 20778 5840
rect 21358 5788 21364 5840
rect 21416 5788 21422 5840
rect 20901 5763 20959 5769
rect 20901 5760 20913 5763
rect 20456 5732 20913 5760
rect 20456 5701 20484 5732
rect 20901 5729 20913 5732
rect 20947 5729 20959 5763
rect 21376 5760 21404 5788
rect 22189 5763 22247 5769
rect 21376 5732 21864 5760
rect 20901 5723 20959 5729
rect 20303 5664 20392 5692
rect 20441 5695 20499 5701
rect 20303 5661 20315 5664
rect 20257 5655 20315 5661
rect 20441 5661 20453 5695
rect 20487 5661 20499 5695
rect 20441 5655 20499 5661
rect 20530 5652 20536 5704
rect 20588 5652 20594 5704
rect 21085 5695 21143 5701
rect 21085 5661 21097 5695
rect 21131 5692 21143 5695
rect 21266 5692 21272 5704
rect 21131 5664 21272 5692
rect 21131 5661 21143 5664
rect 21085 5655 21143 5661
rect 21266 5652 21272 5664
rect 21324 5652 21330 5704
rect 21361 5695 21419 5701
rect 21361 5661 21373 5695
rect 21407 5661 21419 5695
rect 21361 5655 21419 5661
rect 20625 5627 20683 5633
rect 20625 5624 20637 5627
rect 19996 5596 20637 5624
rect 20625 5593 20637 5596
rect 20671 5593 20683 5627
rect 21376 5624 21404 5655
rect 21542 5652 21548 5704
rect 21600 5652 21606 5704
rect 21637 5695 21695 5701
rect 21637 5661 21649 5695
rect 21683 5692 21695 5695
rect 21726 5692 21732 5704
rect 21683 5664 21732 5692
rect 21683 5661 21695 5664
rect 21637 5655 21695 5661
rect 21726 5652 21732 5664
rect 21784 5652 21790 5704
rect 21836 5701 21864 5732
rect 22189 5729 22201 5763
rect 22235 5760 22247 5763
rect 23198 5760 23204 5772
rect 22235 5732 23204 5760
rect 22235 5729 22247 5732
rect 22189 5723 22247 5729
rect 23198 5720 23204 5732
rect 23256 5720 23262 5772
rect 24210 5720 24216 5772
rect 24268 5720 24274 5772
rect 21821 5695 21879 5701
rect 21821 5661 21833 5695
rect 21867 5692 21879 5695
rect 22094 5692 22100 5704
rect 21867 5664 22100 5692
rect 21867 5661 21879 5664
rect 21821 5655 21879 5661
rect 22094 5652 22100 5664
rect 22152 5652 22158 5704
rect 24486 5652 24492 5704
rect 24544 5652 24550 5704
rect 24780 5692 24808 5868
rect 25240 5868 25504 5896
rect 24854 5788 24860 5840
rect 24912 5788 24918 5840
rect 24946 5788 24952 5840
rect 25004 5828 25010 5840
rect 25240 5828 25268 5868
rect 25498 5856 25504 5868
rect 25556 5896 25562 5908
rect 26418 5896 26424 5908
rect 25556 5868 26424 5896
rect 25556 5856 25562 5868
rect 26418 5856 26424 5868
rect 26476 5856 26482 5908
rect 26712 5868 28580 5896
rect 26712 5840 26740 5868
rect 25004 5800 25268 5828
rect 25004 5788 25010 5800
rect 25406 5788 25412 5840
rect 25464 5828 25470 5840
rect 26694 5828 26700 5840
rect 25464 5800 26700 5828
rect 25464 5788 25470 5800
rect 26694 5788 26700 5800
rect 26752 5788 26758 5840
rect 24872 5760 24900 5788
rect 26973 5763 27031 5769
rect 26973 5760 26985 5763
rect 24872 5732 26985 5760
rect 26973 5729 26985 5732
rect 27019 5729 27031 5763
rect 26973 5723 27031 5729
rect 27246 5720 27252 5772
rect 27304 5720 27310 5772
rect 24857 5695 24915 5701
rect 24857 5692 24869 5695
rect 24780 5664 24869 5692
rect 24857 5661 24869 5664
rect 24903 5692 24915 5695
rect 25130 5692 25136 5704
rect 24903 5664 25136 5692
rect 24903 5661 24915 5664
rect 24857 5655 24915 5661
rect 25130 5652 25136 5664
rect 25188 5692 25194 5704
rect 25317 5695 25375 5701
rect 25317 5692 25329 5695
rect 25188 5664 25329 5692
rect 25188 5652 25194 5664
rect 25317 5661 25329 5664
rect 25363 5692 25375 5695
rect 25363 5664 25636 5692
rect 25363 5661 25375 5664
rect 25317 5655 25375 5661
rect 22186 5624 22192 5636
rect 21376 5596 22192 5624
rect 20625 5587 20683 5593
rect 22186 5584 22192 5596
rect 22244 5584 22250 5636
rect 22462 5584 22468 5636
rect 22520 5584 22526 5636
rect 24578 5624 24584 5636
rect 23690 5596 24584 5624
rect 24578 5584 24584 5596
rect 24636 5584 24642 5636
rect 24673 5627 24731 5633
rect 24673 5593 24685 5627
rect 24719 5593 24731 5627
rect 24673 5587 24731 5593
rect 21726 5556 21732 5568
rect 19475 5528 21732 5556
rect 19475 5525 19487 5528
rect 19429 5519 19487 5525
rect 21726 5516 21732 5528
rect 21784 5516 21790 5568
rect 21821 5559 21879 5565
rect 21821 5525 21833 5559
rect 21867 5556 21879 5559
rect 22370 5556 22376 5568
rect 21867 5528 22376 5556
rect 21867 5525 21879 5528
rect 21821 5519 21879 5525
rect 22370 5516 22376 5528
rect 22428 5516 22434 5568
rect 24688 5556 24716 5587
rect 24762 5584 24768 5636
rect 24820 5624 24826 5636
rect 24820 5596 25360 5624
rect 24820 5584 24826 5596
rect 24946 5556 24952 5568
rect 24688 5528 24952 5556
rect 24946 5516 24952 5528
rect 25004 5516 25010 5568
rect 25038 5516 25044 5568
rect 25096 5516 25102 5568
rect 25130 5516 25136 5568
rect 25188 5516 25194 5568
rect 25332 5556 25360 5596
rect 25406 5584 25412 5636
rect 25464 5584 25470 5636
rect 25498 5584 25504 5636
rect 25556 5584 25562 5636
rect 25608 5624 25636 5664
rect 25682 5652 25688 5704
rect 25740 5652 25746 5704
rect 25774 5652 25780 5704
rect 25832 5652 25838 5704
rect 26234 5652 26240 5704
rect 26292 5652 26298 5704
rect 26605 5695 26663 5701
rect 26605 5692 26617 5695
rect 26344 5664 26617 5692
rect 26344 5624 26372 5664
rect 26605 5661 26617 5664
rect 26651 5692 26663 5695
rect 26878 5692 26884 5704
rect 26651 5664 26884 5692
rect 26651 5661 26663 5664
rect 26605 5655 26663 5661
rect 26878 5652 26884 5664
rect 26936 5652 26942 5704
rect 28552 5692 28580 5868
rect 28718 5856 28724 5908
rect 28776 5856 28782 5908
rect 29546 5896 29552 5908
rect 29104 5868 29552 5896
rect 29104 5701 29132 5868
rect 29546 5856 29552 5868
rect 29604 5856 29610 5908
rect 29365 5831 29423 5837
rect 29365 5797 29377 5831
rect 29411 5797 29423 5831
rect 29365 5791 29423 5797
rect 29380 5760 29408 5791
rect 31021 5763 31079 5769
rect 31021 5760 31033 5763
rect 29380 5732 31033 5760
rect 31021 5729 31033 5732
rect 31067 5729 31079 5763
rect 31021 5723 31079 5729
rect 31294 5720 31300 5772
rect 31352 5720 31358 5772
rect 28813 5695 28871 5701
rect 28813 5692 28825 5695
rect 28552 5664 28825 5692
rect 28813 5661 28825 5664
rect 28859 5661 28871 5695
rect 28813 5655 28871 5661
rect 29089 5695 29147 5701
rect 29089 5661 29101 5695
rect 29135 5661 29147 5695
rect 29089 5655 29147 5661
rect 29178 5652 29184 5704
rect 29236 5652 29242 5704
rect 25608 5596 26372 5624
rect 26418 5584 26424 5636
rect 26476 5584 26482 5636
rect 26510 5584 26516 5636
rect 26568 5584 26574 5636
rect 27338 5624 27344 5636
rect 26620 5596 27344 5624
rect 25682 5556 25688 5568
rect 25332 5528 25688 5556
rect 25682 5516 25688 5528
rect 25740 5516 25746 5568
rect 25958 5516 25964 5568
rect 26016 5516 26022 5568
rect 26436 5556 26464 5584
rect 26620 5556 26648 5596
rect 27338 5584 27344 5596
rect 27396 5584 27402 5636
rect 28997 5627 29055 5633
rect 28474 5596 28580 5624
rect 26436 5528 26648 5556
rect 26789 5559 26847 5565
rect 26789 5525 26801 5559
rect 26835 5556 26847 5559
rect 28074 5556 28080 5568
rect 26835 5528 28080 5556
rect 26835 5525 26847 5528
rect 26789 5519 26847 5525
rect 28074 5516 28080 5528
rect 28132 5516 28138 5568
rect 28552 5556 28580 5596
rect 28997 5593 29009 5627
rect 29043 5624 29055 5627
rect 29454 5624 29460 5636
rect 29043 5596 29460 5624
rect 29043 5593 29055 5596
rect 28997 5587 29055 5593
rect 29454 5584 29460 5596
rect 29512 5584 29518 5636
rect 30282 5584 30288 5636
rect 30340 5584 30346 5636
rect 29086 5556 29092 5568
rect 28552 5528 29092 5556
rect 29086 5516 29092 5528
rect 29144 5516 29150 5568
rect 1104 5466 40572 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 40572 5466
rect 1104 5392 40572 5414
rect 13541 5355 13599 5361
rect 13541 5321 13553 5355
rect 13587 5352 13599 5355
rect 13814 5352 13820 5364
rect 13587 5324 13820 5352
rect 13587 5321 13599 5324
rect 13541 5315 13599 5321
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 18417 5355 18475 5361
rect 14292 5324 15240 5352
rect 13354 5284 13360 5296
rect 13294 5256 13360 5284
rect 13354 5244 13360 5256
rect 13412 5284 13418 5296
rect 14292 5284 14320 5324
rect 15212 5284 15240 5324
rect 18417 5321 18429 5355
rect 18463 5352 18475 5355
rect 18506 5352 18512 5364
rect 18463 5324 18512 5352
rect 18463 5321 18475 5324
rect 18417 5315 18475 5321
rect 18506 5312 18512 5324
rect 18564 5312 18570 5364
rect 21358 5312 21364 5364
rect 21416 5352 21422 5364
rect 22278 5352 22284 5364
rect 21416 5324 22284 5352
rect 21416 5312 21422 5324
rect 22278 5312 22284 5324
rect 22336 5312 22342 5364
rect 22462 5312 22468 5364
rect 22520 5352 22526 5364
rect 22557 5355 22615 5361
rect 22557 5352 22569 5355
rect 22520 5324 22569 5352
rect 22520 5312 22526 5324
rect 22557 5321 22569 5324
rect 22603 5321 22615 5355
rect 22557 5315 22615 5321
rect 23569 5355 23627 5361
rect 23569 5321 23581 5355
rect 23615 5352 23627 5355
rect 25774 5352 25780 5364
rect 23615 5324 25780 5352
rect 23615 5321 23627 5324
rect 23569 5315 23627 5321
rect 25774 5312 25780 5324
rect 25832 5312 25838 5364
rect 26786 5312 26792 5364
rect 26844 5352 26850 5364
rect 26973 5355 27031 5361
rect 26973 5352 26985 5355
rect 26844 5324 26985 5352
rect 26844 5312 26850 5324
rect 26973 5321 26985 5324
rect 27019 5321 27031 5355
rect 29086 5352 29092 5364
rect 26973 5315 27031 5321
rect 27080 5324 29092 5352
rect 15378 5284 15384 5296
rect 13412 5256 14320 5284
rect 15134 5256 15384 5284
rect 13412 5244 13418 5256
rect 15378 5244 15384 5256
rect 15436 5244 15442 5296
rect 16945 5287 17003 5293
rect 16945 5253 16957 5287
rect 16991 5284 17003 5287
rect 17034 5284 17040 5296
rect 16991 5256 17040 5284
rect 16991 5253 17003 5256
rect 16945 5247 17003 5253
rect 17034 5244 17040 5256
rect 17092 5244 17098 5296
rect 17678 5244 17684 5296
rect 17736 5244 17742 5296
rect 10962 5176 10968 5228
rect 11020 5216 11026 5228
rect 18524 5225 18552 5312
rect 20070 5244 20076 5296
rect 20128 5284 20134 5296
rect 20128 5256 21312 5284
rect 20128 5244 20134 5256
rect 11793 5219 11851 5225
rect 11793 5216 11805 5219
rect 11020 5188 11805 5216
rect 11020 5176 11026 5188
rect 11793 5185 11805 5188
rect 11839 5185 11851 5219
rect 11793 5179 11851 5185
rect 18509 5219 18567 5225
rect 18509 5185 18521 5219
rect 18555 5185 18567 5219
rect 18509 5179 18567 5185
rect 18598 5176 18604 5228
rect 18656 5216 18662 5228
rect 18785 5219 18843 5225
rect 18785 5216 18797 5219
rect 18656 5188 18797 5216
rect 18656 5176 18662 5188
rect 18785 5185 18797 5188
rect 18831 5185 18843 5219
rect 18785 5179 18843 5185
rect 19334 5176 19340 5228
rect 19392 5176 19398 5228
rect 20349 5219 20407 5225
rect 20349 5185 20361 5219
rect 20395 5216 20407 5219
rect 20622 5216 20628 5228
rect 20395 5188 20628 5216
rect 20395 5185 20407 5188
rect 20349 5179 20407 5185
rect 20622 5176 20628 5188
rect 20680 5176 20686 5228
rect 21284 5225 21312 5256
rect 22370 5244 22376 5296
rect 22428 5284 22434 5296
rect 22925 5287 22983 5293
rect 22925 5284 22937 5287
rect 22428 5256 22937 5284
rect 22428 5244 22434 5256
rect 22925 5253 22937 5256
rect 22971 5253 22983 5287
rect 24210 5284 24216 5296
rect 22925 5247 22983 5253
rect 23124 5256 24216 5284
rect 20717 5219 20775 5225
rect 20717 5185 20729 5219
rect 20763 5185 20775 5219
rect 20717 5179 20775 5185
rect 21269 5219 21327 5225
rect 21269 5185 21281 5219
rect 21315 5185 21327 5219
rect 21269 5179 21327 5185
rect 12066 5108 12072 5160
rect 12124 5108 12130 5160
rect 13633 5151 13691 5157
rect 13633 5117 13645 5151
rect 13679 5117 13691 5151
rect 13633 5111 13691 5117
rect 13909 5151 13967 5157
rect 13909 5117 13921 5151
rect 13955 5148 13967 5151
rect 14274 5148 14280 5160
rect 13955 5120 14280 5148
rect 13955 5117 13967 5120
rect 13909 5111 13967 5117
rect 13648 5012 13676 5111
rect 14274 5108 14280 5120
rect 14332 5108 14338 5160
rect 16025 5151 16083 5157
rect 16025 5148 16037 5151
rect 15580 5120 16037 5148
rect 14918 5040 14924 5092
rect 14976 5080 14982 5092
rect 15473 5083 15531 5089
rect 15473 5080 15485 5083
rect 14976 5052 15485 5080
rect 14976 5040 14982 5052
rect 15473 5049 15485 5052
rect 15519 5049 15531 5083
rect 15473 5043 15531 5049
rect 15194 5012 15200 5024
rect 13648 4984 15200 5012
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 15378 4972 15384 5024
rect 15436 5012 15442 5024
rect 15580 5012 15608 5120
rect 16025 5117 16037 5120
rect 16071 5117 16083 5151
rect 16025 5111 16083 5117
rect 16669 5151 16727 5157
rect 16669 5117 16681 5151
rect 16715 5148 16727 5151
rect 17034 5148 17040 5160
rect 16715 5120 17040 5148
rect 16715 5117 16727 5120
rect 16669 5111 16727 5117
rect 17034 5108 17040 5120
rect 17092 5108 17098 5160
rect 17494 5108 17500 5160
rect 17552 5148 17558 5160
rect 17552 5120 18000 5148
rect 17552 5108 17558 5120
rect 17972 5080 18000 5120
rect 18966 5108 18972 5160
rect 19024 5148 19030 5160
rect 19024 5120 20208 5148
rect 19024 5108 19030 5120
rect 19061 5083 19119 5089
rect 19061 5080 19073 5083
rect 17972 5052 19073 5080
rect 19061 5049 19073 5052
rect 19107 5049 19119 5083
rect 19061 5043 19119 5049
rect 19334 5040 19340 5092
rect 19392 5080 19398 5092
rect 20070 5080 20076 5092
rect 19392 5052 20076 5080
rect 19392 5040 19398 5052
rect 20070 5040 20076 5052
rect 20128 5040 20134 5092
rect 20180 5080 20208 5120
rect 20533 5083 20591 5089
rect 20533 5080 20545 5083
rect 20180 5052 20545 5080
rect 20533 5049 20545 5052
rect 20579 5080 20591 5083
rect 20732 5080 20760 5179
rect 21450 5176 21456 5228
rect 21508 5176 21514 5228
rect 22094 5176 22100 5228
rect 22152 5216 22158 5228
rect 22741 5219 22799 5225
rect 22741 5216 22753 5219
rect 22152 5188 22753 5216
rect 22152 5176 22158 5188
rect 22741 5185 22753 5188
rect 22787 5185 22799 5219
rect 22741 5179 22799 5185
rect 22833 5219 22891 5225
rect 22833 5185 22845 5219
rect 22879 5216 22891 5219
rect 23014 5216 23020 5228
rect 22879 5188 23020 5216
rect 22879 5185 22891 5188
rect 22833 5179 22891 5185
rect 23014 5176 23020 5188
rect 23072 5176 23078 5228
rect 23124 5225 23152 5256
rect 24210 5244 24216 5256
rect 24268 5244 24274 5296
rect 24854 5284 24860 5296
rect 24688 5256 24860 5284
rect 23109 5219 23167 5225
rect 23109 5185 23121 5219
rect 23155 5185 23167 5219
rect 23109 5179 23167 5185
rect 23201 5219 23259 5225
rect 23201 5185 23213 5219
rect 23247 5185 23259 5219
rect 23201 5179 23259 5185
rect 23385 5219 23443 5225
rect 23385 5185 23397 5219
rect 23431 5216 23443 5219
rect 23934 5216 23940 5228
rect 23431 5188 23940 5216
rect 23431 5185 23443 5188
rect 23385 5179 23443 5185
rect 22370 5108 22376 5160
rect 22428 5108 22434 5160
rect 20579 5052 20760 5080
rect 20579 5049 20591 5052
rect 20533 5043 20591 5049
rect 22830 5040 22836 5092
rect 22888 5080 22894 5092
rect 23216 5080 23244 5179
rect 23934 5176 23940 5188
rect 23992 5176 23998 5228
rect 24688 5225 24716 5256
rect 24854 5244 24860 5256
rect 24912 5244 24918 5296
rect 24949 5287 25007 5293
rect 24949 5253 24961 5287
rect 24995 5284 25007 5287
rect 25038 5284 25044 5296
rect 24995 5256 25044 5284
rect 24995 5253 25007 5256
rect 24949 5247 25007 5253
rect 25038 5244 25044 5256
rect 25096 5244 25102 5296
rect 27080 5284 27108 5324
rect 28092 5284 28120 5324
rect 29086 5312 29092 5324
rect 29144 5352 29150 5364
rect 30282 5352 30288 5364
rect 29144 5324 30288 5352
rect 29144 5312 29150 5324
rect 30282 5312 30288 5324
rect 30340 5312 30346 5364
rect 26174 5270 27108 5284
rect 26160 5256 27108 5270
rect 28014 5256 28120 5284
rect 24673 5219 24731 5225
rect 24673 5185 24685 5219
rect 24719 5185 24731 5219
rect 24673 5179 24731 5185
rect 26160 5160 26188 5256
rect 28166 5244 28172 5296
rect 28224 5284 28230 5296
rect 31294 5284 31300 5296
rect 28224 5256 31300 5284
rect 28224 5244 28230 5256
rect 28736 5225 28764 5256
rect 31294 5244 31300 5256
rect 31352 5244 31358 5296
rect 28721 5219 28779 5225
rect 28721 5185 28733 5219
rect 28767 5185 28779 5219
rect 28721 5179 28779 5185
rect 28994 5176 29000 5228
rect 29052 5176 29058 5228
rect 29178 5176 29184 5228
rect 29236 5176 29242 5228
rect 30190 5176 30196 5228
rect 30248 5176 30254 5228
rect 25682 5108 25688 5160
rect 25740 5148 25746 5160
rect 25740 5120 26096 5148
rect 25740 5108 25746 5120
rect 22888 5052 23244 5080
rect 26068 5080 26096 5120
rect 26142 5108 26148 5160
rect 26200 5108 26206 5160
rect 26697 5151 26755 5157
rect 26697 5117 26709 5151
rect 26743 5117 26755 5151
rect 26697 5111 26755 5117
rect 26712 5080 26740 5111
rect 28074 5108 28080 5160
rect 28132 5148 28138 5160
rect 28445 5151 28503 5157
rect 28445 5148 28457 5151
rect 28132 5120 28457 5148
rect 28132 5108 28138 5120
rect 28445 5117 28457 5120
rect 28491 5117 28503 5151
rect 28445 5111 28503 5117
rect 26068 5052 26740 5080
rect 22888 5040 22894 5052
rect 15436 4984 15608 5012
rect 15436 4972 15442 4984
rect 18138 4972 18144 5024
rect 18196 5012 18202 5024
rect 18601 5015 18659 5021
rect 18601 5012 18613 5015
rect 18196 4984 18613 5012
rect 18196 4972 18202 4984
rect 18601 4981 18613 4984
rect 18647 4981 18659 5015
rect 18601 4975 18659 4981
rect 19518 4972 19524 5024
rect 19576 5012 19582 5024
rect 19981 5015 20039 5021
rect 19981 5012 19993 5015
rect 19576 4984 19993 5012
rect 19576 4972 19582 4984
rect 19981 4981 19993 4984
rect 20027 4981 20039 5015
rect 19981 4975 20039 4981
rect 20257 5015 20315 5021
rect 20257 4981 20269 5015
rect 20303 5012 20315 5015
rect 20622 5012 20628 5024
rect 20303 4984 20628 5012
rect 20303 4981 20315 4984
rect 20257 4975 20315 4981
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 20898 4972 20904 5024
rect 20956 4972 20962 5024
rect 21266 4972 21272 5024
rect 21324 5012 21330 5024
rect 21821 5015 21879 5021
rect 21821 5012 21833 5015
rect 21324 4984 21833 5012
rect 21324 4972 21330 4984
rect 21821 4981 21833 4984
rect 21867 4981 21879 5015
rect 21821 4975 21879 4981
rect 28626 4972 28632 5024
rect 28684 5012 28690 5024
rect 28813 5015 28871 5021
rect 28813 5012 28825 5015
rect 28684 4984 28825 5012
rect 28684 4972 28690 4984
rect 28813 4981 28825 4984
rect 28859 4981 28871 5015
rect 28813 4975 28871 4981
rect 1104 4922 40572 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 40572 4922
rect 1104 4848 40572 4870
rect 12066 4768 12072 4820
rect 12124 4808 12130 4820
rect 12345 4811 12403 4817
rect 12345 4808 12357 4811
rect 12124 4780 12357 4808
rect 12124 4768 12130 4780
rect 12345 4777 12357 4780
rect 12391 4777 12403 4811
rect 12345 4771 12403 4777
rect 14274 4768 14280 4820
rect 14332 4768 14338 4820
rect 18966 4808 18972 4820
rect 14660 4780 18972 4808
rect 13906 4700 13912 4752
rect 13964 4740 13970 4752
rect 14660 4740 14688 4780
rect 18966 4768 18972 4780
rect 19024 4768 19030 4820
rect 19061 4811 19119 4817
rect 19061 4777 19073 4811
rect 19107 4808 19119 4811
rect 19702 4808 19708 4820
rect 19107 4780 19708 4808
rect 19107 4777 19119 4780
rect 19061 4771 19119 4777
rect 19702 4768 19708 4780
rect 19760 4808 19766 4820
rect 20530 4808 20536 4820
rect 19760 4780 20536 4808
rect 19760 4768 19766 4780
rect 20530 4768 20536 4780
rect 20588 4768 20594 4820
rect 21177 4811 21235 4817
rect 21177 4777 21189 4811
rect 21223 4808 21235 4811
rect 21450 4808 21456 4820
rect 21223 4780 21456 4808
rect 21223 4777 21235 4780
rect 21177 4771 21235 4777
rect 21450 4768 21456 4780
rect 21508 4768 21514 4820
rect 21560 4780 24808 4808
rect 14918 4740 14924 4752
rect 13964 4712 14688 4740
rect 14752 4712 14924 4740
rect 13964 4700 13970 4712
rect 12986 4632 12992 4684
rect 13044 4632 13050 4684
rect 14752 4681 14780 4712
rect 14918 4700 14924 4712
rect 14976 4700 14982 4752
rect 20622 4700 20628 4752
rect 20680 4740 20686 4752
rect 21560 4740 21588 4780
rect 20680 4712 21588 4740
rect 24780 4740 24808 4780
rect 24780 4712 24900 4740
rect 20680 4700 20686 4712
rect 14737 4675 14795 4681
rect 14737 4641 14749 4675
rect 14783 4641 14795 4675
rect 14737 4635 14795 4641
rect 14829 4675 14887 4681
rect 14829 4641 14841 4675
rect 14875 4672 14887 4675
rect 15010 4672 15016 4684
rect 14875 4644 15016 4672
rect 14875 4641 14887 4644
rect 14829 4635 14887 4641
rect 15010 4632 15016 4644
rect 15068 4632 15074 4684
rect 15194 4632 15200 4684
rect 15252 4672 15258 4684
rect 15289 4675 15347 4681
rect 15289 4672 15301 4675
rect 15252 4644 15301 4672
rect 15252 4632 15258 4644
rect 15289 4641 15301 4644
rect 15335 4641 15347 4675
rect 15289 4635 15347 4641
rect 15565 4675 15623 4681
rect 15565 4641 15577 4675
rect 15611 4672 15623 4675
rect 16574 4672 16580 4684
rect 15611 4644 16580 4672
rect 15611 4641 15623 4644
rect 15565 4635 15623 4641
rect 16574 4632 16580 4644
rect 16632 4632 16638 4684
rect 19245 4675 19303 4681
rect 19245 4672 19257 4675
rect 17328 4644 19257 4672
rect 12250 4564 12256 4616
rect 12308 4564 12314 4616
rect 12342 4564 12348 4616
rect 12400 4604 12406 4616
rect 12713 4607 12771 4613
rect 12713 4604 12725 4607
rect 12400 4576 12725 4604
rect 12400 4564 12406 4576
rect 12713 4573 12725 4576
rect 12759 4573 12771 4607
rect 12713 4567 12771 4573
rect 13814 4564 13820 4616
rect 13872 4604 13878 4616
rect 14274 4604 14280 4616
rect 13872 4576 14280 4604
rect 13872 4564 13878 4576
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 17218 4564 17224 4616
rect 17276 4604 17282 4616
rect 17328 4613 17356 4644
rect 19245 4641 19257 4644
rect 19291 4641 19303 4675
rect 19245 4635 19303 4641
rect 19518 4632 19524 4684
rect 19576 4632 19582 4684
rect 20070 4632 20076 4684
rect 20128 4672 20134 4684
rect 20993 4675 21051 4681
rect 20993 4672 21005 4675
rect 20128 4644 21005 4672
rect 20128 4632 20134 4644
rect 20993 4641 21005 4644
rect 21039 4641 21051 4675
rect 20993 4635 21051 4641
rect 22925 4675 22983 4681
rect 22925 4641 22937 4675
rect 22971 4672 22983 4675
rect 23106 4672 23112 4684
rect 22971 4644 23112 4672
rect 22971 4641 22983 4644
rect 22925 4635 22983 4641
rect 23106 4632 23112 4644
rect 23164 4672 23170 4684
rect 24762 4672 24768 4684
rect 23164 4644 24768 4672
rect 23164 4632 23170 4644
rect 24762 4632 24768 4644
rect 24820 4632 24826 4684
rect 24872 4672 24900 4712
rect 39942 4672 39948 4684
rect 24872 4644 39948 4672
rect 39942 4632 39948 4644
rect 40000 4632 40006 4684
rect 17313 4607 17371 4613
rect 17313 4604 17325 4607
rect 17276 4576 17325 4604
rect 17276 4564 17282 4576
rect 17313 4573 17325 4576
rect 17359 4573 17371 4607
rect 17313 4567 17371 4573
rect 26142 4564 26148 4616
rect 26200 4564 26206 4616
rect 26694 4564 26700 4616
rect 26752 4604 26758 4616
rect 26789 4607 26847 4613
rect 26789 4604 26801 4607
rect 26752 4576 26801 4604
rect 26752 4564 26758 4576
rect 26789 4573 26801 4576
rect 26835 4573 26847 4607
rect 26789 4567 26847 4573
rect 14182 4496 14188 4548
rect 14240 4536 14246 4548
rect 14645 4539 14703 4545
rect 14645 4536 14657 4539
rect 14240 4508 14657 4536
rect 14240 4496 14246 4508
rect 14645 4505 14657 4508
rect 14691 4505 14703 4539
rect 14645 4499 14703 4505
rect 15194 4496 15200 4548
rect 15252 4536 15258 4548
rect 15470 4536 15476 4548
rect 15252 4508 15476 4536
rect 15252 4496 15258 4508
rect 15470 4496 15476 4508
rect 15528 4536 15534 4548
rect 16022 4536 16028 4548
rect 15528 4508 16028 4536
rect 15528 4496 15534 4508
rect 16022 4496 16028 4508
rect 16080 4496 16086 4548
rect 17589 4539 17647 4545
rect 17589 4505 17601 4539
rect 17635 4505 17647 4539
rect 17589 4499 17647 4505
rect 11606 4428 11612 4480
rect 11664 4428 11670 4480
rect 12805 4471 12863 4477
rect 12805 4437 12817 4471
rect 12851 4468 12863 4471
rect 13173 4471 13231 4477
rect 13173 4468 13185 4471
rect 12851 4440 13185 4468
rect 12851 4437 12863 4440
rect 12805 4431 12863 4437
rect 13173 4437 13185 4440
rect 13219 4437 13231 4471
rect 13173 4431 13231 4437
rect 16850 4428 16856 4480
rect 16908 4468 16914 4480
rect 17037 4471 17095 4477
rect 17037 4468 17049 4471
rect 16908 4440 17049 4468
rect 16908 4428 16914 4440
rect 17037 4437 17049 4440
rect 17083 4437 17095 4471
rect 17604 4468 17632 4499
rect 17678 4496 17684 4548
rect 17736 4536 17742 4548
rect 17736 4508 18078 4536
rect 17736 4496 17742 4508
rect 20162 4496 20168 4548
rect 20220 4496 20226 4548
rect 21634 4496 21640 4548
rect 21692 4496 21698 4548
rect 22646 4496 22652 4548
rect 22704 4496 22710 4548
rect 25041 4539 25099 4545
rect 25041 4505 25053 4539
rect 25087 4536 25099 4539
rect 25130 4536 25136 4548
rect 25087 4508 25136 4536
rect 25087 4505 25099 4508
rect 25041 4499 25099 4505
rect 25130 4496 25136 4508
rect 25188 4496 25194 4548
rect 18322 4468 18328 4480
rect 17604 4440 18328 4468
rect 17037 4431 17095 4437
rect 18322 4428 18328 4440
rect 18380 4428 18386 4480
rect 24762 4428 24768 4480
rect 24820 4468 24826 4480
rect 26160 4468 26188 4564
rect 24820 4440 26188 4468
rect 24820 4428 24826 4440
rect 1104 4378 40572 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 40572 4378
rect 1104 4304 40572 4326
rect 11606 4224 11612 4276
rect 11664 4264 11670 4276
rect 11977 4267 12035 4273
rect 11977 4264 11989 4267
rect 11664 4236 11989 4264
rect 11664 4224 11670 4236
rect 11977 4233 11989 4236
rect 12023 4233 12035 4267
rect 11977 4227 12035 4233
rect 12710 4224 12716 4276
rect 12768 4224 12774 4276
rect 16022 4224 16028 4276
rect 16080 4264 16086 4276
rect 16209 4267 16267 4273
rect 16209 4264 16221 4267
rect 16080 4236 16221 4264
rect 16080 4224 16086 4236
rect 16209 4233 16221 4236
rect 16255 4233 16267 4267
rect 16209 4227 16267 4233
rect 17954 4224 17960 4276
rect 18012 4264 18018 4276
rect 20898 4264 20904 4276
rect 18012 4236 20904 4264
rect 18012 4224 18018 4236
rect 11882 4156 11888 4208
rect 11940 4156 11946 4208
rect 16117 4199 16175 4205
rect 16117 4165 16129 4199
rect 16163 4196 16175 4199
rect 16942 4196 16948 4208
rect 16163 4168 16948 4196
rect 16163 4165 16175 4168
rect 16117 4159 16175 4165
rect 16942 4156 16948 4168
rect 17000 4196 17006 4208
rect 17678 4196 17684 4208
rect 17000 4168 17684 4196
rect 17000 4156 17006 4168
rect 17678 4156 17684 4168
rect 17736 4156 17742 4208
rect 19334 4196 19340 4208
rect 18616 4168 19340 4196
rect 12805 4131 12863 4137
rect 12805 4097 12817 4131
rect 12851 4128 12863 4131
rect 14093 4131 14151 4137
rect 14093 4128 14105 4131
rect 12851 4100 14105 4128
rect 12851 4097 12863 4100
rect 12805 4091 12863 4097
rect 14093 4097 14105 4100
rect 14139 4097 14151 4131
rect 14093 4091 14151 4097
rect 16666 4088 16672 4140
rect 16724 4088 16730 4140
rect 18509 4131 18567 4137
rect 18509 4097 18521 4131
rect 18555 4128 18567 4131
rect 18616 4128 18644 4168
rect 19334 4156 19340 4168
rect 19392 4196 19398 4208
rect 19797 4199 19855 4205
rect 19797 4196 19809 4199
rect 19392 4168 19809 4196
rect 19392 4156 19398 4168
rect 19797 4165 19809 4168
rect 19843 4165 19855 4199
rect 19797 4159 19855 4165
rect 20162 4156 20168 4208
rect 20220 4156 20226 4208
rect 20272 4205 20300 4236
rect 20898 4224 20904 4236
rect 20956 4224 20962 4276
rect 21085 4267 21143 4273
rect 21085 4233 21097 4267
rect 21131 4264 21143 4267
rect 21131 4236 21404 4264
rect 21131 4233 21143 4236
rect 21085 4227 21143 4233
rect 20257 4199 20315 4205
rect 20257 4165 20269 4199
rect 20303 4165 20315 4199
rect 20257 4159 20315 4165
rect 21266 4156 21272 4208
rect 21324 4156 21330 4208
rect 21376 4205 21404 4236
rect 22646 4224 22652 4276
rect 22704 4224 22710 4276
rect 23014 4224 23020 4276
rect 23072 4264 23078 4276
rect 29178 4264 29184 4276
rect 23072 4236 29184 4264
rect 23072 4224 23078 4236
rect 29178 4224 29184 4236
rect 29236 4224 29242 4276
rect 21361 4199 21419 4205
rect 21361 4165 21373 4199
rect 21407 4196 21419 4199
rect 21450 4196 21456 4208
rect 21407 4168 21456 4196
rect 21407 4165 21419 4168
rect 21361 4159 21419 4165
rect 21450 4156 21456 4168
rect 21508 4156 21514 4208
rect 23934 4196 23940 4208
rect 21836 4168 23940 4196
rect 18555 4100 18644 4128
rect 18555 4097 18567 4100
rect 18509 4091 18567 4097
rect 18690 4088 18696 4140
rect 18748 4088 18754 4140
rect 18874 4088 18880 4140
rect 18932 4128 18938 4140
rect 18969 4131 19027 4137
rect 18969 4128 18981 4131
rect 18932 4100 18981 4128
rect 18932 4088 18938 4100
rect 18969 4097 18981 4100
rect 19015 4097 19027 4131
rect 18969 4091 19027 4097
rect 19702 4088 19708 4140
rect 19760 4088 19766 4140
rect 19886 4088 19892 4140
rect 19944 4128 19950 4140
rect 19981 4131 20039 4137
rect 19981 4128 19993 4131
rect 19944 4100 19993 4128
rect 19944 4088 19950 4100
rect 19981 4097 19993 4100
rect 20027 4097 20039 4131
rect 19981 4091 20039 4097
rect 20070 4088 20076 4140
rect 20128 4088 20134 4140
rect 12161 4063 12219 4069
rect 12161 4029 12173 4063
rect 12207 4060 12219 4063
rect 12986 4060 12992 4072
rect 12207 4032 12992 4060
rect 12207 4029 12219 4032
rect 12161 4023 12219 4029
rect 12986 4020 12992 4032
rect 13044 4020 13050 4072
rect 13814 4020 13820 4072
rect 13872 4060 13878 4072
rect 13909 4063 13967 4069
rect 13909 4060 13921 4063
rect 13872 4032 13921 4060
rect 13872 4020 13878 4032
rect 13909 4029 13921 4032
rect 13955 4029 13967 4063
rect 13909 4023 13967 4029
rect 13998 4020 14004 4072
rect 14056 4060 14062 4072
rect 14645 4063 14703 4069
rect 14645 4060 14657 4063
rect 14056 4032 14657 4060
rect 14056 4020 14062 4032
rect 14645 4029 14657 4032
rect 14691 4029 14703 4063
rect 14645 4023 14703 4029
rect 15654 4020 15660 4072
rect 15712 4060 15718 4072
rect 15749 4063 15807 4069
rect 15749 4060 15761 4063
rect 15712 4032 15761 4060
rect 15712 4020 15718 4032
rect 15749 4029 15761 4032
rect 15795 4029 15807 4063
rect 15749 4023 15807 4029
rect 16850 4020 16856 4072
rect 16908 4060 16914 4072
rect 17681 4063 17739 4069
rect 17681 4060 17693 4063
rect 16908 4032 17693 4060
rect 16908 4020 16914 4032
rect 17681 4029 17693 4032
rect 17727 4029 17739 4063
rect 17681 4023 17739 4029
rect 18322 4020 18328 4072
rect 18380 4020 18386 4072
rect 18598 4020 18604 4072
rect 18656 4020 18662 4072
rect 18785 4063 18843 4069
rect 18785 4029 18797 4063
rect 18831 4060 18843 4063
rect 19061 4063 19119 4069
rect 19061 4060 19073 4063
rect 18831 4032 19073 4060
rect 18831 4029 18843 4032
rect 18785 4023 18843 4029
rect 19061 4029 19073 4032
rect 19107 4029 19119 4063
rect 19061 4023 19119 4029
rect 13004 3992 13032 4020
rect 15010 3992 15016 4004
rect 13004 3964 15016 3992
rect 15010 3952 15016 3964
rect 15068 3952 15074 4004
rect 19426 3952 19432 4004
rect 19484 3992 19490 4004
rect 19797 3995 19855 4001
rect 19797 3992 19809 3995
rect 19484 3964 19809 3992
rect 19484 3952 19490 3964
rect 19797 3961 19809 3964
rect 19843 3961 19855 3995
rect 19797 3955 19855 3961
rect 11054 3884 11060 3936
rect 11112 3924 11118 3936
rect 11517 3927 11575 3933
rect 11517 3924 11529 3927
rect 11112 3896 11529 3924
rect 11112 3884 11118 3896
rect 11517 3893 11529 3896
rect 11563 3893 11575 3927
rect 11517 3887 11575 3893
rect 11882 3884 11888 3936
rect 11940 3924 11946 3936
rect 12345 3927 12403 3933
rect 12345 3924 12357 3927
rect 11940 3896 12357 3924
rect 11940 3884 11946 3896
rect 12345 3893 12357 3896
rect 12391 3893 12403 3927
rect 12345 3887 12403 3893
rect 12986 3884 12992 3936
rect 13044 3924 13050 3936
rect 13357 3927 13415 3933
rect 13357 3924 13369 3927
rect 13044 3896 13369 3924
rect 13044 3884 13050 3896
rect 13357 3893 13369 3896
rect 13403 3893 13415 3927
rect 13357 3887 13415 3893
rect 14826 3884 14832 3936
rect 14884 3924 14890 3936
rect 15197 3927 15255 3933
rect 15197 3924 15209 3927
rect 14884 3896 15209 3924
rect 14884 3884 14890 3896
rect 15197 3893 15209 3896
rect 15243 3893 15255 3927
rect 15197 3887 15255 3893
rect 16761 3927 16819 3933
rect 16761 3893 16773 3927
rect 16807 3924 16819 3927
rect 17034 3924 17040 3936
rect 16807 3896 17040 3924
rect 16807 3893 16819 3896
rect 16761 3887 16819 3893
rect 17034 3884 17040 3896
rect 17092 3884 17098 3936
rect 17126 3884 17132 3936
rect 17184 3884 17190 3936
rect 18782 3884 18788 3936
rect 18840 3924 18846 3936
rect 20180 3924 20208 4156
rect 21836 4140 21864 4168
rect 23934 4156 23940 4168
rect 23992 4156 23998 4208
rect 30190 4196 30196 4208
rect 29578 4168 30196 4196
rect 30190 4156 30196 4168
rect 30248 4156 30254 4208
rect 20714 4088 20720 4140
rect 20772 4128 20778 4140
rect 20993 4131 21051 4137
rect 20993 4128 21005 4131
rect 20772 4100 21005 4128
rect 20772 4088 20778 4100
rect 20993 4097 21005 4100
rect 21039 4097 21051 4131
rect 20993 4091 21051 4097
rect 21542 4088 21548 4140
rect 21600 4088 21606 4140
rect 21637 4131 21695 4137
rect 21637 4097 21649 4131
rect 21683 4128 21695 4131
rect 21726 4128 21732 4140
rect 21683 4100 21732 4128
rect 21683 4097 21695 4100
rect 21637 4091 21695 4097
rect 21726 4088 21732 4100
rect 21784 4088 21790 4140
rect 21818 4088 21824 4140
rect 21876 4088 21882 4140
rect 21928 4100 22876 4128
rect 21174 4020 21180 4072
rect 21232 4060 21238 4072
rect 21928 4060 21956 4100
rect 22848 4069 22876 4100
rect 23014 4088 23020 4140
rect 23072 4128 23078 4140
rect 23109 4131 23167 4137
rect 23109 4128 23121 4131
rect 23072 4100 23121 4128
rect 23072 4088 23078 4100
rect 23109 4097 23121 4100
rect 23155 4097 23167 4131
rect 23109 4091 23167 4097
rect 23201 4131 23259 4137
rect 23201 4097 23213 4131
rect 23247 4097 23259 4131
rect 23201 4091 23259 4097
rect 21232 4032 21956 4060
rect 22005 4063 22063 4069
rect 21232 4020 21238 4032
rect 22005 4029 22017 4063
rect 22051 4029 22063 4063
rect 22005 4023 22063 4029
rect 22833 4063 22891 4069
rect 22833 4029 22845 4063
rect 22879 4029 22891 4063
rect 23216 4060 23244 4091
rect 23290 4088 23296 4140
rect 23348 4088 23354 4140
rect 23474 4088 23480 4140
rect 23532 4088 23538 4140
rect 28166 4088 28172 4140
rect 28224 4088 28230 4140
rect 28537 4131 28595 4137
rect 28537 4097 28549 4131
rect 28583 4128 28595 4131
rect 28626 4128 28632 4140
rect 28583 4100 28632 4128
rect 28583 4097 28595 4100
rect 28537 4091 28595 4097
rect 28626 4088 28632 4100
rect 28684 4088 28690 4140
rect 23382 4060 23388 4072
rect 23216 4032 23388 4060
rect 22833 4023 22891 4029
rect 21269 3995 21327 4001
rect 21269 3961 21281 3995
rect 21315 3992 21327 3995
rect 22020 3992 22048 4023
rect 23382 4020 23388 4032
rect 23440 4020 23446 4072
rect 21315 3964 22048 3992
rect 21315 3961 21327 3964
rect 21269 3955 21327 3961
rect 29270 3952 29276 4004
rect 29328 3992 29334 4004
rect 29917 3995 29975 4001
rect 29917 3992 29929 3995
rect 29328 3964 29929 3992
rect 29328 3952 29334 3964
rect 29917 3961 29929 3964
rect 29963 3961 29975 3995
rect 29917 3955 29975 3961
rect 20349 3927 20407 3933
rect 20349 3924 20361 3927
rect 18840 3896 20361 3924
rect 18840 3884 18846 3896
rect 20349 3893 20361 3896
rect 20395 3893 20407 3927
rect 20349 3887 20407 3893
rect 21361 3927 21419 3933
rect 21361 3893 21373 3927
rect 21407 3924 21419 3927
rect 22370 3924 22376 3936
rect 21407 3896 22376 3924
rect 21407 3893 21419 3896
rect 21361 3887 21419 3893
rect 22370 3884 22376 3896
rect 22428 3884 22434 3936
rect 1104 3834 40572 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 40572 3834
rect 1104 3760 40572 3782
rect 11606 3680 11612 3732
rect 11664 3720 11670 3732
rect 12250 3720 12256 3732
rect 11664 3692 12256 3720
rect 11664 3680 11670 3692
rect 12250 3680 12256 3692
rect 12308 3720 12314 3732
rect 12437 3723 12495 3729
rect 12437 3720 12449 3723
rect 12308 3692 12449 3720
rect 12308 3680 12314 3692
rect 12437 3689 12449 3692
rect 12483 3689 12495 3723
rect 12437 3683 12495 3689
rect 19889 3723 19947 3729
rect 19889 3689 19901 3723
rect 19935 3720 19947 3723
rect 20070 3720 20076 3732
rect 19935 3692 20076 3720
rect 19935 3689 19947 3692
rect 19889 3683 19947 3689
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 21542 3680 21548 3732
rect 21600 3720 21606 3732
rect 21637 3723 21695 3729
rect 21637 3720 21649 3723
rect 21600 3692 21649 3720
rect 21600 3680 21606 3692
rect 21637 3689 21649 3692
rect 21683 3689 21695 3723
rect 22728 3723 22786 3729
rect 22728 3720 22740 3723
rect 21637 3683 21695 3689
rect 22388 3692 22740 3720
rect 17862 3652 17868 3664
rect 16868 3624 17868 3652
rect 10689 3587 10747 3593
rect 10689 3553 10701 3587
rect 10735 3584 10747 3587
rect 10962 3584 10968 3596
rect 10735 3556 10968 3584
rect 10735 3553 10747 3556
rect 10689 3547 10747 3553
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 12986 3544 12992 3596
rect 13044 3544 13050 3596
rect 13078 3544 13084 3596
rect 13136 3593 13142 3596
rect 13136 3587 13185 3593
rect 13136 3553 13139 3587
rect 13173 3553 13185 3587
rect 13136 3547 13185 3553
rect 13136 3544 13142 3547
rect 14826 3544 14832 3596
rect 14884 3544 14890 3596
rect 15010 3544 15016 3596
rect 15068 3584 15074 3596
rect 16868 3584 16896 3624
rect 17862 3612 17868 3624
rect 17920 3612 17926 3664
rect 15068 3556 16896 3584
rect 17313 3587 17371 3593
rect 15068 3544 15074 3556
rect 17313 3553 17325 3587
rect 17359 3584 17371 3587
rect 17957 3587 18015 3593
rect 17957 3584 17969 3587
rect 17359 3556 17969 3584
rect 17359 3553 17371 3556
rect 17313 3547 17371 3553
rect 17957 3553 17969 3556
rect 18003 3553 18015 3587
rect 17957 3547 18015 3553
rect 12894 3476 12900 3528
rect 12952 3476 12958 3528
rect 13725 3519 13783 3525
rect 13725 3485 13737 3519
rect 13771 3516 13783 3519
rect 13906 3516 13912 3528
rect 13771 3488 13912 3516
rect 13771 3485 13783 3488
rect 13725 3479 13783 3485
rect 13906 3476 13912 3488
rect 13964 3476 13970 3528
rect 14642 3476 14648 3528
rect 14700 3516 14706 3528
rect 14737 3519 14795 3525
rect 14737 3516 14749 3519
rect 14700 3488 14749 3516
rect 14700 3476 14706 3488
rect 14737 3485 14749 3488
rect 14783 3485 14795 3519
rect 14737 3479 14795 3485
rect 15562 3476 15568 3528
rect 15620 3476 15626 3528
rect 16942 3476 16948 3528
rect 17000 3516 17006 3528
rect 18782 3516 18788 3528
rect 17000 3488 18788 3516
rect 17000 3476 17006 3488
rect 18782 3476 18788 3488
rect 18840 3476 18846 3528
rect 19242 3476 19248 3528
rect 19300 3476 19306 3528
rect 21358 3476 21364 3528
rect 21416 3476 21422 3528
rect 21634 3476 21640 3528
rect 21692 3516 21698 3528
rect 22189 3519 22247 3525
rect 22189 3516 22201 3519
rect 21692 3488 22201 3516
rect 21692 3476 21698 3488
rect 22189 3485 22201 3488
rect 22235 3485 22247 3519
rect 22189 3479 22247 3485
rect 10965 3451 11023 3457
rect 10965 3417 10977 3451
rect 11011 3448 11023 3451
rect 11054 3448 11060 3460
rect 11011 3420 11060 3448
rect 11011 3417 11023 3420
rect 10965 3411 11023 3417
rect 11054 3408 11060 3420
rect 11112 3408 11118 3460
rect 13357 3451 13415 3457
rect 13357 3448 13369 3451
rect 11164 3420 11454 3448
rect 12406 3420 13369 3448
rect 10594 3340 10600 3392
rect 10652 3380 10658 3392
rect 11164 3380 11192 3420
rect 12406 3380 12434 3420
rect 13357 3417 13369 3420
rect 13403 3417 13415 3451
rect 13357 3411 13415 3417
rect 15746 3408 15752 3460
rect 15804 3448 15810 3460
rect 15841 3451 15899 3457
rect 15841 3448 15853 3451
rect 15804 3420 15853 3448
rect 15804 3408 15810 3420
rect 15841 3417 15853 3420
rect 15887 3417 15899 3451
rect 15841 3411 15899 3417
rect 21453 3451 21511 3457
rect 21453 3417 21465 3451
rect 21499 3448 21511 3451
rect 22388 3448 22416 3692
rect 22728 3689 22740 3692
rect 22774 3720 22786 3723
rect 22922 3720 22928 3732
rect 22774 3692 22928 3720
rect 22774 3689 22786 3692
rect 22728 3683 22786 3689
rect 22922 3680 22928 3692
rect 22980 3720 22986 3732
rect 23290 3720 23296 3732
rect 22980 3692 23296 3720
rect 22980 3680 22986 3692
rect 23290 3680 23296 3692
rect 23348 3680 23354 3732
rect 39942 3612 39948 3664
rect 40000 3612 40006 3664
rect 22465 3587 22523 3593
rect 22465 3553 22477 3587
rect 22511 3584 22523 3587
rect 22738 3584 22744 3596
rect 22511 3556 22744 3584
rect 22511 3553 22523 3556
rect 22465 3547 22523 3553
rect 22738 3544 22744 3556
rect 22796 3584 22802 3596
rect 23106 3584 23112 3596
rect 22796 3556 23112 3584
rect 22796 3544 22802 3556
rect 23106 3544 23112 3556
rect 23164 3544 23170 3596
rect 24854 3544 24860 3596
rect 24912 3584 24918 3596
rect 26145 3587 26203 3593
rect 26145 3584 26157 3587
rect 24912 3556 26157 3584
rect 24912 3544 24918 3556
rect 26145 3553 26157 3556
rect 26191 3553 26203 3587
rect 26145 3547 26203 3553
rect 24762 3516 24768 3528
rect 23874 3502 24768 3516
rect 21499 3420 22416 3448
rect 23860 3488 24768 3502
rect 21499 3417 21511 3420
rect 21453 3411 21511 3417
rect 10652 3352 12434 3380
rect 10652 3340 10658 3352
rect 12526 3340 12532 3392
rect 12584 3340 12590 3392
rect 14090 3340 14096 3392
rect 14148 3380 14154 3392
rect 14369 3383 14427 3389
rect 14369 3380 14381 3383
rect 14148 3352 14381 3380
rect 14148 3340 14154 3352
rect 14369 3349 14381 3352
rect 14415 3349 14427 3383
rect 14369 3343 14427 3349
rect 17402 3340 17408 3392
rect 17460 3340 17466 3392
rect 21542 3340 21548 3392
rect 21600 3380 21606 3392
rect 23860 3380 23888 3488
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 26786 3476 26792 3528
rect 26844 3476 26850 3528
rect 25869 3451 25927 3457
rect 25869 3417 25881 3451
rect 25915 3448 25927 3451
rect 26237 3451 26295 3457
rect 26237 3448 26249 3451
rect 25915 3420 26249 3448
rect 25915 3417 25927 3420
rect 25869 3411 25927 3417
rect 26237 3417 26249 3420
rect 26283 3417 26295 3451
rect 26237 3411 26295 3417
rect 40126 3408 40132 3460
rect 40184 3408 40190 3460
rect 21600 3352 23888 3380
rect 21600 3340 21606 3352
rect 24210 3340 24216 3392
rect 24268 3340 24274 3392
rect 24302 3340 24308 3392
rect 24360 3380 24366 3392
rect 24397 3383 24455 3389
rect 24397 3380 24409 3383
rect 24360 3352 24409 3380
rect 24360 3340 24366 3352
rect 24397 3349 24409 3352
rect 24443 3349 24455 3383
rect 24397 3343 24455 3349
rect 1104 3290 40572 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 40572 3290
rect 1104 3216 40572 3238
rect 15562 3176 15568 3188
rect 11992 3148 15568 3176
rect 11606 3000 11612 3052
rect 11664 3000 11670 3052
rect 11790 2932 11796 2984
rect 11848 2972 11854 2984
rect 11992 2981 12020 3148
rect 12253 3111 12311 3117
rect 12253 3077 12265 3111
rect 12299 3108 12311 3111
rect 12526 3108 12532 3120
rect 12299 3080 12532 3108
rect 12299 3077 12311 3080
rect 12253 3071 12311 3077
rect 12526 3068 12532 3080
rect 12584 3068 12590 3120
rect 13354 3000 13360 3052
rect 13412 3000 13418 3052
rect 13740 3040 13768 3148
rect 15562 3136 15568 3148
rect 15620 3176 15626 3188
rect 16666 3176 16672 3188
rect 15620 3148 16672 3176
rect 15620 3136 15626 3148
rect 16666 3136 16672 3148
rect 16724 3136 16730 3188
rect 17034 3136 17040 3188
rect 17092 3136 17098 3188
rect 17126 3136 17132 3188
rect 17184 3136 17190 3188
rect 18064 3148 19932 3176
rect 14090 3068 14096 3120
rect 14148 3068 14154 3120
rect 15746 3068 15752 3120
rect 15804 3068 15810 3120
rect 13817 3043 13875 3049
rect 13817 3040 13829 3043
rect 13740 3012 13829 3040
rect 13817 3009 13829 3012
rect 13863 3009 13875 3043
rect 13817 3003 13875 3009
rect 15194 3000 15200 3052
rect 15252 3000 15258 3052
rect 15470 3000 15476 3052
rect 15528 3040 15534 3052
rect 15657 3043 15715 3049
rect 15657 3040 15669 3043
rect 15528 3012 15669 3040
rect 15528 3000 15534 3012
rect 15657 3009 15669 3012
rect 15703 3009 15715 3043
rect 15657 3003 15715 3009
rect 16666 3000 16672 3052
rect 16724 3040 16730 3052
rect 17218 3040 17224 3052
rect 16724 3012 17224 3040
rect 16724 3000 16730 3012
rect 17218 3000 17224 3012
rect 17276 3040 17282 3052
rect 18064 3049 18092 3148
rect 18782 3068 18788 3120
rect 18840 3068 18846 3120
rect 19904 3049 19932 3148
rect 21634 3136 21640 3188
rect 21692 3136 21698 3188
rect 22741 3179 22799 3185
rect 22741 3145 22753 3179
rect 22787 3176 22799 3179
rect 22830 3176 22836 3188
rect 22787 3148 22836 3176
rect 22787 3145 22799 3148
rect 22741 3139 22799 3145
rect 22830 3136 22836 3148
rect 22888 3136 22894 3188
rect 25777 3179 25835 3185
rect 25777 3145 25789 3179
rect 25823 3176 25835 3179
rect 26786 3176 26792 3188
rect 25823 3148 26792 3176
rect 25823 3145 25835 3148
rect 25777 3139 25835 3145
rect 26786 3136 26792 3148
rect 26844 3136 26850 3188
rect 21542 3108 21548 3120
rect 21390 3080 21548 3108
rect 21542 3068 21548 3080
rect 21600 3068 21606 3120
rect 23474 3108 23480 3120
rect 22066 3080 23480 3108
rect 18049 3043 18107 3049
rect 18049 3040 18061 3043
rect 17276 3012 18061 3040
rect 17276 3000 17282 3012
rect 18049 3009 18061 3012
rect 18095 3009 18107 3043
rect 18049 3003 18107 3009
rect 19889 3043 19947 3049
rect 19889 3009 19901 3043
rect 19935 3009 19947 3043
rect 19889 3003 19947 3009
rect 21821 3043 21879 3049
rect 21821 3009 21833 3043
rect 21867 3040 21879 3043
rect 22066 3040 22094 3080
rect 21867 3012 22094 3040
rect 22557 3043 22615 3049
rect 21867 3009 21879 3012
rect 21821 3003 21879 3009
rect 22557 3009 22569 3043
rect 22603 3009 22615 3043
rect 22557 3003 22615 3009
rect 22833 3043 22891 3049
rect 22833 3009 22845 3043
rect 22879 3040 22891 3043
rect 23106 3040 23112 3052
rect 22879 3012 23112 3040
rect 22879 3009 22891 3012
rect 22833 3003 22891 3009
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 11848 2944 11989 2972
rect 11848 2932 11854 2944
rect 11977 2941 11989 2944
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 12802 2932 12808 2984
rect 12860 2972 12866 2984
rect 13372 2972 13400 3000
rect 12860 2944 13400 2972
rect 17313 2975 17371 2981
rect 12860 2932 12866 2944
rect 17313 2941 17325 2975
rect 17359 2972 17371 2975
rect 17862 2972 17868 2984
rect 17359 2944 17868 2972
rect 17359 2941 17371 2944
rect 17313 2935 17371 2941
rect 17862 2932 17868 2944
rect 17920 2932 17926 2984
rect 18325 2975 18383 2981
rect 18325 2941 18337 2975
rect 18371 2972 18383 2975
rect 19334 2972 19340 2984
rect 18371 2944 19340 2972
rect 18371 2941 18383 2944
rect 18325 2935 18383 2941
rect 19334 2932 19340 2944
rect 19392 2932 19398 2984
rect 20162 2932 20168 2984
rect 20220 2932 20226 2984
rect 20806 2932 20812 2984
rect 20864 2972 20870 2984
rect 21836 2972 21864 3003
rect 20864 2944 21864 2972
rect 20864 2932 20870 2944
rect 21910 2932 21916 2984
rect 21968 2972 21974 2984
rect 22189 2975 22247 2981
rect 22189 2972 22201 2975
rect 21968 2944 22201 2972
rect 21968 2932 21974 2944
rect 22189 2941 22201 2944
rect 22235 2941 22247 2975
rect 22189 2935 22247 2941
rect 22462 2932 22468 2984
rect 22520 2972 22526 2984
rect 22572 2972 22600 3003
rect 23106 3000 23112 3012
rect 23164 3000 23170 3052
rect 23216 3049 23244 3080
rect 23474 3068 23480 3080
rect 23532 3068 23538 3120
rect 23934 3068 23940 3120
rect 23992 3068 23998 3120
rect 24210 3068 24216 3120
rect 24268 3108 24274 3120
rect 24489 3111 24547 3117
rect 24489 3108 24501 3111
rect 24268 3080 24501 3108
rect 24268 3068 24274 3080
rect 24489 3077 24501 3080
rect 24535 3108 24547 3111
rect 24535 3080 24624 3108
rect 24535 3077 24547 3080
rect 24489 3071 24547 3077
rect 23201 3043 23259 3049
rect 23201 3009 23213 3043
rect 23247 3009 23259 3043
rect 23201 3003 23259 3009
rect 24302 3000 24308 3052
rect 24360 3000 24366 3052
rect 24596 3049 24624 3080
rect 24581 3043 24639 3049
rect 24581 3009 24593 3043
rect 24627 3009 24639 3043
rect 24581 3003 24639 3009
rect 23382 2972 23388 2984
rect 22520 2944 23388 2972
rect 22520 2932 22526 2944
rect 23382 2932 23388 2944
rect 23440 2972 23446 2984
rect 23477 2975 23535 2981
rect 23477 2972 23489 2975
rect 23440 2944 23489 2972
rect 23440 2932 23446 2944
rect 23477 2941 23489 2944
rect 23523 2941 23535 2975
rect 24320 2972 24348 3000
rect 25317 2975 25375 2981
rect 25317 2972 25329 2975
rect 24320 2944 25329 2972
rect 23477 2935 23535 2941
rect 25317 2941 25329 2944
rect 25363 2941 25375 2975
rect 25317 2935 25375 2941
rect 13725 2907 13783 2913
rect 13725 2873 13737 2907
rect 13771 2904 13783 2907
rect 13814 2904 13820 2916
rect 13771 2876 13820 2904
rect 13771 2873 13783 2876
rect 13725 2867 13783 2873
rect 13814 2864 13820 2876
rect 13872 2864 13878 2916
rect 15565 2907 15623 2913
rect 15565 2873 15577 2907
rect 15611 2904 15623 2907
rect 15654 2904 15660 2916
rect 15611 2876 15660 2904
rect 15611 2873 15623 2876
rect 15565 2867 15623 2873
rect 15654 2864 15660 2876
rect 15712 2864 15718 2916
rect 16574 2864 16580 2916
rect 16632 2904 16638 2916
rect 16669 2907 16727 2913
rect 16669 2904 16681 2907
rect 16632 2876 16681 2904
rect 16632 2864 16638 2876
rect 16669 2873 16681 2876
rect 16715 2873 16727 2907
rect 16669 2867 16727 2873
rect 25225 2907 25283 2913
rect 25225 2873 25237 2907
rect 25271 2904 25283 2907
rect 25593 2907 25651 2913
rect 25593 2904 25605 2907
rect 25271 2876 25605 2904
rect 25271 2873 25283 2876
rect 25225 2867 25283 2873
rect 25593 2873 25605 2876
rect 25639 2873 25651 2907
rect 25593 2867 25651 2873
rect 11793 2839 11851 2845
rect 11793 2805 11805 2839
rect 11839 2836 11851 2839
rect 12342 2836 12348 2848
rect 11839 2808 12348 2836
rect 11839 2805 11851 2808
rect 11793 2799 11851 2805
rect 12342 2796 12348 2808
rect 12400 2796 12406 2848
rect 19794 2796 19800 2848
rect 19852 2796 19858 2848
rect 1104 2746 40572 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 40572 2746
rect 1104 2672 40572 2694
rect 18877 2635 18935 2641
rect 18877 2601 18889 2635
rect 18923 2632 18935 2635
rect 19242 2632 19248 2644
rect 18923 2604 19248 2632
rect 18923 2601 18935 2604
rect 18877 2595 18935 2601
rect 19242 2592 19248 2604
rect 19300 2592 19306 2644
rect 19334 2592 19340 2644
rect 19392 2592 19398 2644
rect 20162 2592 20168 2644
rect 20220 2632 20226 2644
rect 20625 2635 20683 2641
rect 20625 2632 20637 2635
rect 20220 2604 20637 2632
rect 20220 2592 20226 2604
rect 20625 2601 20637 2604
rect 20671 2601 20683 2635
rect 20625 2595 20683 2601
rect 12894 2524 12900 2576
rect 12952 2564 12958 2576
rect 13449 2567 13507 2573
rect 13449 2564 13461 2567
rect 12952 2536 13461 2564
rect 12952 2524 12958 2536
rect 13449 2533 13461 2536
rect 13495 2533 13507 2567
rect 13449 2527 13507 2533
rect 13538 2524 13544 2576
rect 13596 2564 13602 2576
rect 15473 2567 15531 2573
rect 15473 2564 15485 2567
rect 13596 2536 15485 2564
rect 13596 2524 13602 2536
rect 15473 2533 15485 2536
rect 15519 2533 15531 2567
rect 15473 2527 15531 2533
rect 21177 2567 21235 2573
rect 21177 2533 21189 2567
rect 21223 2533 21235 2567
rect 21177 2527 21235 2533
rect 11517 2499 11575 2505
rect 11517 2465 11529 2499
rect 11563 2496 11575 2499
rect 11790 2496 11796 2508
rect 11563 2468 11796 2496
rect 11563 2465 11575 2468
rect 11517 2459 11575 2465
rect 11790 2456 11796 2468
rect 11848 2456 11854 2508
rect 13265 2499 13323 2505
rect 13265 2465 13277 2499
rect 13311 2465 13323 2499
rect 15378 2496 15384 2508
rect 13265 2459 13323 2465
rect 15212 2468 15384 2496
rect 11330 2388 11336 2440
rect 11388 2388 11394 2440
rect 13280 2428 13308 2459
rect 13633 2431 13691 2437
rect 13633 2428 13645 2431
rect 13280 2400 13645 2428
rect 13633 2397 13645 2400
rect 13679 2428 13691 2431
rect 13998 2428 14004 2440
rect 13679 2400 14004 2428
rect 13679 2397 13691 2400
rect 13633 2391 13691 2397
rect 13998 2388 14004 2400
rect 14056 2388 14062 2440
rect 14274 2388 14280 2440
rect 14332 2388 14338 2440
rect 15212 2437 15240 2468
rect 15378 2456 15384 2468
rect 15436 2456 15442 2508
rect 16666 2456 16672 2508
rect 16724 2496 16730 2508
rect 17129 2499 17187 2505
rect 17129 2496 17141 2499
rect 16724 2468 17141 2496
rect 16724 2456 16730 2468
rect 17129 2465 17141 2468
rect 17175 2465 17187 2499
rect 17129 2459 17187 2465
rect 17402 2456 17408 2508
rect 17460 2456 17466 2508
rect 19794 2456 19800 2508
rect 19852 2496 19858 2508
rect 19981 2499 20039 2505
rect 19981 2496 19993 2499
rect 19852 2468 19993 2496
rect 19852 2456 19858 2468
rect 19981 2465 19993 2468
rect 20027 2465 20039 2499
rect 19981 2459 20039 2465
rect 15197 2431 15255 2437
rect 15197 2397 15209 2431
rect 15243 2397 15255 2431
rect 15197 2391 15255 2397
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2397 15347 2431
rect 15289 2391 15347 2397
rect 11793 2363 11851 2369
rect 11793 2329 11805 2363
rect 11839 2360 11851 2363
rect 11882 2360 11888 2372
rect 11839 2332 11888 2360
rect 11839 2329 11851 2332
rect 11793 2323 11851 2329
rect 11882 2320 11888 2332
rect 11940 2320 11946 2372
rect 12802 2320 12808 2372
rect 12860 2320 12866 2372
rect 13814 2320 13820 2372
rect 13872 2360 13878 2372
rect 15304 2360 15332 2391
rect 15562 2388 15568 2440
rect 15620 2428 15626 2440
rect 16209 2431 16267 2437
rect 16209 2428 16221 2431
rect 15620 2400 16221 2428
rect 15620 2388 15626 2400
rect 16209 2397 16221 2400
rect 16255 2397 16267 2431
rect 16209 2391 16267 2397
rect 16850 2388 16856 2440
rect 16908 2428 16914 2440
rect 17037 2431 17095 2437
rect 17037 2428 17049 2431
rect 16908 2400 17049 2428
rect 16908 2388 16914 2400
rect 17037 2397 17049 2400
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 19392 2400 19441 2428
rect 19392 2388 19398 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 20622 2388 20628 2440
rect 20680 2428 20686 2440
rect 20993 2431 21051 2437
rect 20993 2428 21005 2431
rect 20680 2400 21005 2428
rect 20680 2388 20686 2400
rect 20993 2397 21005 2400
rect 21039 2397 21051 2431
rect 21192 2428 21220 2527
rect 22738 2456 22744 2508
rect 22796 2496 22802 2508
rect 23201 2499 23259 2505
rect 23201 2496 23213 2499
rect 22796 2468 23213 2496
rect 22796 2456 22802 2468
rect 23201 2465 23213 2468
rect 23247 2465 23259 2499
rect 23201 2459 23259 2465
rect 21361 2431 21419 2437
rect 21361 2428 21373 2431
rect 21192 2400 21373 2428
rect 20993 2391 21051 2397
rect 21361 2397 21373 2400
rect 21407 2397 21419 2431
rect 21361 2391 21419 2397
rect 23014 2388 23020 2440
rect 23072 2428 23078 2440
rect 23385 2431 23443 2437
rect 23385 2428 23397 2431
rect 23072 2400 23397 2428
rect 23072 2388 23078 2400
rect 23385 2397 23397 2400
rect 23431 2397 23443 2431
rect 23385 2391 23443 2397
rect 13872 2332 15332 2360
rect 13872 2320 13878 2332
rect 17954 2320 17960 2372
rect 18012 2320 18018 2372
rect 20714 2320 20720 2372
rect 20772 2360 20778 2372
rect 21085 2363 21143 2369
rect 21085 2360 21097 2363
rect 20772 2332 21097 2360
rect 20772 2320 20778 2332
rect 21085 2329 21097 2332
rect 21131 2329 21143 2363
rect 21085 2323 21143 2329
rect 21269 2363 21327 2369
rect 21269 2329 21281 2363
rect 21315 2360 21327 2363
rect 22462 2360 22468 2372
rect 21315 2332 22468 2360
rect 21315 2329 21327 2332
rect 21269 2323 21327 2329
rect 22462 2320 22468 2332
rect 22520 2320 22526 2372
rect 11149 2295 11207 2301
rect 11149 2261 11161 2295
rect 11195 2292 11207 2295
rect 11606 2292 11612 2304
rect 11195 2264 11612 2292
rect 11195 2261 11207 2264
rect 11149 2255 11207 2261
rect 11606 2252 11612 2264
rect 11664 2252 11670 2304
rect 14182 2252 14188 2304
rect 14240 2292 14246 2304
rect 14461 2295 14519 2301
rect 14461 2292 14473 2295
rect 14240 2264 14473 2292
rect 14240 2252 14246 2264
rect 14461 2261 14473 2264
rect 14507 2261 14519 2295
rect 14461 2255 14519 2261
rect 14826 2252 14832 2304
rect 14884 2292 14890 2304
rect 15013 2295 15071 2301
rect 15013 2292 15025 2295
rect 14884 2264 15025 2292
rect 14884 2252 14890 2264
rect 15013 2261 15025 2264
rect 15059 2261 15071 2295
rect 15013 2255 15071 2261
rect 16114 2252 16120 2304
rect 16172 2292 16178 2304
rect 16393 2295 16451 2301
rect 16393 2292 16405 2295
rect 16172 2264 16405 2292
rect 16172 2252 16178 2264
rect 16393 2261 16405 2264
rect 16439 2261 16451 2295
rect 16393 2255 16451 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 16853 2295 16911 2301
rect 16853 2292 16865 2295
rect 16816 2264 16865 2292
rect 16816 2252 16822 2264
rect 16853 2261 16865 2264
rect 16899 2261 16911 2295
rect 16853 2255 16911 2261
rect 21358 2252 21364 2304
rect 21416 2292 21422 2304
rect 21545 2295 21603 2301
rect 21545 2292 21557 2295
rect 21416 2264 21557 2292
rect 21416 2252 21422 2264
rect 21545 2261 21557 2264
rect 21591 2261 21603 2295
rect 21545 2255 21603 2261
rect 23569 2295 23627 2301
rect 23569 2261 23581 2295
rect 23615 2292 23627 2295
rect 23842 2292 23848 2304
rect 23615 2264 23848 2292
rect 23615 2261 23627 2264
rect 23569 2255 23627 2261
rect 23842 2252 23848 2264
rect 23900 2252 23906 2304
rect 1104 2202 40572 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 40572 2202
rect 1104 2128 40572 2150
<< via1 >>
rect 4874 41318 4926 41370
rect 4938 41318 4990 41370
rect 5002 41318 5054 41370
rect 5066 41318 5118 41370
rect 5130 41318 5182 41370
rect 35594 41318 35646 41370
rect 35658 41318 35710 41370
rect 35722 41318 35774 41370
rect 35786 41318 35838 41370
rect 35850 41318 35902 41370
rect 30932 41080 30984 41132
rect 31208 41055 31260 41064
rect 31208 41021 31217 41055
rect 31217 41021 31251 41055
rect 31251 41021 31260 41055
rect 31208 41012 31260 41021
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 17040 40604 17092 40656
rect 15016 40536 15068 40588
rect 15752 40511 15804 40520
rect 15752 40477 15761 40511
rect 15761 40477 15795 40511
rect 15795 40477 15804 40511
rect 15752 40468 15804 40477
rect 16396 40468 16448 40520
rect 16580 40511 16632 40520
rect 16580 40477 16589 40511
rect 16589 40477 16623 40511
rect 16623 40477 16632 40511
rect 16580 40468 16632 40477
rect 15936 40332 15988 40384
rect 16488 40375 16540 40384
rect 16488 40341 16497 40375
rect 16497 40341 16531 40375
rect 16531 40341 16540 40375
rect 16488 40332 16540 40341
rect 4874 40230 4926 40282
rect 4938 40230 4990 40282
rect 5002 40230 5054 40282
rect 5066 40230 5118 40282
rect 5130 40230 5182 40282
rect 35594 40230 35646 40282
rect 35658 40230 35710 40282
rect 35722 40230 35774 40282
rect 35786 40230 35838 40282
rect 35850 40230 35902 40282
rect 13452 40103 13504 40112
rect 13452 40069 13461 40103
rect 13461 40069 13495 40103
rect 13495 40069 13504 40103
rect 13452 40060 13504 40069
rect 15476 40128 15528 40180
rect 12256 39924 12308 39976
rect 12164 39788 12216 39840
rect 12532 39788 12584 39840
rect 13636 40035 13688 40044
rect 13636 40001 13645 40035
rect 13645 40001 13679 40035
rect 13679 40001 13688 40035
rect 13636 39992 13688 40001
rect 15016 40035 15068 40044
rect 15016 40001 15025 40035
rect 15025 40001 15059 40035
rect 15059 40001 15068 40035
rect 15016 39992 15068 40001
rect 14464 39924 14516 39976
rect 15568 39992 15620 40044
rect 16396 39992 16448 40044
rect 17132 39992 17184 40044
rect 14280 39899 14332 39908
rect 14280 39865 14289 39899
rect 14289 39865 14323 39899
rect 14323 39865 14332 39899
rect 14280 39856 14332 39865
rect 15752 39856 15804 39908
rect 16304 39924 16356 39976
rect 16856 39856 16908 39908
rect 17868 39856 17920 39908
rect 15200 39831 15252 39840
rect 15200 39797 15209 39831
rect 15209 39797 15243 39831
rect 15243 39797 15252 39831
rect 15200 39788 15252 39797
rect 16396 39831 16448 39840
rect 16396 39797 16405 39831
rect 16405 39797 16439 39831
rect 16439 39797 16448 39831
rect 16396 39788 16448 39797
rect 16948 39788 17000 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 11980 39627 12032 39636
rect 8484 39448 8536 39500
rect 8392 39380 8444 39432
rect 9404 39380 9456 39432
rect 11244 39423 11296 39432
rect 11244 39389 11253 39423
rect 11253 39389 11287 39423
rect 11287 39389 11296 39423
rect 11244 39380 11296 39389
rect 11980 39593 11989 39627
rect 11989 39593 12023 39627
rect 12023 39593 12032 39627
rect 11980 39584 12032 39593
rect 12072 39516 12124 39568
rect 11520 39423 11572 39432
rect 11520 39389 11529 39423
rect 11529 39389 11563 39423
rect 11563 39389 11572 39423
rect 11520 39380 11572 39389
rect 12164 39423 12216 39432
rect 12164 39389 12173 39423
rect 12173 39389 12207 39423
rect 12207 39389 12216 39423
rect 12164 39380 12216 39389
rect 15292 39584 15344 39636
rect 16396 39584 16448 39636
rect 15568 39516 15620 39568
rect 16488 39516 16540 39568
rect 13636 39448 13688 39500
rect 8300 39244 8352 39296
rect 11060 39244 11112 39296
rect 11612 39287 11664 39296
rect 11612 39253 11621 39287
rect 11621 39253 11655 39287
rect 11655 39253 11664 39287
rect 11612 39244 11664 39253
rect 11980 39244 12032 39296
rect 14464 39423 14516 39432
rect 14464 39389 14473 39423
rect 14473 39389 14507 39423
rect 14507 39389 14516 39423
rect 14464 39380 14516 39389
rect 15200 39380 15252 39432
rect 15936 39448 15988 39500
rect 17040 39491 17092 39500
rect 17040 39457 17049 39491
rect 17049 39457 17083 39491
rect 17083 39457 17092 39491
rect 17040 39448 17092 39457
rect 15844 39423 15896 39432
rect 15844 39389 15853 39423
rect 15853 39389 15887 39423
rect 15887 39389 15896 39423
rect 15844 39380 15896 39389
rect 15476 39312 15528 39364
rect 16212 39380 16264 39432
rect 16580 39380 16632 39432
rect 17132 39423 17184 39432
rect 17132 39389 17141 39423
rect 17141 39389 17175 39423
rect 17175 39389 17184 39423
rect 17868 39448 17920 39500
rect 17132 39380 17184 39389
rect 12992 39244 13044 39296
rect 14648 39287 14700 39296
rect 14648 39253 14657 39287
rect 14657 39253 14691 39287
rect 14691 39253 14700 39287
rect 14648 39244 14700 39253
rect 15844 39244 15896 39296
rect 15936 39244 15988 39296
rect 18052 39312 18104 39364
rect 16672 39244 16724 39296
rect 17960 39244 18012 39296
rect 4874 39142 4926 39194
rect 4938 39142 4990 39194
rect 5002 39142 5054 39194
rect 5066 39142 5118 39194
rect 5130 39142 5182 39194
rect 35594 39142 35646 39194
rect 35658 39142 35710 39194
rect 35722 39142 35774 39194
rect 35786 39142 35838 39194
rect 35850 39142 35902 39194
rect 10876 39040 10928 39092
rect 11980 39083 12032 39092
rect 11980 39049 11989 39083
rect 11989 39049 12023 39083
rect 12023 39049 12032 39083
rect 11980 39040 12032 39049
rect 12072 39083 12124 39092
rect 12072 39049 12081 39083
rect 12081 39049 12115 39083
rect 12115 39049 12124 39083
rect 12072 39040 12124 39049
rect 14648 39040 14700 39092
rect 15016 39040 15068 39092
rect 20720 39040 20772 39092
rect 10232 38947 10284 38956
rect 10232 38913 10241 38947
rect 10241 38913 10275 38947
rect 10275 38913 10284 38947
rect 10232 38904 10284 38913
rect 11612 38972 11664 39024
rect 6828 38836 6880 38888
rect 8576 38879 8628 38888
rect 8576 38845 8585 38879
rect 8585 38845 8619 38879
rect 8619 38845 8628 38879
rect 8576 38836 8628 38845
rect 9312 38836 9364 38888
rect 11060 38947 11112 38956
rect 11060 38913 11069 38947
rect 11069 38913 11103 38947
rect 11103 38913 11112 38947
rect 11060 38904 11112 38913
rect 16672 39015 16724 39024
rect 16672 38981 16681 39015
rect 16681 38981 16715 39015
rect 16715 38981 16724 39015
rect 16672 38972 16724 38981
rect 18052 39015 18104 39024
rect 18052 38981 18061 39015
rect 18061 38981 18095 39015
rect 18095 38981 18104 39015
rect 18052 38972 18104 38981
rect 18328 38972 18380 39024
rect 20812 38972 20864 39024
rect 23204 38972 23256 39024
rect 24492 38972 24544 39024
rect 27068 38972 27120 39024
rect 12256 38947 12308 38956
rect 12256 38913 12265 38947
rect 12265 38913 12299 38947
rect 12299 38913 12308 38947
rect 12256 38904 12308 38913
rect 16948 38947 17000 38956
rect 16948 38913 16957 38947
rect 16957 38913 16991 38947
rect 16991 38913 17000 38947
rect 16948 38904 17000 38913
rect 25228 38904 25280 38956
rect 9588 38768 9640 38820
rect 10508 38836 10560 38888
rect 12440 38879 12492 38888
rect 12440 38845 12449 38879
rect 12449 38845 12483 38879
rect 12483 38845 12492 38879
rect 12440 38836 12492 38845
rect 19800 38879 19852 38888
rect 19800 38845 19809 38879
rect 19809 38845 19843 38879
rect 19843 38845 19852 38879
rect 19800 38836 19852 38845
rect 20076 38879 20128 38888
rect 20076 38845 20085 38879
rect 20085 38845 20119 38879
rect 20119 38845 20128 38879
rect 20076 38836 20128 38845
rect 23020 38836 23072 38888
rect 25504 38879 25556 38888
rect 25504 38845 25513 38879
rect 25513 38845 25547 38879
rect 25547 38845 25556 38879
rect 25504 38836 25556 38845
rect 9956 38700 10008 38752
rect 10140 38700 10192 38752
rect 10600 38743 10652 38752
rect 10600 38709 10609 38743
rect 10609 38709 10643 38743
rect 10643 38709 10652 38743
rect 10600 38700 10652 38709
rect 19064 38700 19116 38752
rect 27436 38700 27488 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 8392 38496 8444 38548
rect 8576 38496 8628 38548
rect 9404 38539 9456 38548
rect 9404 38505 9413 38539
rect 9413 38505 9447 38539
rect 9447 38505 9456 38539
rect 9404 38496 9456 38505
rect 10232 38496 10284 38548
rect 10508 38539 10560 38548
rect 10508 38505 10517 38539
rect 10517 38505 10551 38539
rect 10551 38505 10560 38539
rect 10508 38496 10560 38505
rect 11520 38539 11572 38548
rect 11520 38505 11529 38539
rect 11529 38505 11563 38539
rect 11563 38505 11572 38539
rect 11520 38496 11572 38505
rect 13452 38496 13504 38548
rect 15200 38496 15252 38548
rect 19800 38496 19852 38548
rect 19892 38496 19944 38548
rect 8576 38360 8628 38412
rect 8852 38428 8904 38480
rect 5448 38335 5500 38344
rect 5448 38301 5457 38335
rect 5457 38301 5491 38335
rect 5491 38301 5500 38335
rect 5448 38292 5500 38301
rect 5724 38335 5776 38344
rect 5724 38301 5733 38335
rect 5733 38301 5767 38335
rect 5767 38301 5776 38335
rect 5724 38292 5776 38301
rect 8024 38335 8076 38344
rect 8024 38301 8033 38335
rect 8033 38301 8067 38335
rect 8067 38301 8076 38335
rect 8024 38292 8076 38301
rect 8116 38335 8168 38344
rect 8116 38301 8125 38335
rect 8125 38301 8159 38335
rect 8159 38301 8168 38335
rect 8116 38292 8168 38301
rect 8300 38335 8352 38344
rect 8300 38301 8309 38335
rect 8309 38301 8343 38335
rect 8343 38301 8352 38335
rect 8300 38292 8352 38301
rect 8392 38335 8444 38344
rect 8392 38301 8401 38335
rect 8401 38301 8435 38335
rect 8435 38301 8444 38335
rect 8392 38292 8444 38301
rect 7012 38224 7064 38276
rect 8668 38292 8720 38344
rect 9036 38335 9088 38344
rect 9036 38301 9045 38335
rect 9045 38301 9079 38335
rect 9079 38301 9088 38335
rect 9036 38292 9088 38301
rect 9312 38360 9364 38412
rect 9588 38292 9640 38344
rect 10232 38335 10284 38344
rect 10232 38301 10241 38335
rect 10241 38301 10275 38335
rect 10275 38301 10284 38335
rect 10232 38292 10284 38301
rect 11336 38335 11388 38344
rect 11336 38301 11345 38335
rect 11345 38301 11379 38335
rect 11379 38301 11388 38335
rect 11336 38292 11388 38301
rect 12256 38292 12308 38344
rect 12624 38335 12676 38344
rect 12624 38301 12633 38335
rect 12633 38301 12667 38335
rect 12667 38301 12676 38335
rect 12624 38292 12676 38301
rect 12992 38403 13044 38412
rect 12992 38369 13001 38403
rect 13001 38369 13035 38403
rect 13035 38369 13044 38403
rect 12992 38360 13044 38369
rect 13452 38360 13504 38412
rect 13176 38335 13228 38344
rect 13176 38301 13185 38335
rect 13185 38301 13219 38335
rect 13219 38301 13228 38335
rect 13176 38292 13228 38301
rect 4436 38156 4488 38208
rect 12440 38224 12492 38276
rect 20628 38428 20680 38480
rect 20812 38428 20864 38480
rect 21272 38471 21324 38480
rect 16580 38360 16632 38412
rect 21272 38437 21281 38471
rect 21281 38437 21315 38471
rect 21315 38437 21324 38471
rect 21272 38428 21324 38437
rect 17776 38335 17828 38344
rect 17776 38301 17785 38335
rect 17785 38301 17819 38335
rect 17819 38301 17828 38335
rect 17776 38292 17828 38301
rect 17960 38335 18012 38344
rect 17960 38301 17969 38335
rect 17969 38301 18003 38335
rect 18003 38301 18012 38335
rect 17960 38292 18012 38301
rect 18052 38335 18104 38344
rect 18052 38301 18061 38335
rect 18061 38301 18095 38335
rect 18095 38301 18104 38335
rect 18052 38292 18104 38301
rect 18328 38335 18380 38344
rect 18328 38301 18337 38335
rect 18337 38301 18371 38335
rect 18371 38301 18380 38335
rect 18328 38292 18380 38301
rect 19248 38292 19300 38344
rect 18512 38224 18564 38276
rect 11244 38156 11296 38208
rect 12808 38156 12860 38208
rect 13268 38156 13320 38208
rect 14832 38156 14884 38208
rect 18328 38156 18380 38208
rect 19340 38156 19392 38208
rect 21180 38292 21232 38344
rect 22100 38292 22152 38344
rect 23204 38539 23256 38548
rect 23204 38505 23213 38539
rect 23213 38505 23247 38539
rect 23247 38505 23256 38539
rect 23204 38496 23256 38505
rect 25504 38360 25556 38412
rect 26424 38360 26476 38412
rect 27068 38360 27120 38412
rect 27436 38360 27488 38412
rect 23020 38292 23072 38344
rect 28908 38292 28960 38344
rect 21456 38156 21508 38208
rect 21640 38199 21692 38208
rect 21640 38165 21649 38199
rect 21649 38165 21683 38199
rect 21683 38165 21692 38199
rect 21640 38156 21692 38165
rect 24492 38224 24544 38276
rect 24952 38224 25004 38276
rect 25320 38224 25372 38276
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 35594 38054 35646 38106
rect 35658 38054 35710 38106
rect 35722 38054 35774 38106
rect 35786 38054 35838 38106
rect 35850 38054 35902 38106
rect 4436 37927 4488 37936
rect 4436 37893 4445 37927
rect 4445 37893 4479 37927
rect 4479 37893 4488 37927
rect 4436 37884 4488 37893
rect 7012 37952 7064 38004
rect 8668 37995 8720 38004
rect 8668 37961 8677 37995
rect 8677 37961 8711 37995
rect 8711 37961 8720 37995
rect 8668 37952 8720 37961
rect 12808 37952 12860 38004
rect 13176 37952 13228 38004
rect 5908 37816 5960 37868
rect 8944 37816 8996 37868
rect 5540 37612 5592 37664
rect 6644 37791 6696 37800
rect 6644 37757 6653 37791
rect 6653 37757 6687 37791
rect 6687 37757 6696 37791
rect 6644 37748 6696 37757
rect 9312 37859 9364 37868
rect 9312 37825 9321 37859
rect 9321 37825 9355 37859
rect 9355 37825 9364 37859
rect 9312 37816 9364 37825
rect 13268 37927 13320 37936
rect 13268 37893 13277 37927
rect 13277 37893 13311 37927
rect 13311 37893 13320 37927
rect 13268 37884 13320 37893
rect 15016 37884 15068 37936
rect 17776 37952 17828 38004
rect 14832 37816 14884 37868
rect 6828 37612 6880 37664
rect 7932 37612 7984 37664
rect 9128 37612 9180 37664
rect 15200 37748 15252 37800
rect 15384 37816 15436 37868
rect 15844 37859 15896 37868
rect 15844 37825 15853 37859
rect 15853 37825 15887 37859
rect 15887 37825 15896 37859
rect 15844 37816 15896 37825
rect 17408 37816 17460 37868
rect 17684 37859 17736 37868
rect 17684 37825 17693 37859
rect 17693 37825 17727 37859
rect 17727 37825 17736 37859
rect 17684 37816 17736 37825
rect 17316 37748 17368 37800
rect 19248 37884 19300 37936
rect 18144 37816 18196 37868
rect 18972 37859 19024 37868
rect 18972 37825 18981 37859
rect 18981 37825 19015 37859
rect 19015 37825 19024 37859
rect 18972 37816 19024 37825
rect 19156 37859 19208 37868
rect 19156 37825 19165 37859
rect 19165 37825 19199 37859
rect 19199 37825 19208 37859
rect 19156 37816 19208 37825
rect 19340 37859 19392 37868
rect 19340 37825 19349 37859
rect 19349 37825 19383 37859
rect 19383 37825 19392 37859
rect 19340 37816 19392 37825
rect 20076 37952 20128 38004
rect 22376 37952 22428 38004
rect 20628 37884 20680 37936
rect 24952 37995 25004 38004
rect 24952 37961 24961 37995
rect 24961 37961 24995 37995
rect 24995 37961 25004 37995
rect 24952 37952 25004 37961
rect 26424 37952 26476 38004
rect 18052 37748 18104 37800
rect 19248 37791 19300 37800
rect 19248 37757 19257 37791
rect 19257 37757 19291 37791
rect 19291 37757 19300 37791
rect 19248 37748 19300 37757
rect 15568 37680 15620 37732
rect 16764 37680 16816 37732
rect 21548 37816 21600 37868
rect 22100 37859 22152 37868
rect 22100 37825 22109 37859
rect 22109 37825 22143 37859
rect 22143 37825 22152 37859
rect 22100 37816 22152 37825
rect 21824 37791 21876 37800
rect 21824 37757 21833 37791
rect 21833 37757 21867 37791
rect 21867 37757 21876 37791
rect 21824 37748 21876 37757
rect 25228 37816 25280 37868
rect 22376 37791 22428 37800
rect 22376 37757 22385 37791
rect 22385 37757 22419 37791
rect 22419 37757 22428 37791
rect 22376 37748 22428 37757
rect 22652 37791 22704 37800
rect 22652 37757 22661 37791
rect 22661 37757 22695 37791
rect 22695 37757 22704 37791
rect 22652 37748 22704 37757
rect 23848 37748 23900 37800
rect 25504 37791 25556 37800
rect 25504 37757 25513 37791
rect 25513 37757 25547 37791
rect 25547 37757 25556 37791
rect 25504 37748 25556 37757
rect 13728 37612 13780 37664
rect 15292 37612 15344 37664
rect 18604 37612 18656 37664
rect 21456 37612 21508 37664
rect 21916 37655 21968 37664
rect 21916 37621 21925 37655
rect 21925 37621 21959 37655
rect 21959 37621 21968 37655
rect 21916 37612 21968 37621
rect 23020 37612 23072 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 6644 37408 6696 37460
rect 8116 37408 8168 37460
rect 8852 37408 8904 37460
rect 12624 37408 12676 37460
rect 15384 37408 15436 37460
rect 17316 37451 17368 37460
rect 17316 37417 17325 37451
rect 17325 37417 17359 37451
rect 17359 37417 17368 37451
rect 17316 37408 17368 37417
rect 17684 37408 17736 37460
rect 19156 37408 19208 37460
rect 21824 37408 21876 37460
rect 22652 37408 22704 37460
rect 7012 37340 7064 37392
rect 8208 37340 8260 37392
rect 14832 37340 14884 37392
rect 17408 37383 17460 37392
rect 17408 37349 17417 37383
rect 17417 37349 17451 37383
rect 17451 37349 17460 37383
rect 17408 37340 17460 37349
rect 18052 37340 18104 37392
rect 5448 37204 5500 37256
rect 5632 37247 5684 37256
rect 5632 37213 5641 37247
rect 5641 37213 5675 37247
rect 5675 37213 5684 37247
rect 5632 37204 5684 37213
rect 6000 37247 6052 37256
rect 6000 37213 6009 37247
rect 6009 37213 6043 37247
rect 6043 37213 6052 37247
rect 6000 37204 6052 37213
rect 8024 37272 8076 37324
rect 8484 37272 8536 37324
rect 8668 37272 8720 37324
rect 12164 37272 12216 37324
rect 7840 37204 7892 37256
rect 8392 37247 8444 37256
rect 8392 37213 8401 37247
rect 8401 37213 8435 37247
rect 8435 37213 8444 37247
rect 8392 37204 8444 37213
rect 8852 37204 8904 37256
rect 9128 37247 9180 37256
rect 9128 37213 9137 37247
rect 9137 37213 9171 37247
rect 9171 37213 9180 37247
rect 9128 37204 9180 37213
rect 5816 37068 5868 37120
rect 8024 37136 8076 37188
rect 8484 37136 8536 37188
rect 9404 37247 9456 37256
rect 9404 37213 9413 37247
rect 9413 37213 9447 37247
rect 9447 37213 9456 37247
rect 9404 37204 9456 37213
rect 12440 37315 12492 37324
rect 12440 37281 12449 37315
rect 12449 37281 12483 37315
rect 12483 37281 12492 37315
rect 12440 37272 12492 37281
rect 15292 37315 15344 37324
rect 15292 37281 15301 37315
rect 15301 37281 15335 37315
rect 15335 37281 15344 37315
rect 15292 37272 15344 37281
rect 15660 37272 15712 37324
rect 12348 37204 12400 37256
rect 12532 37247 12584 37256
rect 12532 37213 12541 37247
rect 12541 37213 12575 37247
rect 12575 37213 12584 37247
rect 12532 37204 12584 37213
rect 12624 37247 12676 37256
rect 12624 37213 12633 37247
rect 12633 37213 12667 37247
rect 12667 37213 12676 37247
rect 12624 37204 12676 37213
rect 14188 37204 14240 37256
rect 14648 37204 14700 37256
rect 14740 37247 14792 37256
rect 14740 37213 14749 37247
rect 14749 37213 14783 37247
rect 14783 37213 14792 37247
rect 14740 37204 14792 37213
rect 17224 37315 17276 37324
rect 17224 37281 17233 37315
rect 17233 37281 17267 37315
rect 17267 37281 17276 37315
rect 17224 37272 17276 37281
rect 12256 37111 12308 37120
rect 12256 37077 12265 37111
rect 12265 37077 12299 37111
rect 12299 37077 12308 37111
rect 12256 37068 12308 37077
rect 13820 37136 13872 37188
rect 17684 37204 17736 37256
rect 17776 37247 17828 37256
rect 17776 37213 17785 37247
rect 17785 37213 17819 37247
rect 17819 37213 17828 37247
rect 17776 37204 17828 37213
rect 17960 37204 18012 37256
rect 18236 37204 18288 37256
rect 17868 37136 17920 37188
rect 18604 37315 18656 37324
rect 18604 37281 18613 37315
rect 18613 37281 18647 37315
rect 18647 37281 18656 37315
rect 18604 37272 18656 37281
rect 19064 37272 19116 37324
rect 21548 37340 21600 37392
rect 22100 37340 22152 37392
rect 19340 37204 19392 37256
rect 19708 37247 19760 37256
rect 19708 37213 19717 37247
rect 19717 37213 19751 37247
rect 19751 37213 19760 37247
rect 19708 37204 19760 37213
rect 21640 37272 21692 37324
rect 23848 37340 23900 37392
rect 25504 37272 25556 37324
rect 25964 37315 26016 37324
rect 25964 37281 25973 37315
rect 25973 37281 26007 37315
rect 26007 37281 26016 37315
rect 25964 37272 26016 37281
rect 21272 37247 21324 37256
rect 21272 37213 21281 37247
rect 21281 37213 21315 37247
rect 21315 37213 21324 37247
rect 21272 37204 21324 37213
rect 21456 37247 21508 37256
rect 21456 37213 21465 37247
rect 21465 37213 21499 37247
rect 21499 37213 21508 37247
rect 21456 37204 21508 37213
rect 14004 37068 14056 37120
rect 15660 37068 15712 37120
rect 16028 37068 16080 37120
rect 18696 37068 18748 37120
rect 19432 37111 19484 37120
rect 19432 37077 19441 37111
rect 19441 37077 19475 37111
rect 19475 37077 19484 37111
rect 19432 37068 19484 37077
rect 19892 37136 19944 37188
rect 27712 37204 27764 37256
rect 22560 37136 22612 37188
rect 25044 37068 25096 37120
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 6000 36907 6052 36916
rect 6000 36873 6009 36907
rect 6009 36873 6043 36907
rect 6043 36873 6052 36907
rect 6000 36864 6052 36873
rect 8392 36864 8444 36916
rect 9772 36864 9824 36916
rect 10876 36864 10928 36916
rect 11704 36864 11756 36916
rect 12348 36864 12400 36916
rect 12624 36864 12676 36916
rect 9128 36796 9180 36848
rect 10600 36796 10652 36848
rect 5448 36728 5500 36780
rect 5816 36771 5868 36780
rect 5816 36737 5825 36771
rect 5825 36737 5859 36771
rect 5859 36737 5868 36771
rect 5816 36728 5868 36737
rect 6368 36771 6420 36780
rect 6368 36737 6377 36771
rect 6377 36737 6411 36771
rect 6411 36737 6420 36771
rect 6368 36728 6420 36737
rect 8300 36728 8352 36780
rect 8484 36771 8536 36780
rect 8484 36737 8493 36771
rect 8493 36737 8527 36771
rect 8527 36737 8536 36771
rect 8484 36728 8536 36737
rect 8852 36728 8904 36780
rect 9404 36728 9456 36780
rect 10692 36771 10744 36780
rect 10692 36737 10701 36771
rect 10701 36737 10735 36771
rect 10735 36737 10744 36771
rect 10692 36728 10744 36737
rect 6092 36660 6144 36712
rect 8024 36660 8076 36712
rect 11152 36728 11204 36780
rect 11336 36660 11388 36712
rect 11980 36660 12032 36712
rect 3976 36592 4028 36644
rect 9220 36592 9272 36644
rect 12716 36796 12768 36848
rect 13176 36796 13228 36848
rect 15200 36864 15252 36916
rect 15660 36907 15712 36916
rect 15660 36873 15669 36907
rect 15669 36873 15703 36907
rect 15703 36873 15712 36907
rect 15660 36864 15712 36873
rect 16120 36864 16172 36916
rect 13084 36728 13136 36780
rect 13544 36771 13596 36780
rect 13544 36737 13553 36771
rect 13553 36737 13587 36771
rect 13587 36737 13596 36771
rect 13544 36728 13596 36737
rect 14280 36796 14332 36848
rect 14004 36771 14056 36780
rect 14004 36737 14013 36771
rect 14013 36737 14047 36771
rect 14047 36737 14056 36771
rect 18236 36907 18288 36916
rect 18236 36873 18245 36907
rect 18245 36873 18279 36907
rect 18279 36873 18288 36907
rect 18236 36864 18288 36873
rect 18972 36907 19024 36916
rect 18972 36873 18981 36907
rect 18981 36873 19015 36907
rect 19015 36873 19024 36907
rect 18972 36864 19024 36873
rect 24952 36864 25004 36916
rect 25320 36864 25372 36916
rect 14004 36728 14056 36737
rect 15200 36771 15252 36780
rect 15200 36737 15209 36771
rect 15209 36737 15243 36771
rect 15243 36737 15252 36771
rect 15200 36728 15252 36737
rect 15292 36728 15344 36780
rect 16028 36728 16080 36780
rect 16120 36771 16172 36780
rect 16120 36737 16129 36771
rect 16129 36737 16163 36771
rect 16163 36737 16172 36771
rect 16120 36728 16172 36737
rect 20720 36796 20772 36848
rect 25044 36839 25096 36848
rect 25044 36805 25053 36839
rect 25053 36805 25087 36839
rect 25087 36805 25096 36839
rect 25044 36796 25096 36805
rect 27712 36796 27764 36848
rect 17132 36771 17184 36780
rect 17132 36737 17141 36771
rect 17141 36737 17175 36771
rect 17175 36737 17184 36771
rect 17132 36728 17184 36737
rect 17960 36728 18012 36780
rect 18052 36771 18104 36780
rect 18052 36737 18061 36771
rect 18061 36737 18095 36771
rect 18095 36737 18104 36771
rect 18052 36728 18104 36737
rect 18696 36771 18748 36780
rect 18696 36737 18705 36771
rect 18705 36737 18739 36771
rect 18739 36737 18748 36771
rect 18696 36728 18748 36737
rect 23756 36771 23808 36780
rect 23756 36737 23765 36771
rect 23765 36737 23799 36771
rect 23799 36737 23808 36771
rect 23756 36728 23808 36737
rect 12256 36703 12308 36712
rect 12256 36669 12265 36703
rect 12265 36669 12299 36703
rect 12299 36669 12308 36703
rect 12256 36660 12308 36669
rect 14188 36703 14240 36712
rect 14188 36669 14197 36703
rect 14197 36669 14231 36703
rect 14231 36669 14240 36703
rect 14188 36660 14240 36669
rect 5632 36524 5684 36576
rect 9128 36524 9180 36576
rect 10600 36524 10652 36576
rect 12900 36592 12952 36644
rect 11520 36524 11572 36576
rect 17776 36660 17828 36712
rect 19432 36660 19484 36712
rect 23020 36703 23072 36712
rect 23020 36669 23029 36703
rect 23029 36669 23063 36703
rect 23063 36669 23072 36703
rect 23020 36660 23072 36669
rect 24768 36703 24820 36712
rect 24768 36669 24777 36703
rect 24777 36669 24811 36703
rect 24811 36669 24820 36703
rect 24768 36660 24820 36669
rect 17960 36592 18012 36644
rect 20628 36592 20680 36644
rect 14556 36524 14608 36576
rect 15016 36524 15068 36576
rect 18788 36567 18840 36576
rect 18788 36533 18797 36567
rect 18797 36533 18831 36567
rect 18831 36533 18840 36567
rect 18788 36524 18840 36533
rect 19340 36524 19392 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 5448 36320 5500 36372
rect 3976 36159 4028 36168
rect 3976 36125 3985 36159
rect 3985 36125 4019 36159
rect 4019 36125 4028 36159
rect 3976 36116 4028 36125
rect 4620 36116 4672 36168
rect 5724 36116 5776 36168
rect 7472 36320 7524 36372
rect 7840 36363 7892 36372
rect 7840 36329 7849 36363
rect 7849 36329 7883 36363
rect 7883 36329 7892 36363
rect 7840 36320 7892 36329
rect 6368 36116 6420 36168
rect 5816 36048 5868 36100
rect 6276 36091 6328 36100
rect 6276 36057 6285 36091
rect 6285 36057 6319 36091
rect 6319 36057 6328 36091
rect 6276 36048 6328 36057
rect 7288 36159 7340 36168
rect 7288 36125 7297 36159
rect 7297 36125 7331 36159
rect 7331 36125 7340 36159
rect 7288 36116 7340 36125
rect 8576 36320 8628 36372
rect 12164 36320 12216 36372
rect 14740 36320 14792 36372
rect 18052 36320 18104 36372
rect 2964 35980 3016 36032
rect 4252 35980 4304 36032
rect 7564 36091 7616 36100
rect 7564 36057 7573 36091
rect 7573 36057 7607 36091
rect 7607 36057 7616 36091
rect 7564 36048 7616 36057
rect 7748 36048 7800 36100
rect 8208 36116 8260 36168
rect 9496 36252 9548 36304
rect 13084 36252 13136 36304
rect 8576 36184 8628 36236
rect 9128 36159 9180 36168
rect 9128 36125 9137 36159
rect 9137 36125 9171 36159
rect 9171 36125 9180 36159
rect 9128 36116 9180 36125
rect 9220 36159 9272 36168
rect 9220 36125 9229 36159
rect 9229 36125 9263 36159
rect 9263 36125 9272 36159
rect 9220 36116 9272 36125
rect 9680 36116 9732 36168
rect 9956 36184 10008 36236
rect 10692 36184 10744 36236
rect 11612 36184 11664 36236
rect 11888 36184 11940 36236
rect 10140 36048 10192 36100
rect 10416 35980 10468 36032
rect 10600 36091 10652 36100
rect 10600 36057 10609 36091
rect 10609 36057 10643 36091
rect 10643 36057 10652 36091
rect 10600 36048 10652 36057
rect 10876 36048 10928 36100
rect 11612 35980 11664 36032
rect 11980 36116 12032 36168
rect 12440 36091 12492 36100
rect 12440 36057 12449 36091
rect 12449 36057 12483 36091
rect 12483 36057 12492 36091
rect 12440 36048 12492 36057
rect 12716 36159 12768 36168
rect 12716 36125 12725 36159
rect 12725 36125 12759 36159
rect 12759 36125 12768 36159
rect 12716 36116 12768 36125
rect 14556 36227 14608 36236
rect 14556 36193 14565 36227
rect 14565 36193 14599 36227
rect 14599 36193 14608 36227
rect 14556 36184 14608 36193
rect 14832 36184 14884 36236
rect 15292 36295 15344 36304
rect 15292 36261 15301 36295
rect 15301 36261 15335 36295
rect 15335 36261 15344 36295
rect 15292 36252 15344 36261
rect 15200 36184 15252 36236
rect 13544 36048 13596 36100
rect 15660 36252 15712 36304
rect 15844 36227 15896 36236
rect 15844 36193 15853 36227
rect 15853 36193 15887 36227
rect 15887 36193 15896 36227
rect 15844 36184 15896 36193
rect 17224 36184 17276 36236
rect 16120 36048 16172 36100
rect 13360 35980 13412 36032
rect 13728 35980 13780 36032
rect 15476 35980 15528 36032
rect 15844 35980 15896 36032
rect 16396 36116 16448 36168
rect 18788 36184 18840 36236
rect 19248 36184 19300 36236
rect 18236 36116 18288 36168
rect 19616 36159 19668 36168
rect 19616 36125 19625 36159
rect 19625 36125 19659 36159
rect 19659 36125 19668 36159
rect 19616 36116 19668 36125
rect 16304 36048 16356 36100
rect 17132 35980 17184 36032
rect 17960 35980 18012 36032
rect 19892 36091 19944 36100
rect 19892 36057 19901 36091
rect 19901 36057 19935 36091
rect 19935 36057 19944 36091
rect 19892 36048 19944 36057
rect 20628 36048 20680 36100
rect 24768 36184 24820 36236
rect 25780 36184 25832 36236
rect 25964 36184 26016 36236
rect 27160 36227 27212 36236
rect 27160 36193 27169 36227
rect 27169 36193 27203 36227
rect 27203 36193 27212 36227
rect 27160 36184 27212 36193
rect 28356 36184 28408 36236
rect 21916 36159 21968 36168
rect 21916 36125 21925 36159
rect 21925 36125 21959 36159
rect 21959 36125 21968 36159
rect 21916 36116 21968 36125
rect 22284 36159 22336 36168
rect 22284 36125 22293 36159
rect 22293 36125 22327 36159
rect 22327 36125 22336 36159
rect 22284 36116 22336 36125
rect 22468 36159 22520 36168
rect 22468 36125 22477 36159
rect 22477 36125 22511 36159
rect 22511 36125 22520 36159
rect 22468 36116 22520 36125
rect 23020 36116 23072 36168
rect 21364 36023 21416 36032
rect 21364 35989 21373 36023
rect 21373 35989 21407 36023
rect 21407 35989 21416 36023
rect 21364 35980 21416 35989
rect 25136 36048 25188 36100
rect 25412 36091 25464 36100
rect 25412 36057 25421 36091
rect 25421 36057 25455 36091
rect 25455 36057 25464 36091
rect 25412 36048 25464 36057
rect 30472 36048 30524 36100
rect 22560 35980 22612 36032
rect 23480 36023 23532 36032
rect 23480 35989 23489 36023
rect 23489 35989 23523 36023
rect 23523 35989 23532 36023
rect 23480 35980 23532 35989
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 5632 35776 5684 35828
rect 6000 35776 6052 35828
rect 7564 35819 7616 35828
rect 7564 35785 7573 35819
rect 7573 35785 7607 35819
rect 7607 35785 7616 35819
rect 7564 35776 7616 35785
rect 8852 35819 8904 35828
rect 8852 35785 8861 35819
rect 8861 35785 8895 35819
rect 8895 35785 8904 35819
rect 8852 35776 8904 35785
rect 9036 35819 9088 35828
rect 9036 35785 9045 35819
rect 9045 35785 9079 35819
rect 9079 35785 9088 35819
rect 9036 35776 9088 35785
rect 1308 35708 1360 35760
rect 2964 35708 3016 35760
rect 3792 35708 3844 35760
rect 4252 35751 4304 35760
rect 4252 35717 4261 35751
rect 4261 35717 4295 35751
rect 4295 35717 4304 35751
rect 4252 35708 4304 35717
rect 5448 35708 5500 35760
rect 8024 35708 8076 35760
rect 2228 35640 2280 35692
rect 5540 35640 5592 35692
rect 5816 35572 5868 35624
rect 3148 35436 3200 35488
rect 5816 35436 5868 35488
rect 6184 35640 6236 35692
rect 6552 35504 6604 35556
rect 7012 35640 7064 35692
rect 7564 35640 7616 35692
rect 7748 35640 7800 35692
rect 8576 35708 8628 35760
rect 10600 35708 10652 35760
rect 11060 35776 11112 35828
rect 11888 35776 11940 35828
rect 12532 35776 12584 35828
rect 11520 35708 11572 35760
rect 6736 35572 6788 35624
rect 8392 35572 8444 35624
rect 9036 35640 9088 35692
rect 9312 35683 9364 35692
rect 9312 35649 9321 35683
rect 9321 35649 9355 35683
rect 9355 35649 9364 35683
rect 9312 35640 9364 35649
rect 9404 35640 9456 35692
rect 9680 35640 9732 35692
rect 10508 35683 10560 35692
rect 10508 35649 10517 35683
rect 10517 35649 10551 35683
rect 10551 35649 10560 35683
rect 10508 35640 10560 35649
rect 7380 35504 7432 35556
rect 7196 35436 7248 35488
rect 9128 35436 9180 35488
rect 10416 35572 10468 35624
rect 10968 35683 11020 35692
rect 10968 35649 10977 35683
rect 10977 35649 11011 35683
rect 11011 35649 11020 35683
rect 10968 35640 11020 35649
rect 11704 35683 11756 35692
rect 11704 35649 11713 35683
rect 11713 35649 11747 35683
rect 11747 35649 11756 35683
rect 11704 35640 11756 35649
rect 12440 35640 12492 35692
rect 12808 35640 12860 35692
rect 13820 35708 13872 35760
rect 15016 35708 15068 35760
rect 15108 35640 15160 35692
rect 16304 35776 16356 35828
rect 17316 35776 17368 35828
rect 17960 35708 18012 35760
rect 10140 35436 10192 35488
rect 10600 35436 10652 35488
rect 13728 35615 13780 35624
rect 13728 35581 13737 35615
rect 13737 35581 13771 35615
rect 13771 35581 13780 35615
rect 13728 35572 13780 35581
rect 15476 35615 15528 35624
rect 15476 35581 15485 35615
rect 15485 35581 15519 35615
rect 15519 35581 15528 35615
rect 15476 35572 15528 35581
rect 15844 35683 15896 35692
rect 15844 35649 15853 35683
rect 15853 35649 15887 35683
rect 15887 35649 15896 35683
rect 15844 35640 15896 35649
rect 16028 35640 16080 35692
rect 16120 35615 16172 35624
rect 16120 35581 16129 35615
rect 16129 35581 16163 35615
rect 16163 35581 16172 35615
rect 16120 35572 16172 35581
rect 16672 35572 16724 35624
rect 17500 35640 17552 35692
rect 18512 35776 18564 35828
rect 19064 35776 19116 35828
rect 19432 35776 19484 35828
rect 19892 35776 19944 35828
rect 18512 35683 18564 35692
rect 18512 35649 18521 35683
rect 18521 35649 18555 35683
rect 18555 35649 18564 35683
rect 18512 35640 18564 35649
rect 17960 35615 18012 35624
rect 17960 35581 17969 35615
rect 17969 35581 18003 35615
rect 18003 35581 18012 35615
rect 17960 35572 18012 35581
rect 18052 35615 18104 35624
rect 18052 35581 18061 35615
rect 18061 35581 18095 35615
rect 18095 35581 18104 35615
rect 18052 35572 18104 35581
rect 11152 35547 11204 35556
rect 11152 35513 11161 35547
rect 11161 35513 11195 35547
rect 11195 35513 11204 35547
rect 11152 35504 11204 35513
rect 16212 35504 16264 35556
rect 16304 35504 16356 35556
rect 17408 35504 17460 35556
rect 19248 35683 19300 35692
rect 19248 35649 19257 35683
rect 19257 35649 19291 35683
rect 19291 35649 19300 35683
rect 19248 35640 19300 35649
rect 19432 35683 19484 35692
rect 19432 35649 19441 35683
rect 19441 35649 19475 35683
rect 19475 35649 19484 35683
rect 19432 35640 19484 35649
rect 19524 35640 19576 35692
rect 19800 35640 19852 35692
rect 21364 35708 21416 35760
rect 22468 35776 22520 35828
rect 21916 35708 21968 35760
rect 23480 35776 23532 35828
rect 25412 35776 25464 35828
rect 27160 35776 27212 35828
rect 24952 35708 25004 35760
rect 25136 35708 25188 35760
rect 19156 35572 19208 35624
rect 22008 35640 22060 35692
rect 23020 35683 23072 35692
rect 23020 35649 23029 35683
rect 23029 35649 23063 35683
rect 23063 35649 23072 35683
rect 23020 35640 23072 35649
rect 21272 35572 21324 35624
rect 11244 35436 11296 35488
rect 13544 35436 13596 35488
rect 14740 35436 14792 35488
rect 15844 35436 15896 35488
rect 18236 35436 18288 35488
rect 21456 35479 21508 35488
rect 21456 35445 21465 35479
rect 21465 35445 21499 35479
rect 21499 35445 21508 35479
rect 21456 35436 21508 35445
rect 21640 35504 21692 35556
rect 25872 35615 25924 35624
rect 25872 35581 25881 35615
rect 25881 35581 25915 35615
rect 25915 35581 25924 35615
rect 25872 35572 25924 35581
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 5448 35232 5500 35284
rect 6736 35232 6788 35284
rect 7748 35275 7800 35284
rect 7748 35241 7757 35275
rect 7757 35241 7791 35275
rect 7791 35241 7800 35275
rect 7748 35232 7800 35241
rect 9312 35232 9364 35284
rect 16120 35232 16172 35284
rect 16672 35275 16724 35284
rect 16672 35241 16681 35275
rect 16681 35241 16715 35275
rect 16715 35241 16724 35275
rect 16672 35232 16724 35241
rect 9036 35164 9088 35216
rect 3148 35139 3200 35148
rect 3148 35105 3157 35139
rect 3157 35105 3191 35139
rect 3191 35105 3200 35139
rect 3148 35096 3200 35105
rect 5540 35096 5592 35148
rect 6000 35139 6052 35148
rect 6000 35105 6009 35139
rect 6009 35105 6043 35139
rect 6043 35105 6052 35139
rect 6000 35096 6052 35105
rect 6460 35139 6512 35148
rect 6460 35105 6469 35139
rect 6469 35105 6503 35139
rect 6503 35105 6512 35139
rect 6460 35096 6512 35105
rect 6552 35096 6604 35148
rect 6644 35028 6696 35080
rect 8392 35096 8444 35148
rect 8760 35139 8812 35148
rect 8760 35105 8769 35139
rect 8769 35105 8803 35139
rect 8803 35105 8812 35139
rect 11244 35164 11296 35216
rect 17040 35207 17092 35216
rect 17040 35173 17049 35207
rect 17049 35173 17083 35207
rect 17083 35173 17092 35207
rect 17040 35164 17092 35173
rect 17408 35164 17460 35216
rect 8760 35096 8812 35105
rect 13084 35096 13136 35148
rect 13452 35096 13504 35148
rect 16304 35139 16356 35148
rect 16304 35105 16313 35139
rect 16313 35105 16347 35139
rect 16347 35105 16356 35139
rect 16304 35096 16356 35105
rect 17500 35096 17552 35148
rect 1308 34960 1360 35012
rect 2688 34960 2740 35012
rect 5908 34892 5960 34944
rect 6552 34892 6604 34944
rect 7104 35071 7156 35080
rect 7104 35037 7113 35071
rect 7113 35037 7147 35071
rect 7147 35037 7156 35071
rect 7104 35028 7156 35037
rect 7196 35071 7248 35080
rect 7196 35037 7205 35071
rect 7205 35037 7239 35071
rect 7239 35037 7248 35071
rect 7196 35028 7248 35037
rect 7380 35071 7432 35080
rect 7380 35037 7389 35071
rect 7389 35037 7423 35071
rect 7423 35037 7432 35071
rect 7380 35028 7432 35037
rect 7472 35028 7524 35080
rect 8024 35071 8076 35080
rect 8024 35037 8033 35071
rect 8033 35037 8067 35071
rect 8067 35037 8076 35071
rect 8024 35028 8076 35037
rect 8208 35071 8260 35080
rect 8208 35037 8217 35071
rect 8217 35037 8251 35071
rect 8251 35037 8260 35071
rect 8208 35028 8260 35037
rect 8116 34960 8168 35012
rect 9036 35028 9088 35080
rect 9128 35071 9180 35080
rect 9128 35037 9137 35071
rect 9137 35037 9171 35071
rect 9171 35037 9180 35071
rect 9128 35028 9180 35037
rect 9404 35071 9456 35080
rect 9404 35037 9413 35071
rect 9413 35037 9447 35071
rect 9447 35037 9456 35071
rect 9404 35028 9456 35037
rect 12256 35071 12308 35080
rect 12256 35037 12265 35071
rect 12265 35037 12299 35071
rect 12299 35037 12308 35071
rect 12256 35028 12308 35037
rect 12440 35071 12492 35080
rect 12440 35037 12449 35071
rect 12449 35037 12483 35071
rect 12483 35037 12492 35071
rect 12440 35028 12492 35037
rect 12900 35071 12952 35080
rect 12900 35037 12909 35071
rect 12909 35037 12943 35071
rect 12943 35037 12952 35071
rect 12900 35028 12952 35037
rect 16856 35028 16908 35080
rect 17684 35071 17736 35080
rect 17684 35037 17693 35071
rect 17693 35037 17727 35071
rect 17727 35037 17736 35071
rect 17684 35028 17736 35037
rect 17960 35028 18012 35080
rect 19248 35232 19300 35284
rect 20812 35232 20864 35284
rect 22284 35275 22336 35284
rect 18512 35164 18564 35216
rect 18880 35164 18932 35216
rect 19708 35207 19760 35216
rect 19708 35173 19717 35207
rect 19717 35173 19751 35207
rect 19751 35173 19760 35207
rect 19708 35164 19760 35173
rect 22284 35241 22293 35275
rect 22293 35241 22327 35275
rect 22327 35241 22336 35275
rect 22284 35232 22336 35241
rect 21640 35164 21692 35216
rect 19892 35071 19944 35080
rect 19892 35037 19901 35071
rect 19901 35037 19935 35071
rect 19935 35037 19944 35071
rect 19892 35028 19944 35037
rect 20536 35028 20588 35080
rect 21272 35139 21324 35148
rect 21272 35105 21281 35139
rect 21281 35105 21315 35139
rect 21315 35105 21324 35139
rect 21272 35096 21324 35105
rect 21732 35096 21784 35148
rect 20996 35028 21048 35080
rect 11888 34960 11940 35012
rect 15660 34960 15712 35012
rect 15844 34960 15896 35012
rect 16396 34960 16448 35012
rect 16672 34960 16724 35012
rect 10784 34892 10836 34944
rect 11336 34892 11388 34944
rect 12348 34892 12400 34944
rect 17316 35003 17368 35012
rect 17316 34969 17325 35003
rect 17325 34969 17359 35003
rect 17359 34969 17368 35003
rect 17316 34960 17368 34969
rect 17776 35003 17828 35012
rect 17776 34969 17785 35003
rect 17785 34969 17819 35003
rect 17819 34969 17828 35003
rect 17776 34960 17828 34969
rect 18696 34960 18748 35012
rect 22468 35071 22520 35080
rect 22468 35037 22477 35071
rect 22477 35037 22511 35071
rect 22511 35037 22520 35071
rect 22468 35028 22520 35037
rect 17500 34892 17552 34944
rect 18512 34935 18564 34944
rect 18512 34901 18521 34935
rect 18521 34901 18555 34935
rect 18555 34901 18564 34935
rect 18512 34892 18564 34901
rect 18788 34892 18840 34944
rect 19708 34892 19760 34944
rect 20904 34935 20956 34944
rect 20904 34901 20913 34935
rect 20913 34901 20947 34935
rect 20947 34901 20956 34935
rect 20904 34892 20956 34901
rect 21180 34892 21232 34944
rect 22560 34960 22612 35012
rect 22928 35003 22980 35012
rect 22928 34969 22937 35003
rect 22937 34969 22971 35003
rect 22971 34969 22980 35003
rect 22928 34960 22980 34969
rect 22836 34935 22888 34944
rect 22836 34901 22845 34935
rect 22845 34901 22879 34935
rect 22879 34901 22888 34935
rect 22836 34892 22888 34901
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 2688 34688 2740 34740
rect 7104 34688 7156 34740
rect 9404 34688 9456 34740
rect 5908 34620 5960 34672
rect 6184 34620 6236 34672
rect 5540 34552 5592 34604
rect 6092 34552 6144 34604
rect 6552 34595 6604 34604
rect 6552 34561 6561 34595
rect 6561 34561 6595 34595
rect 6595 34561 6604 34595
rect 6552 34552 6604 34561
rect 6644 34595 6696 34604
rect 6644 34561 6653 34595
rect 6653 34561 6687 34595
rect 6687 34561 6696 34595
rect 6644 34552 6696 34561
rect 8208 34620 8260 34672
rect 8484 34620 8536 34672
rect 2320 34527 2372 34536
rect 2320 34493 2329 34527
rect 2329 34493 2363 34527
rect 2363 34493 2372 34527
rect 2320 34484 2372 34493
rect 4068 34527 4120 34536
rect 4068 34493 4077 34527
rect 4077 34493 4111 34527
rect 4111 34493 4120 34527
rect 4068 34484 4120 34493
rect 6828 34484 6880 34536
rect 6092 34416 6144 34468
rect 7104 34416 7156 34468
rect 8576 34552 8628 34604
rect 11428 34620 11480 34672
rect 8944 34552 8996 34604
rect 8484 34484 8536 34536
rect 9588 34552 9640 34604
rect 10140 34595 10192 34604
rect 10140 34561 10149 34595
rect 10149 34561 10183 34595
rect 10183 34561 10192 34595
rect 10140 34552 10192 34561
rect 10600 34595 10652 34604
rect 10600 34561 10609 34595
rect 10609 34561 10643 34595
rect 10643 34561 10652 34595
rect 10600 34552 10652 34561
rect 10784 34552 10836 34604
rect 11060 34595 11112 34604
rect 11060 34561 11069 34595
rect 11069 34561 11103 34595
rect 11103 34561 11112 34595
rect 11060 34552 11112 34561
rect 11244 34595 11296 34604
rect 11244 34561 11252 34595
rect 11252 34561 11286 34595
rect 11286 34561 11296 34595
rect 11244 34552 11296 34561
rect 11336 34595 11388 34604
rect 11336 34561 11345 34595
rect 11345 34561 11379 34595
rect 11379 34561 11388 34595
rect 11336 34552 11388 34561
rect 11888 34595 11940 34604
rect 11888 34561 11897 34595
rect 11897 34561 11931 34595
rect 11931 34561 11940 34595
rect 11888 34552 11940 34561
rect 10324 34527 10376 34536
rect 10324 34493 10333 34527
rect 10333 34493 10367 34527
rect 10367 34493 10376 34527
rect 10324 34484 10376 34493
rect 10692 34484 10744 34536
rect 13820 34688 13872 34740
rect 17408 34731 17460 34740
rect 17408 34697 17417 34731
rect 17417 34697 17451 34731
rect 17451 34697 17460 34731
rect 17408 34688 17460 34697
rect 17500 34688 17552 34740
rect 15016 34620 15068 34672
rect 17776 34620 17828 34672
rect 18512 34688 18564 34740
rect 18788 34688 18840 34740
rect 15292 34552 15344 34604
rect 16028 34552 16080 34604
rect 17316 34595 17368 34604
rect 17316 34561 17325 34595
rect 17325 34561 17359 34595
rect 17359 34561 17368 34595
rect 18236 34595 18288 34604
rect 17316 34552 17368 34561
rect 18236 34561 18245 34595
rect 18245 34561 18279 34595
rect 18279 34561 18288 34595
rect 18236 34552 18288 34561
rect 18604 34552 18656 34604
rect 21548 34688 21600 34740
rect 23756 34688 23808 34740
rect 31116 34688 31168 34740
rect 19064 34620 19116 34672
rect 21180 34620 21232 34672
rect 21640 34620 21692 34672
rect 19248 34552 19300 34604
rect 8392 34416 8444 34468
rect 9772 34416 9824 34468
rect 10968 34416 11020 34468
rect 9128 34348 9180 34400
rect 10140 34391 10192 34400
rect 10140 34357 10149 34391
rect 10149 34357 10183 34391
rect 10183 34357 10192 34391
rect 10140 34348 10192 34357
rect 10232 34348 10284 34400
rect 11704 34391 11756 34400
rect 11704 34357 11713 34391
rect 11713 34357 11747 34391
rect 11747 34357 11756 34391
rect 11704 34348 11756 34357
rect 12072 34348 12124 34400
rect 14280 34527 14332 34536
rect 14280 34493 14289 34527
rect 14289 34493 14323 34527
rect 14323 34493 14332 34527
rect 14280 34484 14332 34493
rect 15660 34484 15712 34536
rect 19616 34527 19668 34536
rect 17684 34416 17736 34468
rect 19616 34493 19625 34527
rect 19625 34493 19659 34527
rect 19659 34493 19668 34527
rect 19616 34484 19668 34493
rect 21456 34552 21508 34604
rect 19248 34416 19300 34468
rect 21088 34484 21140 34536
rect 21824 34484 21876 34536
rect 22192 34595 22244 34604
rect 22192 34561 22201 34595
rect 22201 34561 22235 34595
rect 22235 34561 22244 34595
rect 22192 34552 22244 34561
rect 22560 34595 22612 34604
rect 22560 34561 22569 34595
rect 22569 34561 22603 34595
rect 22603 34561 22612 34595
rect 22560 34552 22612 34561
rect 22836 34552 22888 34604
rect 25688 34620 25740 34672
rect 24952 34552 25004 34604
rect 28264 34552 28316 34604
rect 28908 34552 28960 34604
rect 23848 34527 23900 34536
rect 23848 34493 23857 34527
rect 23857 34493 23891 34527
rect 23891 34493 23900 34527
rect 23848 34484 23900 34493
rect 28356 34527 28408 34536
rect 28356 34493 28365 34527
rect 28365 34493 28399 34527
rect 28399 34493 28408 34527
rect 28356 34484 28408 34493
rect 14740 34348 14792 34400
rect 17408 34348 17460 34400
rect 18144 34348 18196 34400
rect 19064 34348 19116 34400
rect 21824 34391 21876 34400
rect 21824 34357 21833 34391
rect 21833 34357 21867 34391
rect 21867 34357 21876 34391
rect 21824 34348 21876 34357
rect 29000 34391 29052 34400
rect 29000 34357 29009 34391
rect 29009 34357 29043 34391
rect 29043 34357 29052 34391
rect 29000 34348 29052 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 4068 34144 4120 34196
rect 6552 34144 6604 34196
rect 7288 34144 7340 34196
rect 8760 34187 8812 34196
rect 8760 34153 8769 34187
rect 8769 34153 8803 34187
rect 8803 34153 8812 34187
rect 8760 34144 8812 34153
rect 9036 34144 9088 34196
rect 9680 34144 9732 34196
rect 10600 34144 10652 34196
rect 6736 34008 6788 34060
rect 8208 34008 8260 34060
rect 8944 34076 8996 34128
rect 4160 33940 4212 33992
rect 4620 33940 4672 33992
rect 5632 33940 5684 33992
rect 8484 33983 8536 33992
rect 8484 33949 8493 33983
rect 8493 33949 8527 33983
rect 8527 33949 8536 33983
rect 8484 33940 8536 33949
rect 8760 33940 8812 33992
rect 9128 33983 9180 33992
rect 9128 33949 9137 33983
rect 9137 33949 9171 33983
rect 9171 33949 9180 33983
rect 9128 33940 9180 33949
rect 9680 33983 9732 33992
rect 9680 33949 9689 33983
rect 9689 33949 9723 33983
rect 9723 33949 9732 33983
rect 9680 33940 9732 33949
rect 1676 33872 1728 33924
rect 2320 33872 2372 33924
rect 8668 33872 8720 33924
rect 9772 33847 9824 33856
rect 9772 33813 9781 33847
rect 9781 33813 9815 33847
rect 9815 33813 9824 33847
rect 9772 33804 9824 33813
rect 10048 33872 10100 33924
rect 10324 33940 10376 33992
rect 10968 34187 11020 34196
rect 10968 34153 10977 34187
rect 10977 34153 11011 34187
rect 11011 34153 11020 34187
rect 10968 34144 11020 34153
rect 12256 34144 12308 34196
rect 12440 34144 12492 34196
rect 12072 34008 12124 34060
rect 11152 33983 11204 33992
rect 11152 33949 11161 33983
rect 11161 33949 11195 33983
rect 11195 33949 11204 33983
rect 11152 33940 11204 33949
rect 11336 33983 11388 33992
rect 11336 33949 11345 33983
rect 11345 33949 11379 33983
rect 11379 33949 11388 33983
rect 11336 33940 11388 33949
rect 11704 33940 11756 33992
rect 12348 34051 12400 34060
rect 12348 34017 12357 34051
rect 12357 34017 12391 34051
rect 12391 34017 12400 34051
rect 12348 34008 12400 34017
rect 18328 34144 18380 34196
rect 18604 34144 18656 34196
rect 23848 34144 23900 34196
rect 28356 34144 28408 34196
rect 16580 34076 16632 34128
rect 13820 34008 13872 34060
rect 14740 34051 14792 34060
rect 14740 34017 14749 34051
rect 14749 34017 14783 34051
rect 14783 34017 14792 34051
rect 14740 34008 14792 34017
rect 17132 34008 17184 34060
rect 18236 34076 18288 34128
rect 21548 34076 21600 34128
rect 13084 33983 13136 33992
rect 13084 33949 13093 33983
rect 13093 33949 13127 33983
rect 13127 33949 13136 33983
rect 13084 33940 13136 33949
rect 17408 33983 17460 33992
rect 17408 33949 17417 33983
rect 17417 33949 17451 33983
rect 17451 33949 17460 33983
rect 17408 33940 17460 33949
rect 15016 33872 15068 33924
rect 18144 33983 18196 33992
rect 18144 33949 18153 33983
rect 18153 33949 18187 33983
rect 18187 33949 18196 33983
rect 18144 33940 18196 33949
rect 18880 34051 18932 34060
rect 18880 34017 18889 34051
rect 18889 34017 18923 34051
rect 18923 34017 18932 34051
rect 18880 34008 18932 34017
rect 20168 34008 20220 34060
rect 20904 34008 20956 34060
rect 25136 34008 25188 34060
rect 25872 34008 25924 34060
rect 28908 34008 28960 34060
rect 29920 34008 29972 34060
rect 18512 33940 18564 33992
rect 21824 33940 21876 33992
rect 11704 33804 11756 33856
rect 16304 33804 16356 33856
rect 17592 33847 17644 33856
rect 17592 33813 17601 33847
rect 17601 33813 17635 33847
rect 17635 33813 17644 33847
rect 17592 33804 17644 33813
rect 18328 33804 18380 33856
rect 21732 33872 21784 33924
rect 25688 33940 25740 33992
rect 30196 33940 30248 33992
rect 32036 33940 32088 33992
rect 28356 33872 28408 33924
rect 29736 33872 29788 33924
rect 30472 33872 30524 33924
rect 32680 33872 32732 33924
rect 31392 33804 31444 33856
rect 32496 33804 32548 33856
rect 34060 33804 34112 33856
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 2228 33600 2280 33652
rect 4160 33600 4212 33652
rect 5540 33600 5592 33652
rect 9680 33600 9732 33652
rect 1492 33532 1544 33584
rect 2228 33507 2280 33516
rect 2228 33473 2237 33507
rect 2237 33473 2271 33507
rect 2271 33473 2280 33507
rect 2228 33464 2280 33473
rect 6644 33532 6696 33584
rect 1676 33396 1728 33448
rect 2872 33328 2924 33380
rect 5632 33464 5684 33516
rect 6000 33507 6052 33516
rect 6000 33473 6009 33507
rect 6009 33473 6043 33507
rect 6043 33473 6052 33507
rect 6000 33464 6052 33473
rect 6368 33464 6420 33516
rect 7196 33507 7248 33516
rect 7196 33473 7205 33507
rect 7205 33473 7239 33507
rect 7239 33473 7248 33507
rect 7196 33464 7248 33473
rect 7288 33464 7340 33516
rect 7840 33507 7892 33516
rect 7840 33473 7849 33507
rect 7849 33473 7883 33507
rect 7883 33473 7892 33507
rect 7840 33464 7892 33473
rect 10324 33600 10376 33652
rect 14280 33600 14332 33652
rect 14740 33600 14792 33652
rect 8392 33464 8444 33516
rect 8484 33507 8536 33516
rect 8484 33473 8493 33507
rect 8493 33473 8527 33507
rect 8527 33473 8536 33507
rect 8484 33464 8536 33473
rect 9036 33464 9088 33516
rect 9588 33507 9640 33516
rect 9588 33473 9597 33507
rect 9597 33473 9631 33507
rect 9631 33473 9640 33507
rect 9588 33464 9640 33473
rect 4160 33396 4212 33448
rect 5816 33439 5868 33448
rect 5816 33405 5825 33439
rect 5825 33405 5859 33439
rect 5859 33405 5868 33439
rect 5816 33396 5868 33405
rect 6092 33328 6144 33380
rect 6828 33439 6880 33448
rect 6828 33405 6837 33439
rect 6837 33405 6871 33439
rect 6871 33405 6880 33439
rect 6828 33396 6880 33405
rect 7104 33396 7156 33448
rect 7472 33396 7524 33448
rect 8668 33396 8720 33448
rect 8944 33396 8996 33448
rect 10048 33507 10100 33516
rect 10048 33473 10057 33507
rect 10057 33473 10091 33507
rect 10091 33473 10100 33507
rect 10048 33464 10100 33473
rect 10232 33507 10284 33516
rect 10232 33473 10241 33507
rect 10241 33473 10275 33507
rect 10275 33473 10284 33507
rect 10232 33464 10284 33473
rect 15292 33575 15344 33584
rect 15292 33541 15301 33575
rect 15301 33541 15335 33575
rect 15335 33541 15344 33575
rect 15292 33532 15344 33541
rect 15660 33643 15712 33652
rect 15660 33609 15669 33643
rect 15669 33609 15703 33643
rect 15703 33609 15712 33643
rect 15660 33600 15712 33609
rect 16396 33600 16448 33652
rect 16672 33600 16724 33652
rect 18144 33600 18196 33652
rect 18236 33600 18288 33652
rect 18604 33600 18656 33652
rect 20168 33643 20220 33652
rect 20168 33609 20177 33643
rect 20177 33609 20211 33643
rect 20211 33609 20220 33643
rect 20168 33600 20220 33609
rect 29736 33600 29788 33652
rect 30196 33643 30248 33652
rect 30196 33609 30205 33643
rect 30205 33609 30239 33643
rect 30239 33609 30248 33643
rect 30196 33600 30248 33609
rect 32680 33643 32732 33652
rect 32680 33609 32689 33643
rect 32689 33609 32723 33643
rect 32723 33609 32732 33643
rect 32680 33600 32732 33609
rect 16120 33532 16172 33584
rect 17132 33532 17184 33584
rect 7012 33328 7064 33380
rect 7380 33328 7432 33380
rect 9772 33328 9824 33380
rect 10140 33396 10192 33448
rect 13084 33464 13136 33516
rect 11152 33328 11204 33380
rect 3608 33260 3660 33312
rect 5172 33303 5224 33312
rect 5172 33269 5181 33303
rect 5181 33269 5215 33303
rect 5215 33269 5224 33303
rect 5172 33260 5224 33269
rect 7656 33303 7708 33312
rect 7656 33269 7665 33303
rect 7665 33269 7699 33303
rect 7699 33269 7708 33303
rect 7656 33260 7708 33269
rect 9036 33260 9088 33312
rect 14740 33439 14792 33448
rect 14740 33405 14749 33439
rect 14749 33405 14783 33439
rect 14783 33405 14792 33439
rect 14740 33396 14792 33405
rect 16304 33396 16356 33448
rect 17224 33396 17276 33448
rect 17684 33439 17736 33448
rect 17684 33405 17693 33439
rect 17693 33405 17727 33439
rect 17727 33405 17736 33439
rect 17684 33396 17736 33405
rect 17960 33439 18012 33448
rect 17960 33405 17969 33439
rect 17969 33405 18003 33439
rect 18003 33405 18012 33439
rect 17960 33396 18012 33405
rect 18512 33396 18564 33448
rect 19248 33532 19300 33584
rect 28356 33532 28408 33584
rect 29000 33532 29052 33584
rect 18144 33260 18196 33312
rect 28908 33464 28960 33516
rect 29552 33507 29604 33516
rect 29552 33473 29561 33507
rect 29561 33473 29595 33507
rect 29595 33473 29604 33507
rect 29552 33464 29604 33473
rect 29644 33464 29696 33516
rect 19708 33439 19760 33448
rect 19708 33405 19717 33439
rect 19717 33405 19751 33439
rect 19751 33405 19760 33439
rect 19708 33396 19760 33405
rect 28448 33439 28500 33448
rect 28448 33405 28457 33439
rect 28457 33405 28491 33439
rect 28491 33405 28500 33439
rect 28448 33396 28500 33405
rect 19892 33260 19944 33312
rect 24400 33260 24452 33312
rect 28080 33260 28132 33312
rect 29000 33396 29052 33448
rect 29092 33328 29144 33380
rect 30104 33396 30156 33448
rect 29460 33303 29512 33312
rect 29460 33269 29469 33303
rect 29469 33269 29503 33303
rect 29503 33269 29512 33303
rect 29460 33260 29512 33269
rect 31392 33507 31444 33516
rect 31392 33473 31401 33507
rect 31401 33473 31435 33507
rect 31435 33473 31444 33507
rect 31392 33464 31444 33473
rect 31944 33507 31996 33516
rect 31944 33473 31953 33507
rect 31953 33473 31987 33507
rect 31987 33473 31996 33507
rect 31944 33464 31996 33473
rect 32956 33464 33008 33516
rect 34060 33507 34112 33516
rect 34060 33473 34069 33507
rect 34069 33473 34103 33507
rect 34103 33473 34112 33507
rect 34060 33464 34112 33473
rect 34244 33507 34296 33516
rect 34244 33473 34253 33507
rect 34253 33473 34287 33507
rect 34287 33473 34296 33507
rect 34244 33464 34296 33473
rect 30748 33328 30800 33380
rect 38752 33396 38804 33448
rect 31024 33260 31076 33312
rect 33140 33260 33192 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 3792 33056 3844 33108
rect 5632 33099 5684 33108
rect 5632 33065 5641 33099
rect 5641 33065 5675 33099
rect 5675 33065 5684 33099
rect 5632 33056 5684 33065
rect 8392 33056 8444 33108
rect 9220 33056 9272 33108
rect 9588 33056 9640 33108
rect 15292 33056 15344 33108
rect 12440 32988 12492 33040
rect 15844 32988 15896 33040
rect 2872 32920 2924 32972
rect 5172 32920 5224 32972
rect 6552 32920 6604 32972
rect 6920 32963 6972 32972
rect 6920 32929 6929 32963
rect 6929 32929 6963 32963
rect 6963 32929 6972 32963
rect 6920 32920 6972 32929
rect 7656 32920 7708 32972
rect 8392 32920 8444 32972
rect 8668 32920 8720 32972
rect 3884 32895 3936 32904
rect 3884 32861 3893 32895
rect 3893 32861 3927 32895
rect 3927 32861 3936 32895
rect 3884 32852 3936 32861
rect 10600 32852 10652 32904
rect 12532 32852 12584 32904
rect 15568 32895 15620 32904
rect 15568 32861 15577 32895
rect 15577 32861 15611 32895
rect 15611 32861 15620 32895
rect 15568 32852 15620 32861
rect 17960 33056 18012 33108
rect 28448 33056 28500 33108
rect 29552 33056 29604 33108
rect 29736 33056 29788 33108
rect 22560 32988 22612 33040
rect 33232 33056 33284 33108
rect 34244 33056 34296 33108
rect 34336 32988 34388 33040
rect 16120 32852 16172 32904
rect 16488 32895 16540 32904
rect 16488 32861 16497 32895
rect 16497 32861 16531 32895
rect 16531 32861 16540 32895
rect 16488 32852 16540 32861
rect 17592 32895 17644 32904
rect 17592 32861 17601 32895
rect 17601 32861 17635 32895
rect 17635 32861 17644 32895
rect 17592 32852 17644 32861
rect 18328 32920 18380 32972
rect 1492 32827 1544 32836
rect 1492 32793 1501 32827
rect 1501 32793 1535 32827
rect 1535 32793 1544 32827
rect 1492 32784 1544 32793
rect 2780 32784 2832 32836
rect 5540 32784 5592 32836
rect 6276 32784 6328 32836
rect 7288 32784 7340 32836
rect 5816 32716 5868 32768
rect 6552 32759 6604 32768
rect 6552 32725 6561 32759
rect 6561 32725 6595 32759
rect 6595 32725 6604 32759
rect 6552 32716 6604 32725
rect 11060 32716 11112 32768
rect 16028 32716 16080 32768
rect 16672 32784 16724 32836
rect 16396 32716 16448 32768
rect 18144 32895 18196 32904
rect 18144 32861 18153 32895
rect 18153 32861 18187 32895
rect 18187 32861 18196 32895
rect 18144 32852 18196 32861
rect 18236 32852 18288 32904
rect 18604 32784 18656 32836
rect 23664 32827 23716 32836
rect 23664 32793 23673 32827
rect 23673 32793 23707 32827
rect 23707 32793 23716 32827
rect 23664 32784 23716 32793
rect 24124 32852 24176 32904
rect 24676 32852 24728 32904
rect 26792 32920 26844 32972
rect 25780 32852 25832 32904
rect 26148 32895 26200 32904
rect 26148 32861 26161 32895
rect 26161 32861 26200 32895
rect 26148 32852 26200 32861
rect 28908 32920 28960 32972
rect 29460 32920 29512 32972
rect 29920 32963 29972 32972
rect 29920 32929 29929 32963
rect 29929 32929 29963 32963
rect 29963 32929 29972 32963
rect 29920 32920 29972 32929
rect 30196 32920 30248 32972
rect 32036 32920 32088 32972
rect 28816 32895 28868 32904
rect 28816 32861 28825 32895
rect 28825 32861 28859 32895
rect 28859 32861 28868 32895
rect 28816 32852 28868 32861
rect 29092 32852 29144 32904
rect 29552 32895 29604 32904
rect 29552 32861 29561 32895
rect 29561 32861 29595 32895
rect 29595 32861 29604 32895
rect 29552 32852 29604 32861
rect 23756 32759 23808 32768
rect 23756 32725 23771 32759
rect 23771 32725 23805 32759
rect 23805 32725 23808 32759
rect 23756 32716 23808 32725
rect 25044 32716 25096 32768
rect 25596 32716 25648 32768
rect 26424 32716 26476 32768
rect 28816 32716 28868 32768
rect 32220 32852 32272 32904
rect 33692 32895 33744 32904
rect 33692 32861 33701 32895
rect 33701 32861 33735 32895
rect 33735 32861 33744 32895
rect 33692 32852 33744 32861
rect 30472 32784 30524 32836
rect 30932 32784 30984 32836
rect 32496 32784 32548 32836
rect 37280 32852 37332 32904
rect 30288 32716 30340 32768
rect 31668 32759 31720 32768
rect 31668 32725 31677 32759
rect 31677 32725 31711 32759
rect 31711 32725 31720 32759
rect 31668 32716 31720 32725
rect 32404 32716 32456 32768
rect 35992 32784 36044 32836
rect 34428 32759 34480 32768
rect 34428 32725 34437 32759
rect 34437 32725 34471 32759
rect 34471 32725 34480 32759
rect 34428 32716 34480 32725
rect 36452 32827 36504 32836
rect 36452 32793 36461 32827
rect 36461 32793 36495 32827
rect 36495 32793 36504 32827
rect 36452 32784 36504 32793
rect 39672 32716 39724 32768
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 5540 32512 5592 32564
rect 6828 32512 6880 32564
rect 7380 32555 7432 32564
rect 7380 32521 7389 32555
rect 7389 32521 7423 32555
rect 7423 32521 7432 32555
rect 7380 32512 7432 32521
rect 7840 32512 7892 32564
rect 12532 32512 12584 32564
rect 15844 32512 15896 32564
rect 18144 32512 18196 32564
rect 1676 32444 1728 32496
rect 2596 32444 2648 32496
rect 3608 32487 3660 32496
rect 3608 32453 3617 32487
rect 3617 32453 3651 32487
rect 3651 32453 3660 32487
rect 3608 32444 3660 32453
rect 6552 32487 6604 32496
rect 6552 32453 6563 32487
rect 6563 32453 6604 32487
rect 6552 32444 6604 32453
rect 6644 32444 6696 32496
rect 6920 32444 6972 32496
rect 8852 32444 8904 32496
rect 3884 32351 3936 32360
rect 3884 32317 3893 32351
rect 3893 32317 3927 32351
rect 3927 32317 3936 32351
rect 3884 32308 3936 32317
rect 5632 32376 5684 32428
rect 6184 32376 6236 32428
rect 7196 32376 7248 32428
rect 7472 32419 7524 32428
rect 7472 32385 7482 32419
rect 7482 32385 7524 32419
rect 7472 32376 7524 32385
rect 8576 32419 8628 32428
rect 8576 32385 8585 32419
rect 8585 32385 8619 32419
rect 8619 32385 8628 32419
rect 8576 32376 8628 32385
rect 11612 32376 11664 32428
rect 13084 32419 13136 32428
rect 5540 32308 5592 32360
rect 5816 32351 5868 32360
rect 5816 32317 5825 32351
rect 5825 32317 5859 32351
rect 5859 32317 5868 32351
rect 5816 32308 5868 32317
rect 6920 32351 6972 32360
rect 6920 32317 6929 32351
rect 6929 32317 6963 32351
rect 6963 32317 6972 32351
rect 6920 32308 6972 32317
rect 9220 32308 9272 32360
rect 10968 32308 11020 32360
rect 11888 32308 11940 32360
rect 13084 32385 13093 32419
rect 13093 32385 13127 32419
rect 13127 32385 13136 32419
rect 13084 32376 13136 32385
rect 13912 32376 13964 32428
rect 14188 32419 14240 32428
rect 14188 32385 14197 32419
rect 14197 32385 14231 32419
rect 14231 32385 14240 32419
rect 14188 32376 14240 32385
rect 12532 32351 12584 32360
rect 12532 32317 12541 32351
rect 12541 32317 12575 32351
rect 12575 32317 12584 32351
rect 12532 32308 12584 32317
rect 12624 32308 12676 32360
rect 13820 32308 13872 32360
rect 5908 32240 5960 32292
rect 6368 32283 6420 32292
rect 6368 32249 6377 32283
rect 6377 32249 6411 32283
rect 6411 32249 6420 32283
rect 6368 32240 6420 32249
rect 6000 32172 6052 32224
rect 6276 32172 6328 32224
rect 6552 32215 6604 32224
rect 6552 32181 6561 32215
rect 6561 32181 6595 32215
rect 6595 32181 6604 32215
rect 6552 32172 6604 32181
rect 12072 32240 12124 32292
rect 12440 32172 12492 32224
rect 12992 32240 13044 32292
rect 14648 32376 14700 32428
rect 16120 32444 16172 32496
rect 18236 32444 18288 32496
rect 20352 32444 20404 32496
rect 21456 32444 21508 32496
rect 17040 32376 17092 32428
rect 20904 32376 20956 32428
rect 22192 32376 22244 32428
rect 14740 32351 14792 32360
rect 14740 32317 14749 32351
rect 14749 32317 14783 32351
rect 14783 32317 14792 32351
rect 14740 32308 14792 32317
rect 15384 32308 15436 32360
rect 16212 32308 16264 32360
rect 19432 32308 19484 32360
rect 20352 32351 20404 32360
rect 20352 32317 20361 32351
rect 20361 32317 20395 32351
rect 20395 32317 20404 32351
rect 20352 32308 20404 32317
rect 15200 32240 15252 32292
rect 14556 32172 14608 32224
rect 20352 32172 20404 32224
rect 21824 32215 21876 32224
rect 21824 32181 21833 32215
rect 21833 32181 21867 32215
rect 21867 32181 21876 32215
rect 21824 32172 21876 32181
rect 22744 32419 22796 32428
rect 22744 32385 22753 32419
rect 22753 32385 22787 32419
rect 22787 32385 22796 32419
rect 22744 32376 22796 32385
rect 22652 32308 22704 32360
rect 23020 32376 23072 32428
rect 23296 32376 23348 32428
rect 23388 32419 23440 32428
rect 23388 32385 23397 32419
rect 23397 32385 23431 32419
rect 23431 32385 23440 32419
rect 23388 32376 23440 32385
rect 23756 32376 23808 32428
rect 25688 32512 25740 32564
rect 25780 32512 25832 32564
rect 24676 32487 24728 32496
rect 24676 32453 24685 32487
rect 24685 32453 24719 32487
rect 24719 32453 24728 32487
rect 24676 32444 24728 32453
rect 25136 32444 25188 32496
rect 24860 32419 24912 32428
rect 24860 32385 24869 32419
rect 24869 32385 24903 32419
rect 24903 32385 24912 32419
rect 24860 32376 24912 32385
rect 24952 32419 25004 32428
rect 24952 32385 24961 32419
rect 24961 32385 24995 32419
rect 24995 32385 25004 32419
rect 24952 32376 25004 32385
rect 25044 32419 25096 32428
rect 25044 32385 25058 32419
rect 25058 32385 25092 32419
rect 25092 32385 25096 32419
rect 25044 32376 25096 32385
rect 25320 32419 25372 32428
rect 25320 32385 25329 32419
rect 25329 32385 25363 32419
rect 25363 32385 25372 32419
rect 25320 32376 25372 32385
rect 25412 32419 25464 32428
rect 25412 32385 25421 32419
rect 25421 32385 25455 32419
rect 25455 32385 25464 32419
rect 25412 32376 25464 32385
rect 25596 32419 25648 32428
rect 25596 32385 25605 32419
rect 25605 32385 25639 32419
rect 25639 32385 25648 32419
rect 25596 32376 25648 32385
rect 26424 32487 26476 32496
rect 26424 32453 26433 32487
rect 26433 32453 26467 32487
rect 26467 32453 26476 32487
rect 26424 32444 26476 32453
rect 28080 32444 28132 32496
rect 28908 32512 28960 32564
rect 29000 32512 29052 32564
rect 29736 32512 29788 32564
rect 29920 32555 29972 32564
rect 29920 32521 29929 32555
rect 29929 32521 29963 32555
rect 29963 32521 29972 32555
rect 29920 32512 29972 32521
rect 31944 32512 31996 32564
rect 23848 32308 23900 32360
rect 24492 32351 24544 32360
rect 24492 32317 24501 32351
rect 24501 32317 24535 32351
rect 24535 32317 24544 32351
rect 24492 32308 24544 32317
rect 26056 32419 26108 32428
rect 26056 32385 26065 32419
rect 26065 32385 26099 32419
rect 26099 32385 26108 32419
rect 26056 32376 26108 32385
rect 26332 32419 26384 32428
rect 26332 32385 26341 32419
rect 26341 32385 26375 32419
rect 26375 32385 26384 32419
rect 26332 32376 26384 32385
rect 27896 32376 27948 32428
rect 26700 32308 26752 32360
rect 28448 32351 28500 32360
rect 28448 32317 28457 32351
rect 28457 32317 28491 32351
rect 28491 32317 28500 32351
rect 28448 32308 28500 32317
rect 28816 32419 28868 32428
rect 28816 32385 28825 32419
rect 28825 32385 28859 32419
rect 28859 32385 28868 32419
rect 28816 32376 28868 32385
rect 30196 32444 30248 32496
rect 31116 32487 31168 32496
rect 31116 32453 31125 32487
rect 31125 32453 31159 32487
rect 31159 32453 31168 32487
rect 31116 32444 31168 32453
rect 33048 32444 33100 32496
rect 33692 32487 33744 32496
rect 33692 32453 33701 32487
rect 33701 32453 33735 32487
rect 33735 32453 33744 32487
rect 33692 32444 33744 32453
rect 34336 32512 34388 32564
rect 36452 32512 36504 32564
rect 34612 32444 34664 32496
rect 29092 32376 29144 32428
rect 31392 32376 31444 32428
rect 31484 32376 31536 32428
rect 29368 32308 29420 32360
rect 29736 32308 29788 32360
rect 32404 32376 32456 32428
rect 33968 32419 34020 32428
rect 33968 32385 33977 32419
rect 33977 32385 34011 32419
rect 34011 32385 34020 32419
rect 33968 32376 34020 32385
rect 34152 32419 34204 32428
rect 34152 32385 34161 32419
rect 34161 32385 34195 32419
rect 34195 32385 34204 32419
rect 34152 32376 34204 32385
rect 37280 32376 37332 32428
rect 38200 32376 38252 32428
rect 22744 32172 22796 32224
rect 28540 32240 28592 32292
rect 30012 32240 30064 32292
rect 30104 32283 30156 32292
rect 30104 32249 30113 32283
rect 30113 32249 30147 32283
rect 30147 32249 30156 32283
rect 30104 32240 30156 32249
rect 24216 32172 24268 32224
rect 25320 32172 25372 32224
rect 26148 32172 26200 32224
rect 28080 32172 28132 32224
rect 31668 32240 31720 32292
rect 34428 32308 34480 32360
rect 35992 32308 36044 32360
rect 36084 32351 36136 32360
rect 36084 32317 36093 32351
rect 36093 32317 36127 32351
rect 36127 32317 36136 32351
rect 36084 32308 36136 32317
rect 37464 32351 37516 32360
rect 37464 32317 37473 32351
rect 37473 32317 37507 32351
rect 37507 32317 37516 32351
rect 37464 32308 37516 32317
rect 37556 32351 37608 32360
rect 37556 32317 37565 32351
rect 37565 32317 37599 32351
rect 37599 32317 37608 32351
rect 37556 32308 37608 32317
rect 37372 32240 37424 32292
rect 37832 32308 37884 32360
rect 31852 32172 31904 32224
rect 34796 32172 34848 32224
rect 38016 32172 38068 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2596 31968 2648 32020
rect 5724 31968 5776 32020
rect 6276 31968 6328 32020
rect 7380 31968 7432 32020
rect 8668 31968 8720 32020
rect 9036 32011 9088 32020
rect 9036 31977 9045 32011
rect 9045 31977 9079 32011
rect 9079 31977 9088 32011
rect 9036 31968 9088 31977
rect 10968 32011 11020 32020
rect 10968 31977 10977 32011
rect 10977 31977 11011 32011
rect 11011 31977 11020 32011
rect 10968 31968 11020 31977
rect 11060 32011 11112 32020
rect 11060 31977 11069 32011
rect 11069 31977 11103 32011
rect 11103 31977 11112 32011
rect 11060 31968 11112 31977
rect 11704 31968 11756 32020
rect 5540 31900 5592 31952
rect 6644 31900 6696 31952
rect 5816 31832 5868 31884
rect 6092 31832 6144 31884
rect 8024 31875 8076 31884
rect 8024 31841 8033 31875
rect 8033 31841 8067 31875
rect 8067 31841 8076 31875
rect 8024 31832 8076 31841
rect 3792 31764 3844 31816
rect 5908 31764 5960 31816
rect 5264 31696 5316 31748
rect 7840 31696 7892 31748
rect 11888 31832 11940 31884
rect 12532 31900 12584 31952
rect 12256 31832 12308 31884
rect 11244 31764 11296 31816
rect 12164 31807 12216 31816
rect 12164 31773 12173 31807
rect 12173 31773 12207 31807
rect 12207 31773 12216 31807
rect 12164 31764 12216 31773
rect 12716 31764 12768 31816
rect 13728 31807 13780 31816
rect 13728 31773 13737 31807
rect 13737 31773 13771 31807
rect 13771 31773 13780 31807
rect 13728 31764 13780 31773
rect 8208 31696 8260 31748
rect 8300 31628 8352 31680
rect 8760 31739 8812 31748
rect 8760 31705 8769 31739
rect 8769 31705 8803 31739
rect 8803 31705 8812 31739
rect 8760 31696 8812 31705
rect 8944 31696 8996 31748
rect 11152 31696 11204 31748
rect 11428 31739 11480 31748
rect 11428 31705 11437 31739
rect 11437 31705 11471 31739
rect 11471 31705 11480 31739
rect 13912 31807 13964 31816
rect 13912 31773 13921 31807
rect 13921 31773 13955 31807
rect 13955 31773 13964 31807
rect 13912 31764 13964 31773
rect 14556 31968 14608 32020
rect 14924 31968 14976 32020
rect 17224 31968 17276 32020
rect 14740 31875 14792 31884
rect 14740 31841 14749 31875
rect 14749 31841 14783 31875
rect 14783 31841 14792 31875
rect 14740 31832 14792 31841
rect 16120 31875 16172 31884
rect 16120 31841 16129 31875
rect 16129 31841 16163 31875
rect 16163 31841 16172 31875
rect 16120 31832 16172 31841
rect 17224 31875 17276 31884
rect 17224 31841 17233 31875
rect 17233 31841 17267 31875
rect 17267 31841 17276 31875
rect 17224 31832 17276 31841
rect 18052 31832 18104 31884
rect 21088 31968 21140 32020
rect 22560 32011 22612 32020
rect 22560 31977 22569 32011
rect 22569 31977 22603 32011
rect 22603 31977 22612 32011
rect 22560 31968 22612 31977
rect 23020 31968 23072 32020
rect 25320 31968 25372 32020
rect 26608 32011 26660 32020
rect 20628 31832 20680 31884
rect 15292 31807 15344 31816
rect 15292 31773 15301 31807
rect 15301 31773 15335 31807
rect 15335 31773 15344 31807
rect 15292 31764 15344 31773
rect 15476 31764 15528 31816
rect 16304 31807 16356 31816
rect 16304 31773 16313 31807
rect 16313 31773 16347 31807
rect 16347 31773 16356 31807
rect 16304 31764 16356 31773
rect 16396 31807 16448 31816
rect 16396 31773 16405 31807
rect 16405 31773 16439 31807
rect 16439 31773 16448 31807
rect 16396 31764 16448 31773
rect 11428 31696 11480 31705
rect 16764 31696 16816 31748
rect 9036 31628 9088 31680
rect 10508 31671 10560 31680
rect 10508 31637 10517 31671
rect 10517 31637 10551 31671
rect 10551 31637 10560 31671
rect 10508 31628 10560 31637
rect 11888 31628 11940 31680
rect 12992 31628 13044 31680
rect 13636 31628 13688 31680
rect 17960 31696 18012 31748
rect 18512 31628 18564 31680
rect 19248 31696 19300 31748
rect 19616 31739 19668 31748
rect 19616 31705 19625 31739
rect 19625 31705 19659 31739
rect 19659 31705 19668 31739
rect 19616 31696 19668 31705
rect 22100 31832 22152 31884
rect 22192 31807 22244 31816
rect 22192 31773 22201 31807
rect 22201 31773 22235 31807
rect 22235 31773 22244 31807
rect 22192 31764 22244 31773
rect 21364 31696 21416 31748
rect 19064 31628 19116 31680
rect 21180 31671 21232 31680
rect 21180 31637 21189 31671
rect 21189 31637 21223 31671
rect 21223 31637 21232 31671
rect 21180 31628 21232 31637
rect 22192 31628 22244 31680
rect 22652 31832 22704 31884
rect 25780 31900 25832 31952
rect 23020 31807 23072 31816
rect 23020 31773 23029 31807
rect 23029 31773 23063 31807
rect 23063 31773 23072 31807
rect 23020 31764 23072 31773
rect 23756 31832 23808 31884
rect 24860 31832 24912 31884
rect 23848 31764 23900 31816
rect 25228 31807 25280 31816
rect 25228 31773 25237 31807
rect 25237 31773 25271 31807
rect 25271 31773 25280 31807
rect 25228 31764 25280 31773
rect 25596 31764 25648 31816
rect 25688 31807 25740 31816
rect 25688 31773 25697 31807
rect 25697 31773 25731 31807
rect 25731 31773 25740 31807
rect 25688 31764 25740 31773
rect 26608 31977 26617 32011
rect 26617 31977 26651 32011
rect 26651 31977 26660 32011
rect 26608 31968 26660 31977
rect 26424 31900 26476 31952
rect 22836 31628 22888 31680
rect 23204 31671 23256 31680
rect 23204 31637 23213 31671
rect 23213 31637 23247 31671
rect 23247 31637 23256 31671
rect 23204 31628 23256 31637
rect 23296 31628 23348 31680
rect 24124 31739 24176 31748
rect 24124 31705 24133 31739
rect 24133 31705 24167 31739
rect 24167 31705 24176 31739
rect 24124 31696 24176 31705
rect 24584 31696 24636 31748
rect 26148 31764 26200 31816
rect 27344 31832 27396 31884
rect 27252 31807 27304 31816
rect 27252 31773 27261 31807
rect 27261 31773 27295 31807
rect 27295 31773 27304 31807
rect 27896 31968 27948 32020
rect 27988 31900 28040 31952
rect 30472 31968 30524 32020
rect 31668 31968 31720 32020
rect 29000 31900 29052 31952
rect 31392 31900 31444 31952
rect 27252 31764 27304 31773
rect 29092 31832 29144 31884
rect 28080 31807 28132 31816
rect 28080 31773 28089 31807
rect 28089 31773 28123 31807
rect 28123 31773 28132 31807
rect 28080 31764 28132 31773
rect 28264 31807 28316 31816
rect 28264 31773 28272 31807
rect 28272 31773 28306 31807
rect 28306 31773 28316 31807
rect 28264 31764 28316 31773
rect 28540 31764 28592 31816
rect 28632 31807 28684 31816
rect 28632 31773 28641 31807
rect 28641 31773 28675 31807
rect 28675 31773 28684 31807
rect 28632 31764 28684 31773
rect 28816 31807 28868 31816
rect 28816 31773 28825 31807
rect 28825 31773 28859 31807
rect 28859 31773 28868 31807
rect 28816 31764 28868 31773
rect 24216 31628 24268 31680
rect 26148 31628 26200 31680
rect 27068 31671 27120 31680
rect 27068 31637 27077 31671
rect 27077 31637 27111 31671
rect 27111 31637 27120 31671
rect 27068 31628 27120 31637
rect 27344 31628 27396 31680
rect 29000 31764 29052 31816
rect 28080 31628 28132 31680
rect 28632 31628 28684 31680
rect 30012 31764 30064 31816
rect 31024 31764 31076 31816
rect 31576 31832 31628 31884
rect 32128 32011 32180 32020
rect 32128 31977 32137 32011
rect 32137 31977 32171 32011
rect 32171 31977 32180 32011
rect 32128 31968 32180 31977
rect 32220 32011 32272 32020
rect 32220 31977 32229 32011
rect 32229 31977 32263 32011
rect 32263 31977 32272 32011
rect 32220 31968 32272 31977
rect 32404 31968 32456 32020
rect 33140 31968 33192 32020
rect 34612 31968 34664 32020
rect 32496 31900 32548 31952
rect 32956 31900 33008 31952
rect 31392 31807 31444 31816
rect 31392 31773 31401 31807
rect 31401 31773 31435 31807
rect 31435 31773 31444 31807
rect 31392 31764 31444 31773
rect 30656 31739 30708 31748
rect 30656 31705 30665 31739
rect 30665 31705 30699 31739
rect 30699 31705 30708 31739
rect 30656 31696 30708 31705
rect 31576 31696 31628 31748
rect 31484 31628 31536 31680
rect 32220 31764 32272 31816
rect 36084 32011 36136 32020
rect 36084 31977 36093 32011
rect 36093 31977 36127 32011
rect 36127 31977 36136 32011
rect 36084 31968 36136 31977
rect 38016 31968 38068 32020
rect 32036 31696 32088 31748
rect 32956 31764 33008 31816
rect 33232 31807 33284 31816
rect 33232 31773 33241 31807
rect 33241 31773 33275 31807
rect 33275 31773 33284 31807
rect 33232 31764 33284 31773
rect 34796 31875 34848 31884
rect 34796 31841 34805 31875
rect 34805 31841 34839 31875
rect 34839 31841 34848 31875
rect 34796 31832 34848 31841
rect 34888 31832 34940 31884
rect 34152 31764 34204 31816
rect 36728 31900 36780 31952
rect 38660 31900 38712 31952
rect 35992 31832 36044 31884
rect 36176 31832 36228 31884
rect 32772 31696 32824 31748
rect 36728 31764 36780 31816
rect 38200 31764 38252 31816
rect 38292 31807 38344 31816
rect 38292 31773 38301 31807
rect 38301 31773 38335 31807
rect 38335 31773 38344 31807
rect 38292 31764 38344 31773
rect 36544 31696 36596 31748
rect 34244 31628 34296 31680
rect 35440 31628 35492 31680
rect 35992 31628 36044 31680
rect 38568 31807 38620 31816
rect 38568 31773 38577 31807
rect 38577 31773 38611 31807
rect 38611 31773 38620 31807
rect 38568 31764 38620 31773
rect 38660 31807 38712 31816
rect 38660 31773 38669 31807
rect 38669 31773 38703 31807
rect 38703 31773 38712 31807
rect 38660 31764 38712 31773
rect 38384 31696 38436 31748
rect 39488 31696 39540 31748
rect 38844 31671 38896 31680
rect 38844 31637 38853 31671
rect 38853 31637 38887 31671
rect 38887 31637 38896 31671
rect 38844 31628 38896 31637
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 2872 31424 2924 31476
rect 5264 31424 5316 31476
rect 2688 31356 2740 31408
rect 5724 31467 5776 31476
rect 5724 31433 5733 31467
rect 5733 31433 5767 31467
rect 5767 31433 5776 31467
rect 5724 31424 5776 31433
rect 7288 31424 7340 31476
rect 8392 31424 8444 31476
rect 10876 31424 10928 31476
rect 10968 31467 11020 31476
rect 10968 31433 10977 31467
rect 10977 31433 11011 31467
rect 11011 31433 11020 31467
rect 10968 31424 11020 31433
rect 11612 31424 11664 31476
rect 12716 31467 12768 31476
rect 12716 31433 12725 31467
rect 12725 31433 12759 31467
rect 12759 31433 12768 31467
rect 12716 31424 12768 31433
rect 13820 31424 13872 31476
rect 14188 31424 14240 31476
rect 16764 31467 16816 31476
rect 16764 31433 16773 31467
rect 16773 31433 16807 31467
rect 16807 31433 16816 31467
rect 16764 31424 16816 31433
rect 18052 31424 18104 31476
rect 19616 31424 19668 31476
rect 21180 31424 21232 31476
rect 21364 31467 21416 31476
rect 21364 31433 21373 31467
rect 21373 31433 21407 31467
rect 21407 31433 21416 31467
rect 21364 31424 21416 31433
rect 21824 31424 21876 31476
rect 5816 31356 5868 31408
rect 5448 31288 5500 31340
rect 8576 31356 8628 31408
rect 8944 31399 8996 31408
rect 8944 31365 8953 31399
rect 8953 31365 8987 31399
rect 8987 31365 8996 31399
rect 8944 31356 8996 31365
rect 7380 31288 7432 31340
rect 3240 31263 3292 31272
rect 3240 31229 3249 31263
rect 3249 31229 3283 31263
rect 3283 31229 3292 31263
rect 3240 31220 3292 31229
rect 4988 31263 5040 31272
rect 4988 31229 4997 31263
rect 4997 31229 5031 31263
rect 5031 31229 5040 31263
rect 4988 31220 5040 31229
rect 5540 31220 5592 31272
rect 5908 31220 5960 31272
rect 7748 31263 7800 31272
rect 7748 31229 7757 31263
rect 7757 31229 7791 31263
rect 7791 31229 7800 31263
rect 7748 31220 7800 31229
rect 7840 31220 7892 31272
rect 8576 31220 8628 31272
rect 9404 31263 9456 31272
rect 9404 31229 9413 31263
rect 9413 31229 9447 31263
rect 9447 31229 9456 31263
rect 9404 31220 9456 31229
rect 9956 31331 10008 31340
rect 9956 31297 9965 31331
rect 9965 31297 9999 31331
rect 9999 31297 10008 31331
rect 9956 31288 10008 31297
rect 10784 31288 10836 31340
rect 10876 31331 10928 31340
rect 10876 31297 10885 31331
rect 10885 31297 10919 31331
rect 10919 31297 10928 31331
rect 10876 31288 10928 31297
rect 11152 31356 11204 31408
rect 11336 31356 11388 31408
rect 11888 31356 11940 31408
rect 11704 31331 11756 31340
rect 8668 31152 8720 31204
rect 9864 31195 9916 31204
rect 9864 31161 9873 31195
rect 9873 31161 9907 31195
rect 9907 31161 9916 31195
rect 9864 31152 9916 31161
rect 10692 31263 10744 31272
rect 10692 31229 10701 31263
rect 10701 31229 10735 31263
rect 10735 31229 10744 31263
rect 10692 31220 10744 31229
rect 10968 31220 11020 31272
rect 11060 31220 11112 31272
rect 11704 31297 11710 31331
rect 11710 31297 11744 31331
rect 11744 31297 11756 31331
rect 11704 31288 11756 31297
rect 12072 31331 12124 31340
rect 12072 31297 12081 31331
rect 12081 31297 12115 31331
rect 12115 31297 12124 31331
rect 12072 31288 12124 31297
rect 12532 31356 12584 31408
rect 12900 31331 12952 31340
rect 12900 31297 12909 31331
rect 12909 31297 12943 31331
rect 12943 31297 12952 31331
rect 12900 31288 12952 31297
rect 12992 31331 13044 31340
rect 12992 31297 13001 31331
rect 13001 31297 13035 31331
rect 13035 31297 13044 31331
rect 12992 31288 13044 31297
rect 11336 31263 11388 31272
rect 11336 31229 11345 31263
rect 11345 31229 11379 31263
rect 11379 31229 11388 31263
rect 13636 31288 13688 31340
rect 13728 31331 13780 31340
rect 13728 31297 13737 31331
rect 13737 31297 13771 31331
rect 13771 31297 13780 31331
rect 13728 31288 13780 31297
rect 13912 31331 13964 31340
rect 13912 31297 13925 31331
rect 13925 31297 13964 31331
rect 13912 31288 13964 31297
rect 14188 31331 14240 31340
rect 14188 31297 14197 31331
rect 14197 31297 14231 31331
rect 14231 31297 14240 31331
rect 14188 31288 14240 31297
rect 14464 31288 14516 31340
rect 11336 31220 11388 31229
rect 14648 31220 14700 31272
rect 15016 31220 15068 31272
rect 15292 31356 15344 31408
rect 15476 31288 15528 31340
rect 16028 31288 16080 31340
rect 19156 31356 19208 31408
rect 19248 31356 19300 31408
rect 16948 31288 17000 31340
rect 17500 31331 17552 31340
rect 17500 31297 17509 31331
rect 17509 31297 17543 31331
rect 17543 31297 17552 31331
rect 17500 31288 17552 31297
rect 18236 31331 18288 31340
rect 18236 31297 18245 31331
rect 18245 31297 18279 31331
rect 18279 31297 18288 31331
rect 18236 31288 18288 31297
rect 18420 31288 18472 31340
rect 15384 31263 15436 31272
rect 15384 31229 15393 31263
rect 15393 31229 15427 31263
rect 15427 31229 15436 31263
rect 15384 31220 15436 31229
rect 15660 31220 15712 31272
rect 17224 31263 17276 31272
rect 17224 31229 17233 31263
rect 17233 31229 17267 31263
rect 17267 31229 17276 31263
rect 17224 31220 17276 31229
rect 16304 31152 16356 31204
rect 17868 31220 17920 31272
rect 19064 31220 19116 31272
rect 20352 31263 20404 31272
rect 20352 31229 20361 31263
rect 20361 31229 20395 31263
rect 20395 31229 20404 31263
rect 20352 31220 20404 31229
rect 20444 31220 20496 31272
rect 20996 31288 21048 31340
rect 22100 31356 22152 31408
rect 22928 31424 22980 31476
rect 23848 31424 23900 31476
rect 22928 31288 22980 31340
rect 23112 31331 23164 31340
rect 23112 31297 23121 31331
rect 23121 31297 23155 31331
rect 23155 31297 23164 31331
rect 23112 31288 23164 31297
rect 23296 31331 23348 31340
rect 23296 31297 23305 31331
rect 23305 31297 23339 31331
rect 23339 31297 23348 31331
rect 23296 31288 23348 31297
rect 23572 31288 23624 31340
rect 24952 31356 25004 31408
rect 22376 31220 22428 31272
rect 22560 31263 22612 31272
rect 22560 31229 22569 31263
rect 22569 31229 22603 31263
rect 22603 31229 22612 31263
rect 22560 31220 22612 31229
rect 23848 31263 23900 31272
rect 23848 31229 23857 31263
rect 23857 31229 23891 31263
rect 23891 31229 23900 31263
rect 23848 31220 23900 31229
rect 4896 31084 4948 31136
rect 7380 31084 7432 31136
rect 9588 31127 9640 31136
rect 9588 31093 9597 31127
rect 9597 31093 9631 31127
rect 9631 31093 9640 31127
rect 9588 31084 9640 31093
rect 9956 31084 10008 31136
rect 11244 31084 11296 31136
rect 11520 31127 11572 31136
rect 11520 31093 11529 31127
rect 11529 31093 11563 31127
rect 11563 31093 11572 31127
rect 11520 31084 11572 31093
rect 13912 31084 13964 31136
rect 16028 31084 16080 31136
rect 19524 31084 19576 31136
rect 20812 31084 20864 31136
rect 20904 31084 20956 31136
rect 21640 31084 21692 31136
rect 22192 31152 22244 31204
rect 23204 31152 23256 31204
rect 22376 31127 22428 31136
rect 22376 31093 22385 31127
rect 22385 31093 22419 31127
rect 22419 31093 22428 31127
rect 22376 31084 22428 31093
rect 23020 31084 23072 31136
rect 24308 31127 24360 31136
rect 24308 31093 24317 31127
rect 24317 31093 24351 31127
rect 24351 31093 24360 31127
rect 24308 31084 24360 31093
rect 24952 31263 25004 31272
rect 24952 31229 24961 31263
rect 24961 31229 24995 31263
rect 24995 31229 25004 31263
rect 24952 31220 25004 31229
rect 25780 31424 25832 31476
rect 26056 31424 26108 31476
rect 25412 31356 25464 31408
rect 28448 31424 28500 31476
rect 29644 31467 29696 31476
rect 29644 31433 29653 31467
rect 29653 31433 29687 31467
rect 29687 31433 29696 31467
rect 29644 31424 29696 31433
rect 25688 31288 25740 31340
rect 25964 31331 26016 31340
rect 25964 31297 25973 31331
rect 25973 31297 26007 31331
rect 26007 31297 26016 31331
rect 25964 31288 26016 31297
rect 28816 31356 28868 31408
rect 26516 31331 26568 31340
rect 26516 31297 26525 31331
rect 26525 31297 26559 31331
rect 26559 31297 26568 31331
rect 26516 31288 26568 31297
rect 26608 31331 26660 31340
rect 26608 31297 26617 31331
rect 26617 31297 26651 31331
rect 26651 31297 26660 31331
rect 26608 31288 26660 31297
rect 27068 31288 27120 31340
rect 27160 31331 27212 31340
rect 27160 31297 27169 31331
rect 27169 31297 27203 31331
rect 27203 31297 27212 31331
rect 27160 31288 27212 31297
rect 27252 31331 27304 31340
rect 27252 31297 27261 31331
rect 27261 31297 27295 31331
rect 27295 31297 27304 31331
rect 27252 31288 27304 31297
rect 28264 31331 28316 31340
rect 28264 31297 28273 31331
rect 28273 31297 28307 31331
rect 28307 31297 28316 31331
rect 28264 31288 28316 31297
rect 28448 31331 28500 31340
rect 28448 31297 28457 31331
rect 28457 31297 28491 31331
rect 28491 31297 28500 31331
rect 28448 31288 28500 31297
rect 29276 31288 29328 31340
rect 30748 31288 30800 31340
rect 30840 31288 30892 31340
rect 32772 31288 32824 31340
rect 26976 31195 27028 31204
rect 26976 31161 26985 31195
rect 26985 31161 27019 31195
rect 27019 31161 27028 31195
rect 26976 31152 27028 31161
rect 26700 31084 26752 31136
rect 27436 31220 27488 31272
rect 27712 31220 27764 31272
rect 28816 31220 28868 31272
rect 31576 31220 31628 31272
rect 27896 31195 27948 31204
rect 27896 31161 27905 31195
rect 27905 31161 27939 31195
rect 27939 31161 27948 31195
rect 27896 31152 27948 31161
rect 28264 31152 28316 31204
rect 33784 31356 33836 31408
rect 34244 31399 34296 31408
rect 34244 31365 34253 31399
rect 34253 31365 34287 31399
rect 34287 31365 34296 31399
rect 34244 31356 34296 31365
rect 34888 31424 34940 31476
rect 35440 31424 35492 31476
rect 34796 31356 34848 31408
rect 36176 31399 36228 31408
rect 36176 31365 36193 31399
rect 36193 31365 36228 31399
rect 36176 31356 36228 31365
rect 37740 31424 37792 31476
rect 37832 31424 37884 31476
rect 38384 31424 38436 31476
rect 38568 31424 38620 31476
rect 34336 31288 34388 31340
rect 35992 31331 36044 31340
rect 35992 31297 36001 31331
rect 36001 31297 36035 31331
rect 36035 31297 36044 31331
rect 35992 31288 36044 31297
rect 36360 31331 36412 31340
rect 36360 31297 36369 31331
rect 36369 31297 36403 31331
rect 36403 31297 36412 31331
rect 36360 31288 36412 31297
rect 36452 31331 36504 31340
rect 36452 31297 36461 31331
rect 36461 31297 36495 31331
rect 36495 31297 36504 31331
rect 36452 31288 36504 31297
rect 37188 31356 37240 31408
rect 37372 31288 37424 31340
rect 35440 31220 35492 31272
rect 38844 31356 38896 31408
rect 39488 31356 39540 31408
rect 37556 31220 37608 31272
rect 37464 31152 37516 31204
rect 38200 31288 38252 31340
rect 28080 31084 28132 31136
rect 28724 31084 28776 31136
rect 31576 31084 31628 31136
rect 33324 31084 33376 31136
rect 33600 31127 33652 31136
rect 33600 31093 33609 31127
rect 33609 31093 33643 31127
rect 33643 31093 33652 31127
rect 33600 31084 33652 31093
rect 34152 31084 34204 31136
rect 34796 31084 34848 31136
rect 37280 31084 37332 31136
rect 38568 31084 38620 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 4988 30880 5040 30932
rect 8024 30880 8076 30932
rect 8576 30923 8628 30932
rect 8576 30889 8585 30923
rect 8585 30889 8619 30923
rect 8619 30889 8628 30923
rect 8576 30880 8628 30889
rect 10784 30923 10836 30932
rect 10784 30889 10793 30923
rect 10793 30889 10827 30923
rect 10827 30889 10836 30923
rect 10784 30880 10836 30889
rect 11336 30923 11388 30932
rect 11336 30889 11345 30923
rect 11345 30889 11379 30923
rect 11379 30889 11388 30923
rect 11336 30880 11388 30889
rect 11888 30880 11940 30932
rect 15476 30880 15528 30932
rect 17408 30880 17460 30932
rect 17868 30880 17920 30932
rect 18420 30923 18472 30932
rect 18420 30889 18429 30923
rect 18429 30889 18463 30923
rect 18463 30889 18472 30923
rect 18420 30880 18472 30889
rect 18696 30923 18748 30932
rect 18696 30889 18705 30923
rect 18705 30889 18739 30923
rect 18739 30889 18748 30923
rect 18696 30880 18748 30889
rect 20996 30880 21048 30932
rect 22836 30923 22888 30932
rect 22836 30889 22845 30923
rect 22845 30889 22879 30923
rect 22879 30889 22888 30923
rect 22836 30880 22888 30889
rect 23204 30880 23256 30932
rect 23664 30923 23716 30932
rect 23664 30889 23673 30923
rect 23673 30889 23707 30923
rect 23707 30889 23716 30923
rect 23664 30880 23716 30889
rect 23848 30880 23900 30932
rect 26516 30880 26568 30932
rect 26700 30880 26752 30932
rect 3240 30744 3292 30796
rect 4804 30787 4856 30796
rect 4804 30753 4813 30787
rect 4813 30753 4847 30787
rect 4847 30753 4856 30787
rect 4804 30744 4856 30753
rect 3792 30676 3844 30728
rect 4896 30676 4948 30728
rect 6092 30719 6144 30728
rect 6092 30685 6101 30719
rect 6101 30685 6135 30719
rect 6135 30685 6144 30719
rect 6092 30676 6144 30685
rect 6552 30676 6604 30728
rect 7656 30676 7708 30728
rect 8392 30812 8444 30864
rect 8760 30812 8812 30864
rect 9128 30812 9180 30864
rect 8300 30744 8352 30796
rect 8208 30719 8260 30728
rect 8208 30685 8217 30719
rect 8217 30685 8251 30719
rect 8251 30685 8260 30719
rect 8208 30676 8260 30685
rect 9680 30787 9732 30796
rect 9680 30753 9689 30787
rect 9689 30753 9723 30787
rect 9723 30753 9732 30787
rect 9680 30744 9732 30753
rect 10508 30812 10560 30864
rect 10968 30812 11020 30864
rect 11520 30744 11572 30796
rect 1584 30651 1636 30660
rect 1584 30617 1593 30651
rect 1593 30617 1627 30651
rect 1627 30617 1636 30651
rect 1584 30608 1636 30617
rect 2688 30608 2740 30660
rect 3332 30651 3384 30660
rect 3332 30617 3341 30651
rect 3341 30617 3375 30651
rect 3375 30617 3384 30651
rect 3332 30608 3384 30617
rect 6184 30583 6236 30592
rect 6184 30549 6193 30583
rect 6193 30549 6227 30583
rect 6227 30549 6236 30583
rect 6184 30540 6236 30549
rect 10692 30719 10744 30728
rect 10692 30685 10701 30719
rect 10701 30685 10735 30719
rect 10735 30685 10744 30719
rect 10692 30676 10744 30685
rect 11060 30676 11112 30728
rect 11428 30719 11480 30728
rect 11428 30685 11437 30719
rect 11437 30685 11471 30719
rect 11471 30685 11480 30719
rect 11428 30676 11480 30685
rect 13084 30719 13136 30728
rect 13084 30685 13093 30719
rect 13093 30685 13127 30719
rect 13127 30685 13136 30719
rect 13084 30676 13136 30685
rect 12164 30608 12216 30660
rect 14188 30676 14240 30728
rect 15016 30676 15068 30728
rect 16672 30744 16724 30796
rect 15568 30719 15620 30728
rect 15568 30685 15577 30719
rect 15577 30685 15611 30719
rect 15611 30685 15620 30719
rect 15568 30676 15620 30685
rect 15660 30719 15712 30728
rect 15660 30685 15669 30719
rect 15669 30685 15703 30719
rect 15703 30685 15712 30719
rect 15660 30676 15712 30685
rect 10324 30540 10376 30592
rect 10600 30540 10652 30592
rect 12900 30540 12952 30592
rect 13268 30583 13320 30592
rect 13268 30549 13277 30583
rect 13277 30549 13311 30583
rect 13311 30549 13320 30583
rect 13268 30540 13320 30549
rect 15292 30540 15344 30592
rect 16488 30540 16540 30592
rect 17684 30608 17736 30660
rect 18328 30676 18380 30728
rect 18604 30608 18656 30660
rect 22928 30812 22980 30864
rect 27528 30812 27580 30864
rect 27712 30812 27764 30864
rect 27804 30855 27856 30864
rect 27804 30821 27813 30855
rect 27813 30821 27847 30855
rect 27847 30821 27856 30855
rect 27804 30812 27856 30821
rect 28356 30812 28408 30864
rect 28908 30812 28960 30864
rect 33600 30923 33652 30932
rect 33600 30889 33609 30923
rect 33609 30889 33643 30923
rect 33643 30889 33652 30923
rect 33600 30880 33652 30889
rect 34704 30880 34756 30932
rect 36360 30880 36412 30932
rect 37464 30880 37516 30932
rect 38292 30880 38344 30932
rect 20444 30744 20496 30796
rect 20812 30787 20864 30796
rect 20812 30753 20821 30787
rect 20821 30753 20855 30787
rect 20855 30753 20864 30787
rect 20812 30744 20864 30753
rect 21088 30787 21140 30796
rect 21088 30753 21097 30787
rect 21097 30753 21131 30787
rect 21131 30753 21140 30787
rect 21088 30744 21140 30753
rect 21732 30719 21784 30728
rect 21732 30685 21741 30719
rect 21741 30685 21775 30719
rect 21775 30685 21784 30719
rect 21732 30676 21784 30685
rect 23204 30719 23256 30728
rect 23204 30685 23213 30719
rect 23213 30685 23247 30719
rect 23247 30685 23256 30719
rect 23204 30676 23256 30685
rect 23572 30719 23624 30728
rect 23572 30685 23581 30719
rect 23581 30685 23615 30719
rect 23615 30685 23624 30719
rect 23572 30676 23624 30685
rect 23756 30676 23808 30728
rect 19432 30608 19484 30660
rect 21364 30608 21416 30660
rect 17776 30540 17828 30592
rect 20996 30540 21048 30592
rect 21824 30608 21876 30660
rect 26516 30744 26568 30796
rect 26240 30676 26292 30728
rect 22100 30540 22152 30592
rect 23388 30540 23440 30592
rect 23848 30540 23900 30592
rect 25872 30608 25924 30660
rect 26884 30719 26936 30728
rect 26884 30685 26893 30719
rect 26893 30685 26927 30719
rect 26927 30685 26936 30719
rect 26884 30676 26936 30685
rect 27620 30676 27672 30728
rect 28632 30744 28684 30796
rect 30472 30744 30524 30796
rect 27896 30676 27948 30728
rect 28172 30608 28224 30660
rect 28632 30608 28684 30660
rect 29000 30719 29052 30728
rect 29000 30685 29009 30719
rect 29009 30685 29043 30719
rect 29043 30685 29052 30719
rect 29000 30676 29052 30685
rect 29552 30719 29604 30728
rect 29552 30685 29561 30719
rect 29561 30685 29595 30719
rect 29595 30685 29604 30719
rect 29552 30676 29604 30685
rect 30380 30676 30432 30728
rect 30748 30676 30800 30728
rect 30104 30608 30156 30660
rect 30564 30608 30616 30660
rect 31208 30719 31260 30728
rect 31208 30685 31217 30719
rect 31217 30685 31251 30719
rect 31251 30685 31260 30719
rect 31208 30676 31260 30685
rect 34612 30812 34664 30864
rect 32128 30744 32180 30796
rect 32680 30744 32732 30796
rect 33692 30744 33744 30796
rect 36084 30812 36136 30864
rect 36820 30812 36872 30864
rect 37004 30812 37056 30864
rect 31576 30719 31628 30728
rect 31576 30685 31585 30719
rect 31585 30685 31619 30719
rect 31619 30685 31628 30719
rect 31576 30676 31628 30685
rect 31668 30651 31720 30660
rect 31668 30617 31677 30651
rect 31677 30617 31711 30651
rect 31711 30617 31720 30651
rect 31668 30608 31720 30617
rect 30288 30540 30340 30592
rect 31116 30540 31168 30592
rect 32036 30676 32088 30728
rect 33876 30719 33928 30728
rect 33876 30685 33885 30719
rect 33885 30685 33919 30719
rect 33919 30685 33928 30719
rect 33876 30676 33928 30685
rect 34336 30676 34388 30728
rect 36268 30787 36320 30796
rect 36268 30753 36277 30787
rect 36277 30753 36311 30787
rect 36311 30753 36320 30787
rect 36268 30744 36320 30753
rect 32312 30608 32364 30660
rect 32588 30608 32640 30660
rect 33324 30608 33376 30660
rect 36176 30676 36228 30728
rect 36820 30719 36872 30728
rect 36820 30685 36829 30719
rect 36829 30685 36863 30719
rect 36863 30685 36872 30719
rect 36820 30676 36872 30685
rect 37556 30744 37608 30796
rect 37372 30719 37424 30728
rect 37372 30685 37381 30719
rect 37381 30685 37415 30719
rect 37415 30685 37424 30719
rect 37372 30676 37424 30685
rect 37648 30676 37700 30728
rect 38292 30676 38344 30728
rect 33600 30540 33652 30592
rect 34244 30540 34296 30592
rect 36176 30540 36228 30592
rect 37464 30608 37516 30660
rect 38108 30608 38160 30660
rect 38752 30608 38804 30660
rect 39028 30608 39080 30660
rect 36728 30540 36780 30592
rect 37648 30583 37700 30592
rect 37648 30549 37657 30583
rect 37657 30549 37691 30583
rect 37691 30549 37700 30583
rect 37648 30540 37700 30549
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 1584 30336 1636 30388
rect 7840 30336 7892 30388
rect 8576 30336 8628 30388
rect 10692 30336 10744 30388
rect 13084 30336 13136 30388
rect 14280 30336 14332 30388
rect 3332 30268 3384 30320
rect 848 30200 900 30252
rect 2872 30243 2924 30252
rect 2872 30209 2881 30243
rect 2881 30209 2915 30243
rect 2915 30209 2924 30243
rect 2872 30200 2924 30209
rect 4804 30268 4856 30320
rect 4896 30268 4948 30320
rect 9404 30268 9456 30320
rect 11336 30268 11388 30320
rect 11612 30268 11664 30320
rect 11704 30268 11756 30320
rect 7380 30243 7432 30252
rect 7380 30209 7389 30243
rect 7389 30209 7423 30243
rect 7423 30209 7432 30243
rect 7380 30200 7432 30209
rect 10876 30243 10928 30252
rect 10876 30209 10885 30243
rect 10885 30209 10919 30243
rect 10919 30209 10928 30243
rect 10876 30200 10928 30209
rect 4620 30175 4672 30184
rect 4620 30141 4629 30175
rect 4629 30141 4663 30175
rect 4663 30141 4672 30175
rect 4620 30132 4672 30141
rect 4804 30175 4856 30184
rect 4804 30141 4813 30175
rect 4813 30141 4847 30175
rect 4847 30141 4856 30175
rect 4804 30132 4856 30141
rect 4896 30132 4948 30184
rect 5264 30132 5316 30184
rect 9864 30132 9916 30184
rect 11888 30175 11940 30184
rect 11888 30141 11897 30175
rect 11897 30141 11931 30175
rect 11931 30141 11940 30175
rect 11888 30132 11940 30141
rect 12440 30243 12492 30252
rect 12440 30209 12449 30243
rect 12449 30209 12483 30243
rect 12483 30209 12492 30243
rect 12440 30200 12492 30209
rect 5908 30064 5960 30116
rect 6184 30064 6236 30116
rect 7840 30064 7892 30116
rect 11980 30064 12032 30116
rect 12532 30064 12584 30116
rect 12900 30064 12952 30116
rect 13268 30268 13320 30320
rect 14188 30200 14240 30252
rect 14372 30200 14424 30252
rect 14648 30243 14700 30252
rect 14648 30209 14657 30243
rect 14657 30209 14691 30243
rect 14691 30209 14700 30243
rect 14648 30200 14700 30209
rect 15016 30200 15068 30252
rect 15108 30200 15160 30252
rect 15660 30268 15712 30320
rect 18236 30336 18288 30388
rect 13176 30132 13228 30184
rect 15568 30200 15620 30252
rect 21180 30268 21232 30320
rect 22376 30268 22428 30320
rect 23296 30336 23348 30388
rect 16028 30243 16080 30252
rect 16028 30209 16037 30243
rect 16037 30209 16071 30243
rect 16071 30209 16080 30243
rect 16028 30200 16080 30209
rect 4068 29996 4120 30048
rect 7656 29996 7708 30048
rect 9772 29996 9824 30048
rect 12348 29996 12400 30048
rect 15476 30132 15528 30184
rect 16304 30243 16356 30252
rect 16304 30209 16313 30243
rect 16313 30209 16347 30243
rect 16347 30209 16356 30243
rect 16304 30200 16356 30209
rect 16764 30200 16816 30252
rect 17132 30200 17184 30252
rect 18420 30200 18472 30252
rect 22100 30200 22152 30252
rect 23112 30200 23164 30252
rect 24216 30268 24268 30320
rect 23388 30243 23440 30252
rect 23388 30209 23433 30243
rect 23433 30209 23440 30243
rect 23388 30200 23440 30209
rect 23664 30200 23716 30252
rect 27528 30336 27580 30388
rect 29276 30336 29328 30388
rect 29920 30336 29972 30388
rect 25872 30311 25924 30320
rect 25872 30277 25881 30311
rect 25881 30277 25915 30311
rect 25915 30277 25924 30311
rect 25872 30268 25924 30277
rect 28080 30268 28132 30320
rect 28908 30268 28960 30320
rect 31760 30268 31812 30320
rect 31944 30268 31996 30320
rect 26424 30243 26476 30252
rect 26424 30209 26433 30243
rect 26433 30209 26467 30243
rect 26467 30209 26476 30243
rect 26424 30200 26476 30209
rect 17684 30132 17736 30184
rect 18604 30175 18656 30184
rect 18604 30141 18613 30175
rect 18613 30141 18647 30175
rect 18647 30141 18656 30175
rect 18604 30132 18656 30141
rect 21732 30132 21784 30184
rect 24492 30132 24544 30184
rect 24676 30132 24728 30184
rect 25596 30132 25648 30184
rect 26056 30132 26108 30184
rect 26240 30175 26292 30184
rect 26240 30141 26249 30175
rect 26249 30141 26283 30175
rect 26283 30141 26292 30175
rect 26240 30132 26292 30141
rect 30288 30243 30340 30252
rect 30288 30209 30297 30243
rect 30297 30209 30331 30243
rect 30331 30209 30340 30243
rect 30288 30200 30340 30209
rect 30472 30243 30524 30252
rect 30472 30209 30489 30243
rect 30489 30209 30524 30243
rect 30472 30200 30524 30209
rect 30564 30243 30616 30252
rect 30564 30209 30573 30243
rect 30573 30209 30607 30243
rect 30607 30209 30616 30243
rect 30564 30200 30616 30209
rect 31116 30200 31168 30252
rect 26884 30132 26936 30184
rect 29552 30132 29604 30184
rect 14280 29996 14332 30048
rect 15568 29996 15620 30048
rect 15936 29996 15988 30048
rect 16028 30039 16080 30048
rect 16028 30005 16037 30039
rect 16037 30005 16071 30039
rect 16071 30005 16080 30039
rect 16028 29996 16080 30005
rect 16948 30064 17000 30116
rect 16580 29996 16632 30048
rect 16764 30039 16816 30048
rect 16764 30005 16773 30039
rect 16773 30005 16807 30039
rect 16807 30005 16816 30039
rect 16764 29996 16816 30005
rect 17040 29996 17092 30048
rect 18696 30064 18748 30116
rect 25780 30064 25832 30116
rect 25964 30064 26016 30116
rect 30196 30175 30248 30184
rect 30196 30141 30205 30175
rect 30205 30141 30239 30175
rect 30239 30141 30248 30175
rect 30196 30132 30248 30141
rect 31300 30200 31352 30252
rect 31760 30132 31812 30184
rect 32128 30243 32180 30252
rect 32128 30209 32137 30243
rect 32137 30209 32171 30243
rect 32171 30209 32180 30243
rect 32128 30200 32180 30209
rect 32680 30336 32732 30388
rect 36360 30336 36412 30388
rect 36544 30336 36596 30388
rect 37924 30336 37976 30388
rect 33692 30268 33744 30320
rect 32312 30200 32364 30252
rect 33140 30200 33192 30252
rect 31392 30064 31444 30116
rect 32036 30064 32088 30116
rect 33416 30107 33468 30116
rect 33416 30073 33425 30107
rect 33425 30073 33459 30107
rect 33459 30073 33468 30107
rect 33416 30064 33468 30073
rect 23388 29996 23440 30048
rect 24216 29996 24268 30048
rect 25044 29996 25096 30048
rect 25412 29996 25464 30048
rect 26240 29996 26292 30048
rect 26976 29996 27028 30048
rect 31576 29996 31628 30048
rect 31668 30039 31720 30048
rect 31668 30005 31677 30039
rect 31677 30005 31711 30039
rect 31711 30005 31720 30039
rect 31668 29996 31720 30005
rect 32680 29996 32732 30048
rect 33600 29996 33652 30048
rect 34060 30132 34112 30184
rect 34152 30064 34204 30116
rect 36268 30243 36320 30252
rect 36268 30209 36277 30243
rect 36277 30209 36311 30243
rect 36311 30209 36320 30243
rect 36268 30200 36320 30209
rect 36820 30200 36872 30252
rect 37372 30200 37424 30252
rect 37556 30243 37608 30252
rect 37556 30209 37565 30243
rect 37565 30209 37599 30243
rect 37599 30209 37608 30243
rect 37556 30200 37608 30209
rect 39488 30268 39540 30320
rect 40040 30268 40092 30320
rect 36176 30132 36228 30184
rect 38016 30132 38068 30184
rect 38200 30243 38252 30252
rect 38200 30209 38209 30243
rect 38209 30209 38243 30243
rect 38243 30209 38252 30243
rect 38200 30200 38252 30209
rect 38476 30175 38528 30184
rect 38476 30141 38485 30175
rect 38485 30141 38519 30175
rect 38519 30141 38528 30175
rect 38476 30132 38528 30141
rect 34336 29996 34388 30048
rect 35348 29996 35400 30048
rect 36084 29996 36136 30048
rect 36360 29996 36412 30048
rect 37280 29996 37332 30048
rect 37372 30039 37424 30048
rect 37372 30005 37381 30039
rect 37381 30005 37415 30039
rect 37415 30005 37424 30039
rect 37372 29996 37424 30005
rect 37832 30039 37884 30048
rect 37832 30005 37841 30039
rect 37841 30005 37875 30039
rect 37875 30005 37884 30039
rect 37832 29996 37884 30005
rect 38292 29996 38344 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 4620 29792 4672 29844
rect 6828 29792 6880 29844
rect 11060 29792 11112 29844
rect 12256 29792 12308 29844
rect 14556 29792 14608 29844
rect 16304 29792 16356 29844
rect 18328 29835 18380 29844
rect 18328 29801 18337 29835
rect 18337 29801 18371 29835
rect 18371 29801 18380 29835
rect 18328 29792 18380 29801
rect 18512 29792 18564 29844
rect 21456 29792 21508 29844
rect 21916 29792 21968 29844
rect 4068 29699 4120 29708
rect 4068 29665 4077 29699
rect 4077 29665 4111 29699
rect 4111 29665 4120 29699
rect 4068 29656 4120 29665
rect 4804 29656 4856 29708
rect 6552 29656 6604 29708
rect 9404 29656 9456 29708
rect 10692 29724 10744 29776
rect 13452 29724 13504 29776
rect 14740 29724 14792 29776
rect 19156 29724 19208 29776
rect 10784 29656 10836 29708
rect 3792 29631 3844 29640
rect 3792 29597 3801 29631
rect 3801 29597 3835 29631
rect 3835 29597 3844 29631
rect 3792 29588 3844 29597
rect 6000 29588 6052 29640
rect 9956 29588 10008 29640
rect 10692 29588 10744 29640
rect 11336 29588 11388 29640
rect 11796 29631 11848 29640
rect 11796 29597 11805 29631
rect 11805 29597 11839 29631
rect 11839 29597 11848 29631
rect 11796 29588 11848 29597
rect 7196 29520 7248 29572
rect 5724 29452 5776 29504
rect 6184 29452 6236 29504
rect 9680 29520 9732 29572
rect 11520 29520 11572 29572
rect 9496 29452 9548 29504
rect 13084 29656 13136 29708
rect 12348 29631 12400 29640
rect 12348 29597 12357 29631
rect 12357 29597 12391 29631
rect 12391 29597 12400 29631
rect 12348 29588 12400 29597
rect 12532 29588 12584 29640
rect 12164 29452 12216 29504
rect 12348 29452 12400 29504
rect 12900 29631 12952 29640
rect 12900 29597 12909 29631
rect 12909 29597 12943 29631
rect 12943 29597 12952 29631
rect 12900 29588 12952 29597
rect 15476 29699 15528 29708
rect 15476 29665 15485 29699
rect 15485 29665 15519 29699
rect 15519 29665 15528 29699
rect 15476 29656 15528 29665
rect 14096 29631 14148 29640
rect 14096 29597 14105 29631
rect 14105 29597 14139 29631
rect 14139 29597 14148 29631
rect 14096 29588 14148 29597
rect 14372 29631 14424 29640
rect 14372 29597 14381 29631
rect 14381 29597 14415 29631
rect 14415 29597 14424 29631
rect 14372 29588 14424 29597
rect 14648 29588 14700 29640
rect 14924 29588 14976 29640
rect 15016 29588 15068 29640
rect 14188 29520 14240 29572
rect 15752 29588 15804 29640
rect 16488 29631 16540 29640
rect 16488 29597 16497 29631
rect 16497 29597 16531 29631
rect 16531 29597 16540 29631
rect 16488 29588 16540 29597
rect 16948 29588 17000 29640
rect 17132 29631 17184 29640
rect 17132 29597 17141 29631
rect 17141 29597 17175 29631
rect 17175 29597 17184 29631
rect 17132 29588 17184 29597
rect 19984 29656 20036 29708
rect 13176 29495 13228 29504
rect 13176 29461 13185 29495
rect 13185 29461 13219 29495
rect 13219 29461 13228 29495
rect 13176 29452 13228 29461
rect 13820 29452 13872 29504
rect 16764 29520 16816 29572
rect 18512 29631 18564 29640
rect 18512 29597 18521 29631
rect 18521 29597 18555 29631
rect 18555 29597 18564 29631
rect 18512 29588 18564 29597
rect 18788 29631 18840 29640
rect 18788 29597 18797 29631
rect 18797 29597 18831 29631
rect 18831 29597 18840 29631
rect 18788 29588 18840 29597
rect 18880 29631 18932 29640
rect 18880 29597 18889 29631
rect 18889 29597 18923 29631
rect 18923 29597 18932 29631
rect 18880 29588 18932 29597
rect 18972 29588 19024 29640
rect 19432 29563 19484 29572
rect 19432 29529 19441 29563
rect 19441 29529 19475 29563
rect 19475 29529 19484 29563
rect 23020 29656 23072 29708
rect 22284 29631 22336 29640
rect 22284 29597 22293 29631
rect 22293 29597 22327 29631
rect 22327 29597 22336 29631
rect 22284 29588 22336 29597
rect 22652 29631 22704 29640
rect 22652 29597 22661 29631
rect 22661 29597 22695 29631
rect 22695 29597 22704 29631
rect 22652 29588 22704 29597
rect 22744 29588 22796 29640
rect 23480 29724 23532 29776
rect 23848 29724 23900 29776
rect 24124 29724 24176 29776
rect 23388 29631 23440 29640
rect 23388 29597 23397 29631
rect 23397 29597 23431 29631
rect 23431 29597 23440 29631
rect 23388 29588 23440 29597
rect 23572 29588 23624 29640
rect 24216 29656 24268 29708
rect 23848 29588 23900 29640
rect 24032 29588 24084 29640
rect 26424 29724 26476 29776
rect 27436 29792 27488 29844
rect 33876 29792 33928 29844
rect 35256 29792 35308 29844
rect 36452 29792 36504 29844
rect 38384 29835 38436 29844
rect 38384 29801 38393 29835
rect 38393 29801 38427 29835
rect 38427 29801 38436 29835
rect 38384 29792 38436 29801
rect 27804 29724 27856 29776
rect 27896 29724 27948 29776
rect 31024 29724 31076 29776
rect 25044 29656 25096 29708
rect 19432 29520 19484 29529
rect 22560 29520 22612 29572
rect 25136 29631 25188 29640
rect 25136 29597 25145 29631
rect 25145 29597 25179 29631
rect 25179 29597 25188 29631
rect 25136 29588 25188 29597
rect 25320 29631 25372 29640
rect 25320 29597 25329 29631
rect 25329 29597 25363 29631
rect 25363 29597 25372 29631
rect 25320 29588 25372 29597
rect 28540 29656 28592 29708
rect 19524 29452 19576 29504
rect 20720 29452 20772 29504
rect 21916 29452 21968 29504
rect 22468 29452 22520 29504
rect 23572 29495 23624 29504
rect 23572 29461 23581 29495
rect 23581 29461 23615 29495
rect 23615 29461 23624 29495
rect 23572 29452 23624 29461
rect 24216 29452 24268 29504
rect 24860 29520 24912 29572
rect 25688 29520 25740 29572
rect 26240 29631 26292 29640
rect 26240 29597 26249 29631
rect 26249 29597 26283 29631
rect 26283 29597 26292 29631
rect 26240 29588 26292 29597
rect 26516 29631 26568 29640
rect 26516 29597 26525 29631
rect 26525 29597 26559 29631
rect 26559 29597 26568 29631
rect 26516 29588 26568 29597
rect 26884 29588 26936 29640
rect 26148 29520 26200 29572
rect 27528 29520 27580 29572
rect 28264 29588 28316 29640
rect 28356 29631 28408 29640
rect 28356 29597 28365 29631
rect 28365 29597 28399 29631
rect 28399 29597 28408 29631
rect 28356 29588 28408 29597
rect 31760 29656 31812 29708
rect 31852 29656 31904 29708
rect 33048 29656 33100 29708
rect 33600 29724 33652 29776
rect 34244 29724 34296 29776
rect 34888 29767 34940 29776
rect 34888 29733 34897 29767
rect 34897 29733 34931 29767
rect 34931 29733 34940 29767
rect 34888 29724 34940 29733
rect 35164 29724 35216 29776
rect 36084 29724 36136 29776
rect 33508 29656 33560 29708
rect 28540 29520 28592 29572
rect 24676 29452 24728 29504
rect 28264 29452 28316 29504
rect 30472 29631 30524 29640
rect 30472 29597 30481 29631
rect 30481 29597 30515 29631
rect 30515 29597 30524 29631
rect 30472 29588 30524 29597
rect 30748 29495 30800 29504
rect 30748 29461 30757 29495
rect 30757 29461 30791 29495
rect 30791 29461 30800 29495
rect 30748 29452 30800 29461
rect 32772 29631 32824 29640
rect 32772 29597 32781 29631
rect 32781 29597 32815 29631
rect 32815 29597 32824 29631
rect 32772 29588 32824 29597
rect 32864 29631 32916 29640
rect 32864 29597 32873 29631
rect 32873 29597 32907 29631
rect 32907 29597 32916 29631
rect 32864 29588 32916 29597
rect 33324 29588 33376 29640
rect 33968 29588 34020 29640
rect 36176 29656 36228 29708
rect 34152 29631 34204 29640
rect 34152 29597 34161 29631
rect 34161 29597 34195 29631
rect 34195 29597 34204 29631
rect 34152 29588 34204 29597
rect 34244 29588 34296 29640
rect 30932 29520 30984 29572
rect 33048 29520 33100 29572
rect 31852 29452 31904 29504
rect 31944 29452 31996 29504
rect 33232 29452 33284 29504
rect 33784 29452 33836 29504
rect 34704 29631 34756 29640
rect 34704 29597 34713 29631
rect 34713 29597 34747 29631
rect 34747 29597 34756 29631
rect 34704 29588 34756 29597
rect 35440 29588 35492 29640
rect 36544 29724 36596 29776
rect 38016 29724 38068 29776
rect 36636 29656 36688 29708
rect 34152 29452 34204 29504
rect 35072 29520 35124 29572
rect 35624 29563 35676 29572
rect 35624 29529 35633 29563
rect 35633 29529 35667 29563
rect 35667 29529 35676 29563
rect 35624 29520 35676 29529
rect 36820 29588 36872 29640
rect 37464 29588 37516 29640
rect 37648 29588 37700 29640
rect 37832 29588 37884 29640
rect 38384 29656 38436 29708
rect 37372 29520 37424 29572
rect 35992 29452 36044 29504
rect 36176 29452 36228 29504
rect 38016 29452 38068 29504
rect 38384 29563 38436 29572
rect 38384 29529 38393 29563
rect 38393 29529 38427 29563
rect 38427 29529 38436 29563
rect 38384 29520 38436 29529
rect 38660 29631 38712 29640
rect 38660 29597 38669 29631
rect 38669 29597 38703 29631
rect 38703 29597 38712 29631
rect 38660 29588 38712 29597
rect 38936 29588 38988 29640
rect 39120 29631 39172 29640
rect 39120 29597 39129 29631
rect 39129 29597 39163 29631
rect 39163 29597 39172 29631
rect 39120 29588 39172 29597
rect 38660 29452 38712 29504
rect 38844 29563 38896 29572
rect 38844 29529 38853 29563
rect 38853 29529 38887 29563
rect 38887 29529 38896 29563
rect 38844 29520 38896 29529
rect 39212 29452 39264 29504
rect 39304 29495 39356 29504
rect 39304 29461 39313 29495
rect 39313 29461 39347 29495
rect 39347 29461 39356 29495
rect 39304 29452 39356 29461
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 3792 29248 3844 29300
rect 5540 29248 5592 29300
rect 6828 29248 6880 29300
rect 7196 29180 7248 29232
rect 7748 29180 7800 29232
rect 6184 29112 6236 29164
rect 4804 29044 4856 29096
rect 6828 29087 6880 29096
rect 6828 29053 6837 29087
rect 6837 29053 6871 29087
rect 6871 29053 6880 29087
rect 6828 29044 6880 29053
rect 7104 29087 7156 29096
rect 7104 29053 7113 29087
rect 7113 29053 7147 29087
rect 7147 29053 7156 29087
rect 7104 29044 7156 29053
rect 7196 29044 7248 29096
rect 7748 29044 7800 29096
rect 6000 28976 6052 29028
rect 6184 29019 6236 29028
rect 6184 28985 6193 29019
rect 6193 28985 6227 29019
rect 6227 28985 6236 29019
rect 6184 28976 6236 28985
rect 8760 28976 8812 29028
rect 9496 29180 9548 29232
rect 9772 29223 9824 29232
rect 9772 29189 9781 29223
rect 9781 29189 9815 29223
rect 9815 29189 9824 29223
rect 9772 29180 9824 29189
rect 11060 29180 11112 29232
rect 11336 29291 11388 29300
rect 11336 29257 11345 29291
rect 11345 29257 11379 29291
rect 11379 29257 11388 29291
rect 11336 29248 11388 29257
rect 11704 29248 11756 29300
rect 12440 29248 12492 29300
rect 14372 29248 14424 29300
rect 16764 29248 16816 29300
rect 19524 29291 19576 29300
rect 19524 29257 19533 29291
rect 19533 29257 19567 29291
rect 19567 29257 19576 29291
rect 19524 29248 19576 29257
rect 9496 29044 9548 29096
rect 9956 29019 10008 29028
rect 9956 28985 9965 29019
rect 9965 28985 9999 29019
rect 9999 28985 10008 29019
rect 9956 28976 10008 28985
rect 10784 29044 10836 29096
rect 11336 29112 11388 29164
rect 11980 29180 12032 29232
rect 12348 29180 12400 29232
rect 12624 29180 12676 29232
rect 14648 29180 14700 29232
rect 11704 29112 11756 29164
rect 12164 29112 12216 29164
rect 12440 29155 12492 29164
rect 12440 29121 12449 29155
rect 12449 29121 12483 29155
rect 12483 29121 12492 29155
rect 12440 29112 12492 29121
rect 11336 28976 11388 29028
rect 12532 29044 12584 29096
rect 15016 29087 15068 29096
rect 15016 29053 15025 29087
rect 15025 29053 15059 29087
rect 15059 29053 15068 29087
rect 15016 29044 15068 29053
rect 15292 29087 15344 29096
rect 15292 29053 15301 29087
rect 15301 29053 15335 29087
rect 15335 29053 15344 29087
rect 15292 29044 15344 29053
rect 5724 28908 5776 28960
rect 8668 28951 8720 28960
rect 8668 28917 8677 28951
rect 8677 28917 8711 28951
rect 8711 28917 8720 28951
rect 8668 28908 8720 28917
rect 9496 28951 9548 28960
rect 9496 28917 9505 28951
rect 9505 28917 9539 28951
rect 9539 28917 9548 28951
rect 9496 28908 9548 28917
rect 9680 28908 9732 28960
rect 10416 28951 10468 28960
rect 10416 28917 10425 28951
rect 10425 28917 10459 28951
rect 10459 28917 10468 28951
rect 10416 28908 10468 28917
rect 10692 28908 10744 28960
rect 11704 28908 11756 28960
rect 13820 28976 13872 29028
rect 16028 29180 16080 29232
rect 15844 29155 15896 29164
rect 15844 29121 15853 29155
rect 15853 29121 15887 29155
rect 15887 29121 15896 29155
rect 15844 29112 15896 29121
rect 16488 29112 16540 29164
rect 16764 29044 16816 29096
rect 17040 29155 17092 29164
rect 17040 29121 17049 29155
rect 17049 29121 17083 29155
rect 17083 29121 17092 29155
rect 17040 29112 17092 29121
rect 18788 29180 18840 29232
rect 17592 29155 17644 29164
rect 17592 29121 17601 29155
rect 17601 29121 17635 29155
rect 17635 29121 17644 29155
rect 17592 29112 17644 29121
rect 17868 29155 17920 29164
rect 17868 29121 17877 29155
rect 17877 29121 17911 29155
rect 17911 29121 17920 29155
rect 17868 29112 17920 29121
rect 18972 29087 19024 29096
rect 18972 29053 18981 29087
rect 18981 29053 19015 29087
rect 19015 29053 19024 29087
rect 20720 29112 20772 29164
rect 20904 29155 20956 29164
rect 20904 29121 20913 29155
rect 20913 29121 20947 29155
rect 20947 29121 20956 29155
rect 20904 29112 20956 29121
rect 18972 29044 19024 29053
rect 20812 29044 20864 29096
rect 16948 29019 17000 29028
rect 16948 28985 16957 29019
rect 16957 28985 16991 29019
rect 16991 28985 17000 29019
rect 16948 28976 17000 28985
rect 18604 28976 18656 29028
rect 20720 29019 20772 29028
rect 20720 28985 20729 29019
rect 20729 28985 20763 29019
rect 20763 28985 20772 29019
rect 20720 28976 20772 28985
rect 21180 29180 21232 29232
rect 26976 29248 27028 29300
rect 22652 29180 22704 29232
rect 23664 29180 23716 29232
rect 21088 29155 21140 29164
rect 21088 29121 21097 29155
rect 21097 29121 21131 29155
rect 21131 29121 21140 29155
rect 21088 29112 21140 29121
rect 21456 29112 21508 29164
rect 21548 29155 21600 29164
rect 21548 29121 21557 29155
rect 21557 29121 21591 29155
rect 21591 29121 21600 29155
rect 21548 29112 21600 29121
rect 21272 29087 21324 29096
rect 21272 29053 21281 29087
rect 21281 29053 21315 29087
rect 21315 29053 21324 29087
rect 23020 29112 23072 29164
rect 23480 29112 23532 29164
rect 23572 29155 23624 29164
rect 23572 29121 23581 29155
rect 23581 29121 23615 29155
rect 23615 29121 23624 29155
rect 23572 29112 23624 29121
rect 23848 29155 23900 29164
rect 23848 29121 23857 29155
rect 23857 29121 23891 29155
rect 23891 29121 23900 29155
rect 23848 29112 23900 29121
rect 24032 29155 24084 29164
rect 24032 29121 24041 29155
rect 24041 29121 24075 29155
rect 24075 29121 24084 29155
rect 24032 29112 24084 29121
rect 21272 29044 21324 29053
rect 22376 29044 22428 29096
rect 22560 29044 22612 29096
rect 24492 29112 24544 29164
rect 16028 28908 16080 28960
rect 19156 28951 19208 28960
rect 19156 28917 19184 28951
rect 19184 28917 19208 28951
rect 21732 28976 21784 29028
rect 22284 28976 22336 29028
rect 19156 28908 19208 28917
rect 23020 28908 23072 28960
rect 23848 28976 23900 29028
rect 23480 28908 23532 28960
rect 23664 28951 23716 28960
rect 23664 28917 23673 28951
rect 23673 28917 23707 28951
rect 23707 28917 23716 28951
rect 23664 28908 23716 28917
rect 24492 28908 24544 28960
rect 24768 29155 24820 29164
rect 24768 29121 24777 29155
rect 24777 29121 24811 29155
rect 24811 29121 24820 29155
rect 24768 29112 24820 29121
rect 25136 29180 25188 29232
rect 25780 29180 25832 29232
rect 27436 29248 27488 29300
rect 29736 29248 29788 29300
rect 30748 29248 30800 29300
rect 31484 29248 31536 29300
rect 28540 29223 28592 29232
rect 25412 29155 25464 29164
rect 25412 29121 25421 29155
rect 25421 29121 25455 29155
rect 25455 29121 25464 29155
rect 25412 29112 25464 29121
rect 25504 29112 25556 29164
rect 25596 29155 25648 29164
rect 25596 29121 25605 29155
rect 25605 29121 25639 29155
rect 25639 29121 25648 29155
rect 25596 29112 25648 29121
rect 26240 29112 26292 29164
rect 26424 29155 26476 29164
rect 26424 29121 26433 29155
rect 26433 29121 26467 29155
rect 26467 29121 26476 29155
rect 26424 29112 26476 29121
rect 28540 29189 28575 29223
rect 28575 29189 28592 29223
rect 28540 29180 28592 29189
rect 31760 29223 31812 29232
rect 31760 29189 31769 29223
rect 31769 29189 31803 29223
rect 31803 29189 31812 29223
rect 31760 29180 31812 29189
rect 32772 29248 32824 29300
rect 33692 29248 33744 29300
rect 35072 29248 35124 29300
rect 33508 29180 33560 29232
rect 27528 29155 27580 29164
rect 27528 29121 27537 29155
rect 27537 29121 27571 29155
rect 27571 29121 27580 29155
rect 27528 29112 27580 29121
rect 28264 29155 28316 29164
rect 28264 29121 28273 29155
rect 28273 29121 28307 29155
rect 28307 29121 28316 29155
rect 28264 29112 28316 29121
rect 28356 29155 28408 29164
rect 28356 29121 28365 29155
rect 28365 29121 28399 29155
rect 28399 29121 28408 29155
rect 28356 29112 28408 29121
rect 28448 29155 28500 29164
rect 28448 29121 28457 29155
rect 28457 29121 28491 29155
rect 28491 29121 28500 29155
rect 28448 29112 28500 29121
rect 30380 29112 30432 29164
rect 32404 29155 32456 29164
rect 25136 29087 25188 29096
rect 25136 29053 25145 29087
rect 25145 29053 25179 29087
rect 25179 29053 25188 29087
rect 25136 29044 25188 29053
rect 27436 29087 27488 29096
rect 27436 29053 27445 29087
rect 27445 29053 27479 29087
rect 27479 29053 27488 29087
rect 27436 29044 27488 29053
rect 28724 29087 28776 29096
rect 28724 29053 28733 29087
rect 28733 29053 28767 29087
rect 28767 29053 28776 29087
rect 28724 29044 28776 29053
rect 32404 29121 32408 29155
rect 32408 29121 32442 29155
rect 32442 29121 32456 29155
rect 32404 29112 32456 29121
rect 32680 29155 32732 29164
rect 32680 29121 32725 29155
rect 32725 29121 32732 29155
rect 32680 29112 32732 29121
rect 33048 29112 33100 29164
rect 34336 29180 34388 29232
rect 34520 29180 34572 29232
rect 33692 29155 33744 29164
rect 33692 29121 33701 29155
rect 33701 29121 33735 29155
rect 33735 29121 33744 29155
rect 33692 29112 33744 29121
rect 34152 29112 34204 29164
rect 34612 29155 34664 29164
rect 34612 29121 34621 29155
rect 34621 29121 34655 29155
rect 34655 29121 34664 29155
rect 34612 29112 34664 29121
rect 34980 29155 35032 29164
rect 34980 29121 34989 29155
rect 34989 29121 35023 29155
rect 35023 29121 35032 29155
rect 34980 29112 35032 29121
rect 24860 28976 24912 29028
rect 25320 28976 25372 29028
rect 26700 28976 26752 29028
rect 28816 29019 28868 29028
rect 28816 28985 28825 29019
rect 28825 28985 28859 29019
rect 28859 28985 28868 29019
rect 28816 28976 28868 28985
rect 32220 28976 32272 29028
rect 28264 28908 28316 28960
rect 32864 28976 32916 29028
rect 35532 29223 35584 29232
rect 35532 29189 35541 29223
rect 35541 29189 35575 29223
rect 35575 29189 35584 29223
rect 35532 29180 35584 29189
rect 36084 29248 36136 29300
rect 36452 29180 36504 29232
rect 36728 29223 36780 29232
rect 36728 29189 36755 29223
rect 36755 29189 36780 29223
rect 36728 29180 36780 29189
rect 36912 29223 36964 29232
rect 36912 29189 36921 29223
rect 36921 29189 36955 29223
rect 36955 29189 36964 29223
rect 36912 29180 36964 29189
rect 36084 29112 36136 29164
rect 36268 29112 36320 29164
rect 36544 29112 36596 29164
rect 37280 29155 37332 29164
rect 37280 29121 37289 29155
rect 37289 29121 37323 29155
rect 37323 29121 37332 29155
rect 37280 29112 37332 29121
rect 39212 29248 39264 29300
rect 38476 29223 38528 29232
rect 38476 29189 38485 29223
rect 38485 29189 38519 29223
rect 38519 29189 38528 29223
rect 38476 29180 38528 29189
rect 39488 29180 39540 29232
rect 37832 29112 37884 29164
rect 38200 29155 38252 29164
rect 38200 29121 38209 29155
rect 38209 29121 38243 29155
rect 38243 29121 38252 29155
rect 38200 29112 38252 29121
rect 33876 29019 33928 29028
rect 33876 28985 33885 29019
rect 33885 28985 33919 29019
rect 33919 28985 33928 29019
rect 33876 28976 33928 28985
rect 34060 28976 34112 29028
rect 34152 28976 34204 29028
rect 38936 29044 38988 29096
rect 33140 28908 33192 28960
rect 33600 28908 33652 28960
rect 34244 28951 34296 28960
rect 34244 28917 34253 28951
rect 34253 28917 34287 28951
rect 34287 28917 34296 28951
rect 34244 28908 34296 28917
rect 34428 28908 34480 28960
rect 35256 29019 35308 29028
rect 35256 28985 35265 29019
rect 35265 28985 35299 29019
rect 35299 28985 35308 29019
rect 35256 28976 35308 28985
rect 35808 29019 35860 29028
rect 35808 28985 35817 29019
rect 35817 28985 35851 29019
rect 35851 28985 35860 29019
rect 35808 28976 35860 28985
rect 36268 28976 36320 29028
rect 37556 28976 37608 29028
rect 37740 28976 37792 29028
rect 38200 28976 38252 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 6184 28704 6236 28756
rect 7104 28704 7156 28756
rect 9864 28636 9916 28688
rect 11796 28704 11848 28756
rect 11888 28704 11940 28756
rect 14372 28704 14424 28756
rect 16396 28704 16448 28756
rect 20904 28704 20956 28756
rect 24032 28747 24084 28756
rect 24032 28713 24041 28747
rect 24041 28713 24075 28747
rect 24075 28713 24084 28747
rect 24032 28704 24084 28713
rect 24400 28704 24452 28756
rect 26240 28747 26292 28756
rect 26240 28713 26249 28747
rect 26249 28713 26283 28747
rect 26283 28713 26292 28747
rect 26240 28704 26292 28713
rect 26700 28747 26752 28756
rect 26700 28713 26709 28747
rect 26709 28713 26743 28747
rect 26743 28713 26752 28747
rect 26700 28704 26752 28713
rect 27068 28704 27120 28756
rect 29644 28704 29696 28756
rect 29920 28704 29972 28756
rect 32404 28704 32456 28756
rect 32588 28704 32640 28756
rect 34152 28704 34204 28756
rect 34428 28704 34480 28756
rect 36452 28704 36504 28756
rect 38108 28704 38160 28756
rect 38384 28704 38436 28756
rect 5540 28611 5592 28620
rect 5540 28577 5549 28611
rect 5549 28577 5583 28611
rect 5583 28577 5592 28611
rect 5540 28568 5592 28577
rect 6828 28568 6880 28620
rect 8484 28568 8536 28620
rect 8668 28500 8720 28552
rect 9680 28500 9732 28552
rect 10416 28543 10468 28552
rect 10416 28509 10425 28543
rect 10425 28509 10459 28543
rect 10459 28509 10468 28543
rect 10416 28500 10468 28509
rect 10692 28500 10744 28552
rect 11612 28568 11664 28620
rect 13912 28636 13964 28688
rect 15568 28636 15620 28688
rect 17592 28636 17644 28688
rect 11704 28500 11756 28552
rect 14740 28568 14792 28620
rect 16948 28568 17000 28620
rect 3884 28432 3936 28484
rect 4620 28432 4672 28484
rect 5816 28475 5868 28484
rect 5816 28441 5825 28475
rect 5825 28441 5859 28475
rect 5859 28441 5868 28475
rect 5816 28432 5868 28441
rect 4068 28364 4120 28416
rect 6460 28364 6512 28416
rect 10784 28475 10836 28484
rect 10784 28441 10793 28475
rect 10793 28441 10827 28475
rect 10827 28441 10836 28475
rect 10784 28432 10836 28441
rect 12256 28500 12308 28552
rect 13360 28500 13412 28552
rect 14280 28543 14332 28552
rect 14280 28509 14289 28543
rect 14289 28509 14323 28543
rect 14323 28509 14332 28543
rect 14280 28500 14332 28509
rect 14648 28543 14700 28552
rect 14648 28509 14657 28543
rect 14657 28509 14691 28543
rect 14691 28509 14700 28543
rect 14648 28500 14700 28509
rect 17868 28611 17920 28620
rect 17868 28577 17877 28611
rect 17877 28577 17911 28611
rect 17911 28577 17920 28611
rect 17868 28568 17920 28577
rect 21180 28543 21232 28552
rect 21180 28509 21189 28543
rect 21189 28509 21223 28543
rect 21223 28509 21232 28543
rect 21180 28500 21232 28509
rect 21364 28500 21416 28552
rect 22100 28543 22152 28552
rect 22100 28509 22109 28543
rect 22109 28509 22143 28543
rect 22143 28509 22152 28543
rect 22100 28500 22152 28509
rect 7288 28407 7340 28416
rect 7288 28373 7297 28407
rect 7297 28373 7331 28407
rect 7331 28373 7340 28407
rect 7288 28364 7340 28373
rect 8300 28364 8352 28416
rect 8852 28364 8904 28416
rect 10232 28364 10284 28416
rect 12440 28432 12492 28484
rect 11704 28364 11756 28416
rect 11796 28364 11848 28416
rect 12072 28364 12124 28416
rect 14096 28407 14148 28416
rect 14096 28373 14105 28407
rect 14105 28373 14139 28407
rect 14139 28373 14148 28407
rect 14096 28364 14148 28373
rect 15016 28432 15068 28484
rect 16120 28364 16172 28416
rect 20904 28364 20956 28416
rect 21088 28364 21140 28416
rect 23572 28568 23624 28620
rect 24676 28636 24728 28688
rect 22468 28543 22520 28552
rect 22468 28509 22477 28543
rect 22477 28509 22511 28543
rect 22511 28509 22520 28543
rect 22468 28500 22520 28509
rect 23388 28500 23440 28552
rect 23480 28543 23532 28552
rect 23480 28509 23489 28543
rect 23489 28509 23523 28543
rect 23523 28509 23532 28543
rect 23480 28500 23532 28509
rect 23756 28500 23808 28552
rect 24676 28500 24728 28552
rect 24768 28543 24820 28552
rect 24768 28509 24777 28543
rect 24777 28509 24811 28543
rect 24811 28509 24820 28543
rect 24768 28500 24820 28509
rect 25044 28500 25096 28552
rect 25136 28543 25188 28552
rect 25136 28509 25145 28543
rect 25145 28509 25179 28543
rect 25179 28509 25188 28543
rect 25136 28500 25188 28509
rect 25596 28568 25648 28620
rect 25872 28568 25924 28620
rect 25504 28543 25556 28552
rect 25504 28509 25513 28543
rect 25513 28509 25547 28543
rect 25547 28509 25556 28543
rect 25504 28500 25556 28509
rect 25780 28543 25832 28552
rect 25780 28509 25789 28543
rect 25789 28509 25823 28543
rect 25823 28509 25832 28543
rect 25780 28500 25832 28509
rect 27344 28636 27396 28688
rect 27528 28568 27580 28620
rect 24216 28475 24268 28484
rect 24216 28441 24225 28475
rect 24225 28441 24259 28475
rect 24259 28441 24268 28475
rect 24216 28432 24268 28441
rect 26148 28500 26200 28552
rect 26516 28543 26568 28552
rect 26516 28509 26525 28543
rect 26525 28509 26559 28543
rect 26559 28509 26568 28543
rect 26516 28500 26568 28509
rect 27436 28500 27488 28552
rect 27896 28500 27948 28552
rect 38292 28636 38344 28688
rect 28264 28543 28316 28552
rect 28264 28509 28273 28543
rect 28273 28509 28307 28543
rect 28307 28509 28316 28543
rect 28264 28500 28316 28509
rect 28816 28500 28868 28552
rect 29736 28543 29788 28552
rect 29736 28509 29745 28543
rect 29745 28509 29779 28543
rect 29779 28509 29788 28543
rect 29736 28500 29788 28509
rect 29920 28543 29972 28552
rect 29920 28509 29929 28543
rect 29929 28509 29963 28543
rect 29963 28509 29972 28543
rect 29920 28500 29972 28509
rect 31944 28568 31996 28620
rect 32680 28568 32732 28620
rect 32956 28568 33008 28620
rect 35440 28568 35492 28620
rect 35808 28568 35860 28620
rect 38844 28611 38896 28620
rect 38844 28577 38853 28611
rect 38853 28577 38887 28611
rect 38887 28577 38896 28611
rect 38844 28568 38896 28577
rect 39764 28568 39816 28620
rect 22652 28364 22704 28416
rect 23112 28407 23164 28416
rect 23112 28373 23121 28407
rect 23121 28373 23155 28407
rect 23155 28373 23164 28407
rect 23112 28364 23164 28373
rect 23756 28364 23808 28416
rect 29276 28432 29328 28484
rect 26516 28407 26568 28416
rect 26516 28373 26525 28407
rect 26525 28373 26559 28407
rect 26559 28373 26568 28407
rect 26516 28364 26568 28373
rect 28540 28407 28592 28416
rect 28540 28373 28549 28407
rect 28549 28373 28583 28407
rect 28583 28373 28592 28407
rect 28540 28364 28592 28373
rect 29184 28364 29236 28416
rect 29828 28475 29880 28484
rect 29828 28441 29837 28475
rect 29837 28441 29871 28475
rect 29871 28441 29880 28475
rect 29828 28432 29880 28441
rect 30012 28432 30064 28484
rect 30656 28432 30708 28484
rect 32220 28500 32272 28552
rect 32588 28543 32640 28552
rect 32588 28509 32597 28543
rect 32597 28509 32631 28543
rect 32631 28509 32640 28543
rect 32588 28500 32640 28509
rect 33600 28543 33652 28552
rect 33600 28509 33609 28543
rect 33609 28509 33643 28543
rect 33643 28509 33652 28543
rect 33600 28500 33652 28509
rect 34244 28500 34296 28552
rect 35532 28500 35584 28552
rect 35992 28543 36044 28552
rect 35992 28509 36001 28543
rect 36001 28509 36035 28543
rect 36035 28509 36044 28543
rect 35992 28500 36044 28509
rect 38016 28500 38068 28552
rect 39212 28500 39264 28552
rect 33508 28432 33560 28484
rect 33692 28432 33744 28484
rect 34336 28432 34388 28484
rect 36176 28432 36228 28484
rect 38108 28432 38160 28484
rect 30380 28364 30432 28416
rect 33416 28364 33468 28416
rect 34244 28364 34296 28416
rect 35624 28364 35676 28416
rect 36084 28364 36136 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 4068 28092 4120 28144
rect 5816 28160 5868 28212
rect 6460 28160 6512 28212
rect 14648 28160 14700 28212
rect 6000 28092 6052 28144
rect 4712 28067 4764 28076
rect 4712 28033 4721 28067
rect 4721 28033 4755 28067
rect 4755 28033 4764 28067
rect 4712 28024 4764 28033
rect 6368 28024 6420 28076
rect 6552 28092 6604 28144
rect 4620 27888 4672 27940
rect 3792 27820 3844 27872
rect 7104 28092 7156 28144
rect 8484 27956 8536 28008
rect 7564 27888 7616 27940
rect 9864 28024 9916 28076
rect 11152 28024 11204 28076
rect 11336 28024 11388 28076
rect 11704 28067 11756 28076
rect 11704 28033 11713 28067
rect 11713 28033 11747 28067
rect 11747 28033 11756 28067
rect 11704 28024 11756 28033
rect 11796 28024 11848 28076
rect 12624 28024 12676 28076
rect 12716 28024 12768 28076
rect 8852 27956 8904 28008
rect 9680 27888 9732 27940
rect 13360 28024 13412 28076
rect 13544 28067 13596 28076
rect 13544 28033 13553 28067
rect 13553 28033 13587 28067
rect 13587 28033 13596 28067
rect 13544 28024 13596 28033
rect 13912 28135 13964 28144
rect 13912 28101 13921 28135
rect 13921 28101 13955 28135
rect 13955 28101 13964 28135
rect 13912 28092 13964 28101
rect 14832 28160 14884 28212
rect 15016 28160 15068 28212
rect 15476 28160 15528 28212
rect 15752 28135 15804 28144
rect 15752 28101 15761 28135
rect 15761 28101 15795 28135
rect 15795 28101 15804 28135
rect 15752 28092 15804 28101
rect 16028 28092 16080 28144
rect 13820 28067 13872 28076
rect 13820 28033 13829 28067
rect 13829 28033 13863 28067
rect 13863 28033 13872 28067
rect 13820 28024 13872 28033
rect 14280 28024 14332 28076
rect 14372 27956 14424 28008
rect 13820 27888 13872 27940
rect 13912 27888 13964 27940
rect 14556 27956 14608 28008
rect 14740 28024 14792 28076
rect 15200 28024 15252 28076
rect 15016 27956 15068 28008
rect 14740 27888 14792 27940
rect 6920 27820 6972 27872
rect 7288 27820 7340 27872
rect 12532 27820 12584 27872
rect 14004 27820 14056 27872
rect 14280 27863 14332 27872
rect 14280 27829 14289 27863
rect 14289 27829 14323 27863
rect 14323 27829 14332 27863
rect 14280 27820 14332 27829
rect 14372 27820 14424 27872
rect 15752 27956 15804 28008
rect 16672 28067 16724 28076
rect 16672 28033 16681 28067
rect 16681 28033 16715 28067
rect 16715 28033 16724 28067
rect 16672 28024 16724 28033
rect 17500 28092 17552 28144
rect 17684 28024 17736 28076
rect 18144 27956 18196 28008
rect 18696 27956 18748 28008
rect 19432 28092 19484 28144
rect 19708 28024 19760 28076
rect 21456 28092 21508 28144
rect 19156 27956 19208 28008
rect 19248 27956 19300 28008
rect 19616 27956 19668 28008
rect 19524 27888 19576 27940
rect 16120 27820 16172 27872
rect 17316 27863 17368 27872
rect 17316 27829 17325 27863
rect 17325 27829 17359 27863
rect 17359 27829 17368 27863
rect 17316 27820 17368 27829
rect 17408 27820 17460 27872
rect 17868 27820 17920 27872
rect 19156 27820 19208 27872
rect 21640 28024 21692 28076
rect 21824 28067 21876 28076
rect 21824 28033 21833 28067
rect 21833 28033 21867 28067
rect 21867 28033 21876 28067
rect 21824 28024 21876 28033
rect 22100 28067 22152 28076
rect 22100 28033 22109 28067
rect 22109 28033 22143 28067
rect 22143 28033 22152 28067
rect 22100 28024 22152 28033
rect 20812 27999 20864 28008
rect 20812 27965 20821 27999
rect 20821 27965 20855 27999
rect 20855 27965 20864 27999
rect 20812 27956 20864 27965
rect 21456 27956 21508 28008
rect 25412 28203 25464 28212
rect 25412 28169 25421 28203
rect 25421 28169 25455 28203
rect 25455 28169 25464 28203
rect 25412 28160 25464 28169
rect 25504 28160 25556 28212
rect 32496 28203 32548 28212
rect 32496 28169 32505 28203
rect 32505 28169 32539 28203
rect 32539 28169 32548 28203
rect 32496 28160 32548 28169
rect 22468 28024 22520 28076
rect 22744 28024 22796 28076
rect 24768 28092 24820 28144
rect 30104 28092 30156 28144
rect 30840 28135 30892 28144
rect 30840 28101 30849 28135
rect 30849 28101 30883 28135
rect 30883 28101 30892 28135
rect 30840 28092 30892 28101
rect 31392 28135 31444 28144
rect 31392 28101 31401 28135
rect 31401 28101 31435 28135
rect 31435 28101 31444 28135
rect 31392 28092 31444 28101
rect 23020 28067 23072 28076
rect 23020 28033 23029 28067
rect 23029 28033 23063 28067
rect 23063 28033 23072 28067
rect 23020 28024 23072 28033
rect 26056 28024 26108 28076
rect 20352 27888 20404 27940
rect 21088 27888 21140 27940
rect 23664 27956 23716 28008
rect 23756 27956 23808 28008
rect 22744 27888 22796 27940
rect 25780 27956 25832 28008
rect 29184 27999 29236 28008
rect 29184 27965 29193 27999
rect 29193 27965 29227 27999
rect 29227 27965 29236 27999
rect 29184 27956 29236 27965
rect 30748 28024 30800 28076
rect 32404 28024 32456 28076
rect 32588 28024 32640 28076
rect 30196 27956 30248 28008
rect 30564 27956 30616 28008
rect 25872 27888 25924 27940
rect 20536 27820 20588 27872
rect 23296 27820 23348 27872
rect 24216 27820 24268 27872
rect 25136 27820 25188 27872
rect 29920 27820 29972 27872
rect 30104 27820 30156 27872
rect 30288 27820 30340 27872
rect 30656 27820 30708 27872
rect 31668 27956 31720 28008
rect 32772 27956 32824 28008
rect 31484 27888 31536 27940
rect 31944 27888 31996 27940
rect 37004 27888 37056 27940
rect 32128 27820 32180 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 8392 27616 8444 27668
rect 5540 27591 5592 27600
rect 5540 27557 5549 27591
rect 5549 27557 5583 27591
rect 5583 27557 5592 27591
rect 5540 27548 5592 27557
rect 6460 27548 6512 27600
rect 3792 27523 3844 27532
rect 3792 27489 3801 27523
rect 3801 27489 3835 27523
rect 3835 27489 3844 27523
rect 3792 27480 3844 27489
rect 6828 27480 6880 27532
rect 9588 27523 9640 27532
rect 9588 27489 9597 27523
rect 9597 27489 9631 27523
rect 9631 27489 9640 27523
rect 9588 27480 9640 27489
rect 11520 27616 11572 27668
rect 11796 27616 11848 27668
rect 12716 27616 12768 27668
rect 13820 27616 13872 27668
rect 14556 27616 14608 27668
rect 14740 27616 14792 27668
rect 15752 27616 15804 27668
rect 17684 27659 17736 27668
rect 17684 27625 17693 27659
rect 17693 27625 17727 27659
rect 17727 27625 17736 27659
rect 17684 27616 17736 27625
rect 17868 27659 17920 27668
rect 17868 27625 17877 27659
rect 17877 27625 17911 27659
rect 17911 27625 17920 27659
rect 17868 27616 17920 27625
rect 12992 27591 13044 27600
rect 12992 27557 13001 27591
rect 13001 27557 13035 27591
rect 13035 27557 13044 27591
rect 12992 27548 13044 27557
rect 13544 27548 13596 27600
rect 12256 27480 12308 27532
rect 9864 27412 9916 27464
rect 10692 27412 10744 27464
rect 10876 27412 10928 27464
rect 11152 27412 11204 27464
rect 13268 27455 13320 27464
rect 13268 27421 13277 27455
rect 13277 27421 13311 27455
rect 13311 27421 13320 27455
rect 13268 27412 13320 27421
rect 4068 27387 4120 27396
rect 4068 27353 4077 27387
rect 4077 27353 4111 27387
rect 4111 27353 4120 27387
rect 4068 27344 4120 27353
rect 7748 27344 7800 27396
rect 9772 27344 9824 27396
rect 13452 27455 13504 27464
rect 13452 27421 13461 27455
rect 13461 27421 13495 27455
rect 13495 27421 13504 27455
rect 13452 27412 13504 27421
rect 15200 27548 15252 27600
rect 16672 27548 16724 27600
rect 15016 27480 15068 27532
rect 14096 27344 14148 27396
rect 4344 27276 4396 27328
rect 11152 27276 11204 27328
rect 14556 27455 14608 27464
rect 14556 27421 14565 27455
rect 14565 27421 14599 27455
rect 14599 27421 14608 27455
rect 14556 27412 14608 27421
rect 14648 27455 14700 27464
rect 14648 27421 14657 27455
rect 14657 27421 14691 27455
rect 14691 27421 14700 27455
rect 14648 27412 14700 27421
rect 14740 27455 14792 27464
rect 14740 27421 14749 27455
rect 14749 27421 14783 27455
rect 14783 27421 14792 27455
rect 14740 27412 14792 27421
rect 14832 27344 14884 27396
rect 15476 27455 15528 27464
rect 15476 27421 15485 27455
rect 15485 27421 15519 27455
rect 15519 27421 15528 27455
rect 15476 27412 15528 27421
rect 15844 27480 15896 27532
rect 15936 27480 15988 27532
rect 19892 27548 19944 27600
rect 20904 27548 20956 27600
rect 24492 27548 24544 27600
rect 30380 27616 30432 27668
rect 31208 27616 31260 27668
rect 36084 27616 36136 27668
rect 37096 27616 37148 27668
rect 15752 27412 15804 27464
rect 17408 27412 17460 27464
rect 18512 27412 18564 27464
rect 18696 27455 18748 27464
rect 18696 27421 18705 27455
rect 18705 27421 18739 27455
rect 18739 27421 18748 27455
rect 18696 27412 18748 27421
rect 18788 27455 18840 27464
rect 18788 27421 18797 27455
rect 18797 27421 18831 27455
rect 18831 27421 18840 27455
rect 18788 27412 18840 27421
rect 17776 27344 17828 27396
rect 18236 27387 18288 27396
rect 18236 27353 18245 27387
rect 18245 27353 18279 27387
rect 18279 27353 18288 27387
rect 18236 27344 18288 27353
rect 18972 27455 19024 27464
rect 18972 27421 18981 27455
rect 18981 27421 19015 27455
rect 19015 27421 19024 27455
rect 20812 27480 20864 27532
rect 22836 27480 22888 27532
rect 23204 27480 23256 27532
rect 18972 27412 19024 27421
rect 19616 27412 19668 27464
rect 19708 27412 19760 27464
rect 20352 27412 20404 27464
rect 20628 27455 20680 27464
rect 20628 27421 20637 27455
rect 20637 27421 20671 27455
rect 20671 27421 20680 27455
rect 20628 27412 20680 27421
rect 27896 27480 27948 27532
rect 28172 27480 28224 27532
rect 19432 27344 19484 27396
rect 14372 27276 14424 27328
rect 14924 27276 14976 27328
rect 16028 27276 16080 27328
rect 16212 27276 16264 27328
rect 18052 27276 18104 27328
rect 19708 27319 19760 27328
rect 19708 27285 19717 27319
rect 19717 27285 19751 27319
rect 19751 27285 19760 27319
rect 19708 27276 19760 27285
rect 19892 27387 19944 27396
rect 19892 27353 19901 27387
rect 19901 27353 19935 27387
rect 19935 27353 19944 27387
rect 19892 27344 19944 27353
rect 24860 27344 24912 27396
rect 26516 27412 26568 27464
rect 27344 27412 27396 27464
rect 27712 27412 27764 27464
rect 28080 27412 28132 27464
rect 30748 27548 30800 27600
rect 30932 27591 30984 27600
rect 30932 27557 30941 27591
rect 30941 27557 30975 27591
rect 30975 27557 30984 27591
rect 30932 27548 30984 27557
rect 29736 27523 29788 27532
rect 29736 27489 29745 27523
rect 29745 27489 29779 27523
rect 29779 27489 29788 27523
rect 29736 27480 29788 27489
rect 30564 27480 30616 27532
rect 31024 27523 31076 27532
rect 31024 27489 31033 27523
rect 31033 27489 31067 27523
rect 31067 27489 31076 27523
rect 31024 27480 31076 27489
rect 28724 27412 28776 27464
rect 29644 27412 29696 27464
rect 31852 27548 31904 27600
rect 32312 27548 32364 27600
rect 32588 27548 32640 27600
rect 32128 27523 32180 27532
rect 32128 27489 32137 27523
rect 32137 27489 32171 27523
rect 32171 27489 32180 27523
rect 32128 27480 32180 27489
rect 32956 27480 33008 27532
rect 38660 27548 38712 27600
rect 34428 27480 34480 27532
rect 32588 27455 32640 27464
rect 32588 27421 32597 27455
rect 32597 27421 32631 27455
rect 32631 27421 32640 27455
rect 32588 27412 32640 27421
rect 32772 27412 32824 27464
rect 33140 27455 33192 27464
rect 33140 27421 33149 27455
rect 33149 27421 33183 27455
rect 33183 27421 33192 27455
rect 33140 27412 33192 27421
rect 25596 27344 25648 27396
rect 25780 27344 25832 27396
rect 20260 27319 20312 27328
rect 20260 27285 20269 27319
rect 20269 27285 20303 27319
rect 20303 27285 20312 27319
rect 20260 27276 20312 27285
rect 24308 27276 24360 27328
rect 24584 27276 24636 27328
rect 31208 27387 31260 27396
rect 31208 27353 31217 27387
rect 31217 27353 31251 27387
rect 31251 27353 31260 27387
rect 31208 27344 31260 27353
rect 31392 27344 31444 27396
rect 32128 27344 32180 27396
rect 32404 27387 32456 27396
rect 32404 27353 32413 27387
rect 32413 27353 32447 27387
rect 32447 27353 32456 27387
rect 32404 27344 32456 27353
rect 33784 27412 33836 27464
rect 37188 27480 37240 27532
rect 38108 27480 38160 27532
rect 36820 27455 36872 27464
rect 36820 27421 36829 27455
rect 36829 27421 36863 27455
rect 36863 27421 36872 27455
rect 36820 27412 36872 27421
rect 37372 27455 37424 27464
rect 37372 27421 37381 27455
rect 37381 27421 37415 27455
rect 37415 27421 37424 27455
rect 37372 27412 37424 27421
rect 38016 27412 38068 27464
rect 38844 27344 38896 27396
rect 39580 27387 39632 27396
rect 39580 27353 39589 27387
rect 39589 27353 39623 27387
rect 39623 27353 39632 27387
rect 39580 27344 39632 27353
rect 32772 27319 32824 27328
rect 32772 27285 32781 27319
rect 32781 27285 32815 27319
rect 32815 27285 32824 27319
rect 32772 27276 32824 27285
rect 32956 27276 33008 27328
rect 35992 27276 36044 27328
rect 36544 27276 36596 27328
rect 36912 27276 36964 27328
rect 37464 27276 37516 27328
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 4068 27072 4120 27124
rect 4344 27115 4396 27124
rect 4344 27081 4353 27115
rect 4353 27081 4387 27115
rect 4387 27081 4396 27115
rect 4344 27072 4396 27081
rect 5540 27072 5592 27124
rect 5908 27072 5960 27124
rect 6736 27072 6788 27124
rect 8392 27115 8444 27124
rect 8392 27081 8401 27115
rect 8401 27081 8435 27115
rect 8435 27081 8444 27115
rect 8392 27072 8444 27081
rect 9680 27072 9732 27124
rect 9772 27115 9824 27124
rect 9772 27081 9781 27115
rect 9781 27081 9815 27115
rect 9815 27081 9824 27115
rect 9772 27072 9824 27081
rect 10232 27115 10284 27124
rect 10232 27081 10241 27115
rect 10241 27081 10275 27115
rect 10275 27081 10284 27115
rect 10232 27072 10284 27081
rect 3148 27004 3200 27056
rect 6092 27004 6144 27056
rect 7288 27004 7340 27056
rect 7932 27004 7984 27056
rect 11060 27072 11112 27124
rect 11244 27072 11296 27124
rect 4620 26911 4672 26920
rect 4620 26877 4629 26911
rect 4629 26877 4663 26911
rect 4663 26877 4672 26911
rect 4620 26868 4672 26877
rect 5816 26979 5868 26988
rect 5816 26945 5825 26979
rect 5825 26945 5859 26979
rect 5859 26945 5868 26979
rect 5816 26936 5868 26945
rect 5908 26979 5960 26988
rect 5908 26945 5917 26979
rect 5917 26945 5951 26979
rect 5951 26945 5960 26979
rect 5908 26936 5960 26945
rect 6368 26936 6420 26988
rect 6828 26979 6880 26988
rect 6828 26945 6837 26979
rect 6837 26945 6871 26979
rect 6871 26945 6880 26979
rect 6828 26936 6880 26945
rect 8484 26868 8536 26920
rect 8760 26868 8812 26920
rect 10232 26936 10284 26988
rect 10692 27047 10744 27056
rect 10692 27013 10701 27047
rect 10701 27013 10735 27047
rect 10735 27013 10744 27047
rect 10692 27004 10744 27013
rect 10968 27004 11020 27056
rect 13728 27072 13780 27124
rect 14648 27072 14700 27124
rect 15108 27072 15160 27124
rect 15292 27072 15344 27124
rect 15844 27072 15896 27124
rect 16488 27072 16540 27124
rect 12440 27004 12492 27056
rect 9772 26868 9824 26920
rect 6276 26800 6328 26852
rect 9496 26800 9548 26852
rect 10140 26800 10192 26852
rect 10508 26979 10560 26988
rect 10508 26945 10517 26979
rect 10517 26945 10551 26979
rect 10551 26945 10560 26979
rect 10508 26936 10560 26945
rect 11520 26979 11572 26988
rect 11520 26945 11529 26979
rect 11529 26945 11563 26979
rect 11563 26945 11572 26979
rect 11520 26936 11572 26945
rect 13360 26979 13412 26988
rect 13360 26945 13369 26979
rect 13369 26945 13403 26979
rect 13403 26945 13412 26979
rect 13360 26936 13412 26945
rect 13820 26936 13872 26988
rect 14556 26936 14608 26988
rect 14924 26979 14976 26988
rect 14924 26945 14933 26979
rect 14933 26945 14967 26979
rect 14967 26945 14976 26979
rect 14924 26936 14976 26945
rect 15292 26979 15344 26988
rect 15292 26945 15301 26979
rect 15301 26945 15335 26979
rect 15335 26945 15344 26979
rect 15292 26936 15344 26945
rect 10600 26911 10652 26920
rect 10600 26877 10628 26911
rect 10628 26877 10652 26911
rect 10600 26868 10652 26877
rect 11152 26868 11204 26920
rect 11336 26868 11388 26920
rect 12532 26868 12584 26920
rect 13912 26868 13964 26920
rect 14740 26868 14792 26920
rect 14832 26911 14884 26920
rect 14832 26877 14841 26911
rect 14841 26877 14875 26911
rect 14875 26877 14884 26911
rect 14832 26868 14884 26877
rect 11980 26800 12032 26852
rect 6000 26732 6052 26784
rect 6460 26732 6512 26784
rect 9772 26732 9824 26784
rect 10600 26732 10652 26784
rect 11888 26732 11940 26784
rect 12072 26775 12124 26784
rect 12072 26741 12081 26775
rect 12081 26741 12115 26775
rect 12115 26741 12124 26775
rect 12072 26732 12124 26741
rect 13268 26800 13320 26852
rect 15108 26911 15160 26920
rect 15108 26877 15117 26911
rect 15117 26877 15151 26911
rect 15151 26877 15160 26911
rect 15108 26868 15160 26877
rect 14188 26732 14240 26784
rect 14924 26732 14976 26784
rect 16212 26936 16264 26988
rect 16764 26936 16816 26988
rect 16948 26979 17000 26988
rect 16948 26945 16957 26979
rect 16957 26945 16991 26979
rect 16991 26945 17000 26979
rect 16948 26936 17000 26945
rect 17224 26979 17276 26988
rect 16396 26868 16448 26920
rect 17224 26945 17232 26979
rect 17232 26945 17266 26979
rect 17266 26945 17276 26979
rect 17224 26936 17276 26945
rect 17316 26979 17368 26988
rect 17316 26945 17325 26979
rect 17325 26945 17359 26979
rect 17359 26945 17368 26979
rect 17316 26936 17368 26945
rect 17776 26936 17828 26988
rect 18052 26868 18104 26920
rect 18328 26979 18380 26988
rect 18328 26945 18337 26979
rect 18337 26945 18371 26979
rect 18371 26945 18380 26979
rect 18328 26936 18380 26945
rect 18696 27004 18748 27056
rect 18696 26868 18748 26920
rect 18788 26911 18840 26920
rect 18788 26877 18797 26911
rect 18797 26877 18831 26911
rect 18831 26877 18840 26911
rect 18788 26868 18840 26877
rect 19156 26979 19208 26988
rect 19156 26945 19165 26979
rect 19165 26945 19199 26979
rect 19199 26945 19208 26979
rect 19708 27072 19760 27124
rect 19892 27072 19944 27124
rect 20812 27115 20864 27124
rect 20812 27081 20821 27115
rect 20821 27081 20855 27115
rect 20855 27081 20864 27115
rect 20812 27072 20864 27081
rect 24124 27072 24176 27124
rect 19156 26936 19208 26945
rect 19248 26911 19300 26920
rect 19248 26877 19257 26911
rect 19257 26877 19291 26911
rect 19291 26877 19300 26911
rect 19248 26868 19300 26877
rect 19892 26936 19944 26988
rect 20076 26979 20128 26988
rect 20076 26945 20085 26979
rect 20085 26945 20119 26979
rect 20119 26945 20128 26979
rect 20076 26936 20128 26945
rect 20260 26936 20312 26988
rect 20628 26936 20680 26988
rect 21824 26936 21876 26988
rect 22192 26979 22244 26988
rect 22192 26945 22201 26979
rect 22201 26945 22235 26979
rect 22235 26945 22244 26979
rect 22192 26936 22244 26945
rect 21456 26868 21508 26920
rect 18604 26800 18656 26852
rect 22652 26979 22704 26988
rect 22652 26945 22661 26979
rect 22661 26945 22695 26979
rect 22695 26945 22704 26979
rect 22652 26936 22704 26945
rect 22744 26936 22796 26988
rect 25964 27072 26016 27124
rect 30012 27072 30064 27124
rect 25228 27004 25280 27056
rect 28632 27004 28684 27056
rect 31024 27072 31076 27124
rect 31116 27072 31168 27124
rect 31576 27072 31628 27124
rect 23296 26979 23348 26988
rect 23296 26945 23305 26979
rect 23305 26945 23339 26979
rect 23339 26945 23348 26979
rect 23296 26936 23348 26945
rect 24124 26936 24176 26988
rect 25320 26936 25372 26988
rect 20720 26732 20772 26784
rect 21364 26732 21416 26784
rect 22744 26775 22796 26784
rect 22744 26741 22753 26775
rect 22753 26741 22787 26775
rect 22787 26741 22796 26775
rect 22744 26732 22796 26741
rect 23480 26868 23532 26920
rect 24584 26868 24636 26920
rect 24676 26868 24728 26920
rect 23204 26800 23256 26852
rect 25780 26979 25832 26988
rect 25780 26945 25789 26979
rect 25789 26945 25823 26979
rect 25823 26945 25832 26979
rect 25780 26936 25832 26945
rect 26792 26936 26844 26988
rect 30748 26936 30800 26988
rect 32128 27047 32180 27056
rect 32128 27013 32137 27047
rect 32137 27013 32171 27047
rect 32171 27013 32180 27047
rect 32128 27004 32180 27013
rect 31760 26979 31812 26988
rect 31760 26945 31769 26979
rect 31769 26945 31803 26979
rect 31803 26945 31812 26979
rect 31760 26936 31812 26945
rect 31944 26936 31996 26988
rect 34428 26979 34480 26988
rect 34428 26945 34437 26979
rect 34437 26945 34471 26979
rect 34471 26945 34480 26979
rect 34428 26936 34480 26945
rect 36544 27072 36596 27124
rect 37832 27072 37884 27124
rect 38016 27072 38068 27124
rect 38752 27072 38804 27124
rect 37556 27047 37608 27056
rect 37556 27013 37565 27047
rect 37565 27013 37599 27047
rect 37599 27013 37608 27047
rect 37556 27004 37608 27013
rect 30012 26868 30064 26920
rect 29920 26800 29972 26852
rect 24216 26775 24268 26784
rect 24216 26741 24225 26775
rect 24225 26741 24259 26775
rect 24259 26741 24268 26775
rect 24216 26732 24268 26741
rect 32036 26868 32088 26920
rect 32588 26868 32640 26920
rect 36360 26868 36412 26920
rect 36820 26979 36872 26988
rect 36820 26945 36829 26979
rect 36829 26945 36863 26979
rect 36863 26945 36872 26979
rect 36820 26936 36872 26945
rect 37096 26936 37148 26988
rect 37464 26979 37516 26988
rect 37464 26945 37473 26979
rect 37473 26945 37507 26979
rect 37507 26945 37516 26979
rect 37464 26936 37516 26945
rect 37648 26979 37700 26988
rect 37648 26945 37657 26979
rect 37657 26945 37691 26979
rect 37691 26945 37700 26979
rect 37648 26936 37700 26945
rect 37740 26979 37792 26988
rect 37740 26945 37775 26979
rect 37775 26945 37792 26979
rect 37740 26936 37792 26945
rect 38384 26979 38436 26988
rect 38384 26945 38393 26979
rect 38393 26945 38427 26979
rect 38427 26945 38436 26979
rect 38384 26936 38436 26945
rect 38660 26979 38712 26988
rect 38660 26945 38669 26979
rect 38669 26945 38703 26979
rect 38703 26945 38712 26979
rect 38660 26936 38712 26945
rect 38936 26979 38988 26988
rect 38936 26945 38945 26979
rect 38945 26945 38979 26979
rect 38979 26945 38988 26979
rect 38936 26936 38988 26945
rect 34060 26800 34112 26852
rect 35532 26800 35584 26852
rect 38752 26911 38804 26920
rect 38752 26877 38761 26911
rect 38761 26877 38795 26911
rect 38795 26877 38804 26911
rect 38752 26868 38804 26877
rect 38844 26911 38896 26920
rect 38844 26877 38853 26911
rect 38853 26877 38887 26911
rect 38887 26877 38896 26911
rect 38844 26868 38896 26877
rect 38016 26800 38068 26852
rect 38292 26800 38344 26852
rect 39304 27004 39356 27056
rect 39764 26936 39816 26988
rect 40224 26979 40276 26988
rect 40224 26945 40233 26979
rect 40233 26945 40267 26979
rect 40267 26945 40276 26979
rect 40224 26936 40276 26945
rect 39856 26800 39908 26852
rect 32312 26775 32364 26784
rect 32312 26741 32321 26775
rect 32321 26741 32355 26775
rect 32355 26741 32364 26775
rect 32312 26732 32364 26741
rect 34428 26732 34480 26784
rect 35348 26732 35400 26784
rect 37372 26732 37424 26784
rect 38844 26732 38896 26784
rect 39212 26732 39264 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 3056 26528 3108 26580
rect 5264 26528 5316 26580
rect 5356 26528 5408 26580
rect 6460 26528 6512 26580
rect 6828 26528 6880 26580
rect 9312 26528 9364 26580
rect 2780 26392 2832 26444
rect 3148 26435 3200 26444
rect 3148 26401 3157 26435
rect 3157 26401 3191 26435
rect 3191 26401 3200 26435
rect 3148 26392 3200 26401
rect 5264 26392 5316 26444
rect 4344 26367 4396 26376
rect 4344 26333 4353 26367
rect 4353 26333 4387 26367
rect 4387 26333 4396 26367
rect 4344 26324 4396 26333
rect 7012 26460 7064 26512
rect 8944 26503 8996 26512
rect 8944 26469 8953 26503
rect 8953 26469 8987 26503
rect 8987 26469 8996 26503
rect 8944 26460 8996 26469
rect 6368 26392 6420 26444
rect 6644 26392 6696 26444
rect 10508 26528 10560 26580
rect 10600 26571 10652 26580
rect 10600 26537 10609 26571
rect 10609 26537 10643 26571
rect 10643 26537 10652 26571
rect 10600 26528 10652 26537
rect 10784 26528 10836 26580
rect 10232 26460 10284 26512
rect 10876 26460 10928 26512
rect 12072 26571 12124 26580
rect 12072 26537 12081 26571
rect 12081 26537 12115 26571
rect 12115 26537 12124 26571
rect 12072 26528 12124 26537
rect 12256 26571 12308 26580
rect 12256 26537 12265 26571
rect 12265 26537 12299 26571
rect 12299 26537 12308 26571
rect 12256 26528 12308 26537
rect 12624 26571 12676 26580
rect 12624 26537 12633 26571
rect 12633 26537 12667 26571
rect 12667 26537 12676 26571
rect 12624 26528 12676 26537
rect 6000 26367 6052 26376
rect 6000 26333 6009 26367
rect 6009 26333 6043 26367
rect 6043 26333 6052 26367
rect 6000 26324 6052 26333
rect 6092 26367 6144 26376
rect 6092 26333 6102 26367
rect 6102 26333 6136 26367
rect 6136 26333 6144 26367
rect 6092 26324 6144 26333
rect 6828 26324 6880 26376
rect 7288 26324 7340 26376
rect 8024 26367 8076 26376
rect 8024 26333 8033 26367
rect 8033 26333 8067 26367
rect 8067 26333 8076 26367
rect 8024 26324 8076 26333
rect 9496 26392 9548 26444
rect 8392 26367 8444 26376
rect 8392 26333 8401 26367
rect 8401 26333 8435 26367
rect 8435 26333 8444 26367
rect 8392 26324 8444 26333
rect 8484 26324 8536 26376
rect 1860 26188 1912 26240
rect 5632 26299 5684 26308
rect 5632 26265 5641 26299
rect 5641 26265 5675 26299
rect 5675 26265 5684 26299
rect 5632 26256 5684 26265
rect 6276 26299 6328 26308
rect 6276 26265 6285 26299
rect 6285 26265 6319 26299
rect 6319 26265 6328 26299
rect 6276 26256 6328 26265
rect 6736 26256 6788 26308
rect 7104 26299 7156 26308
rect 7104 26265 7113 26299
rect 7113 26265 7147 26299
rect 7147 26265 7156 26299
rect 7104 26256 7156 26265
rect 9036 26256 9088 26308
rect 9312 26367 9364 26376
rect 9312 26333 9321 26367
rect 9321 26333 9355 26367
rect 9355 26333 9364 26367
rect 9312 26324 9364 26333
rect 10968 26392 11020 26444
rect 9496 26256 9548 26308
rect 10324 26324 10376 26376
rect 11152 26324 11204 26376
rect 11704 26460 11756 26512
rect 14280 26528 14332 26580
rect 14556 26528 14608 26580
rect 14832 26528 14884 26580
rect 18328 26528 18380 26580
rect 18696 26528 18748 26580
rect 19156 26528 19208 26580
rect 20076 26528 20128 26580
rect 22468 26571 22520 26580
rect 22468 26537 22477 26571
rect 22477 26537 22511 26571
rect 22511 26537 22520 26571
rect 22468 26528 22520 26537
rect 22652 26528 22704 26580
rect 22928 26528 22980 26580
rect 24032 26528 24084 26580
rect 14096 26503 14148 26512
rect 14096 26469 14105 26503
rect 14105 26469 14139 26503
rect 14139 26469 14148 26503
rect 14096 26460 14148 26469
rect 11336 26392 11388 26444
rect 10048 26256 10100 26308
rect 11060 26256 11112 26308
rect 11980 26256 12032 26308
rect 12164 26324 12216 26376
rect 12440 26367 12492 26376
rect 12440 26333 12449 26367
rect 12449 26333 12483 26367
rect 12483 26333 12492 26367
rect 12440 26324 12492 26333
rect 14372 26392 14424 26444
rect 15476 26460 15528 26512
rect 14648 26367 14700 26376
rect 12624 26256 12676 26308
rect 14648 26333 14656 26367
rect 14656 26333 14690 26367
rect 14690 26333 14700 26367
rect 14648 26324 14700 26333
rect 14740 26367 14792 26376
rect 14740 26333 14749 26367
rect 14749 26333 14783 26367
rect 14783 26333 14792 26367
rect 14740 26324 14792 26333
rect 14832 26256 14884 26308
rect 15844 26367 15896 26376
rect 15844 26333 15889 26367
rect 15889 26333 15896 26367
rect 15844 26324 15896 26333
rect 16028 26367 16080 26376
rect 16028 26333 16037 26367
rect 16037 26333 16071 26367
rect 16071 26333 16080 26367
rect 16028 26324 16080 26333
rect 16120 26367 16172 26376
rect 16120 26333 16129 26367
rect 16129 26333 16163 26367
rect 16163 26333 16172 26367
rect 16120 26324 16172 26333
rect 16304 26367 16356 26376
rect 16304 26333 16311 26367
rect 16311 26333 16356 26367
rect 16304 26324 16356 26333
rect 16396 26367 16448 26376
rect 16396 26333 16405 26367
rect 16405 26333 16439 26367
rect 16439 26333 16448 26367
rect 16396 26324 16448 26333
rect 16764 26324 16816 26376
rect 5816 26188 5868 26240
rect 8208 26188 8260 26240
rect 9772 26188 9824 26240
rect 14280 26188 14332 26240
rect 15660 26299 15712 26308
rect 15660 26265 15669 26299
rect 15669 26265 15703 26299
rect 15703 26265 15712 26299
rect 15660 26256 15712 26265
rect 15384 26231 15436 26240
rect 15384 26197 15393 26231
rect 15393 26197 15427 26231
rect 15427 26197 15436 26231
rect 15384 26188 15436 26197
rect 15476 26188 15528 26240
rect 16212 26188 16264 26240
rect 16856 26299 16908 26308
rect 16856 26265 16865 26299
rect 16865 26265 16899 26299
rect 16899 26265 16908 26299
rect 16856 26256 16908 26265
rect 16764 26231 16816 26240
rect 16764 26197 16773 26231
rect 16773 26197 16807 26231
rect 16807 26197 16816 26231
rect 16764 26188 16816 26197
rect 17132 26299 17184 26308
rect 17132 26265 17141 26299
rect 17141 26265 17175 26299
rect 17175 26265 17184 26299
rect 17132 26256 17184 26265
rect 18052 26324 18104 26376
rect 18144 26367 18196 26376
rect 18144 26333 18153 26367
rect 18153 26333 18187 26367
rect 18187 26333 18196 26367
rect 18144 26324 18196 26333
rect 18236 26324 18288 26376
rect 24676 26528 24728 26580
rect 20444 26392 20496 26444
rect 22836 26392 22888 26444
rect 25044 26528 25096 26580
rect 25136 26460 25188 26512
rect 25228 26460 25280 26512
rect 25504 26503 25556 26512
rect 25504 26469 25513 26503
rect 25513 26469 25547 26503
rect 25547 26469 25556 26503
rect 25504 26460 25556 26469
rect 25872 26528 25924 26580
rect 26792 26571 26844 26580
rect 26792 26537 26801 26571
rect 26801 26537 26835 26571
rect 26835 26537 26844 26571
rect 26792 26528 26844 26537
rect 19340 26324 19392 26376
rect 20352 26324 20404 26376
rect 17868 26299 17920 26308
rect 17868 26265 17877 26299
rect 17877 26265 17911 26299
rect 17911 26265 17920 26299
rect 17868 26256 17920 26265
rect 21364 26324 21416 26376
rect 22192 26367 22244 26376
rect 22192 26333 22201 26367
rect 22201 26333 22235 26367
rect 22235 26333 22244 26367
rect 22192 26324 22244 26333
rect 22376 26367 22428 26376
rect 22376 26333 22385 26367
rect 22385 26333 22419 26367
rect 22419 26333 22428 26367
rect 22376 26324 22428 26333
rect 26700 26435 26752 26444
rect 26700 26401 26709 26435
rect 26709 26401 26743 26435
rect 26743 26401 26752 26435
rect 26700 26392 26752 26401
rect 17316 26188 17368 26240
rect 18696 26188 18748 26240
rect 20812 26188 20864 26240
rect 23388 26256 23440 26308
rect 23572 26367 23624 26376
rect 23572 26333 23581 26367
rect 23581 26333 23615 26367
rect 23615 26333 23624 26367
rect 23572 26324 23624 26333
rect 24216 26324 24268 26376
rect 24492 26324 24544 26376
rect 24676 26367 24728 26376
rect 24676 26333 24685 26367
rect 24685 26333 24719 26367
rect 24719 26333 24728 26367
rect 24676 26324 24728 26333
rect 24768 26324 24820 26376
rect 25504 26324 25556 26376
rect 25044 26256 25096 26308
rect 25688 26299 25740 26308
rect 25688 26265 25715 26299
rect 25715 26265 25740 26299
rect 25688 26256 25740 26265
rect 26056 26256 26108 26308
rect 27068 26324 27120 26376
rect 29736 26571 29788 26580
rect 29736 26537 29745 26571
rect 29745 26537 29779 26571
rect 29779 26537 29788 26571
rect 29736 26528 29788 26537
rect 27988 26460 28040 26512
rect 28540 26460 28592 26512
rect 27620 26435 27672 26444
rect 27620 26401 27629 26435
rect 27629 26401 27663 26435
rect 27663 26401 27672 26435
rect 27620 26392 27672 26401
rect 28172 26392 28224 26444
rect 29276 26392 29328 26444
rect 31760 26528 31812 26580
rect 34520 26571 34572 26580
rect 34520 26537 34529 26571
rect 34529 26537 34563 26571
rect 34563 26537 34572 26571
rect 34520 26528 34572 26537
rect 27712 26324 27764 26376
rect 27804 26367 27856 26376
rect 27804 26333 27813 26367
rect 27813 26333 27847 26367
rect 27847 26333 27856 26367
rect 27804 26324 27856 26333
rect 27896 26367 27948 26376
rect 27896 26333 27905 26367
rect 27905 26333 27939 26367
rect 27939 26333 27948 26367
rect 27896 26324 27948 26333
rect 27988 26367 28040 26376
rect 27988 26333 27997 26367
rect 27997 26333 28031 26367
rect 28031 26333 28040 26367
rect 27988 26324 28040 26333
rect 22836 26231 22888 26240
rect 22836 26197 22845 26231
rect 22845 26197 22879 26231
rect 22879 26197 22888 26231
rect 22836 26188 22888 26197
rect 23112 26188 23164 26240
rect 24032 26188 24084 26240
rect 24400 26188 24452 26240
rect 24584 26188 24636 26240
rect 28264 26188 28316 26240
rect 28448 26367 28500 26376
rect 28448 26333 28457 26367
rect 28457 26333 28491 26367
rect 28491 26333 28500 26367
rect 28448 26324 28500 26333
rect 28816 26367 28868 26376
rect 28816 26333 28825 26367
rect 28825 26333 28859 26367
rect 28859 26333 28868 26367
rect 28816 26324 28868 26333
rect 29920 26367 29972 26376
rect 29920 26333 29929 26367
rect 29929 26333 29963 26367
rect 29963 26333 29972 26367
rect 29920 26324 29972 26333
rect 30748 26324 30800 26376
rect 32496 26460 32548 26512
rect 33600 26460 33652 26512
rect 33876 26460 33928 26512
rect 31944 26392 31996 26444
rect 31392 26367 31444 26376
rect 31392 26333 31401 26367
rect 31401 26333 31435 26367
rect 31435 26333 31444 26367
rect 31392 26324 31444 26333
rect 31576 26367 31628 26376
rect 31576 26333 31585 26367
rect 31585 26333 31619 26367
rect 31619 26333 31628 26367
rect 31576 26324 31628 26333
rect 31852 26367 31904 26376
rect 31852 26333 31861 26367
rect 31861 26333 31895 26367
rect 31895 26333 31904 26367
rect 31852 26324 31904 26333
rect 32036 26324 32088 26376
rect 32404 26324 32456 26376
rect 32496 26367 32548 26376
rect 32496 26333 32505 26367
rect 32505 26333 32539 26367
rect 32539 26333 32548 26367
rect 32496 26324 32548 26333
rect 32588 26367 32640 26376
rect 32588 26333 32597 26367
rect 32597 26333 32631 26367
rect 32631 26333 32640 26367
rect 32588 26324 32640 26333
rect 33508 26324 33560 26376
rect 33876 26324 33928 26376
rect 34428 26324 34480 26376
rect 35348 26460 35400 26512
rect 36360 26528 36412 26580
rect 38384 26528 38436 26580
rect 37556 26460 37608 26512
rect 38476 26460 38528 26512
rect 38936 26460 38988 26512
rect 39304 26460 39356 26512
rect 37096 26392 37148 26444
rect 37280 26392 37332 26444
rect 38108 26435 38160 26444
rect 38108 26401 38117 26435
rect 38117 26401 38151 26435
rect 38151 26401 38160 26435
rect 38108 26392 38160 26401
rect 28632 26256 28684 26308
rect 29736 26256 29788 26308
rect 31208 26299 31260 26308
rect 31208 26265 31217 26299
rect 31217 26265 31251 26299
rect 31251 26265 31260 26299
rect 31208 26256 31260 26265
rect 31116 26188 31168 26240
rect 32772 26299 32824 26308
rect 32772 26265 32781 26299
rect 32781 26265 32815 26299
rect 32815 26265 32824 26299
rect 35532 26324 35584 26376
rect 37740 26324 37792 26376
rect 37832 26324 37884 26376
rect 32772 26256 32824 26265
rect 35624 26299 35676 26308
rect 35624 26265 35633 26299
rect 35633 26265 35667 26299
rect 35667 26265 35676 26299
rect 35624 26256 35676 26265
rect 35992 26256 36044 26308
rect 39764 26324 39816 26376
rect 39948 26324 40000 26376
rect 38384 26299 38436 26308
rect 38384 26265 38393 26299
rect 38393 26265 38427 26299
rect 38427 26265 38436 26299
rect 38384 26256 38436 26265
rect 31852 26231 31904 26240
rect 31852 26197 31861 26231
rect 31861 26197 31895 26231
rect 31895 26197 31904 26231
rect 31852 26188 31904 26197
rect 33140 26188 33192 26240
rect 34888 26188 34940 26240
rect 35072 26188 35124 26240
rect 36544 26188 36596 26240
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 4344 25984 4396 26036
rect 5356 25984 5408 26036
rect 5632 25984 5684 26036
rect 7104 25984 7156 26036
rect 9220 25984 9272 26036
rect 11888 25984 11940 26036
rect 12256 25984 12308 26036
rect 1860 25959 1912 25968
rect 1860 25925 1869 25959
rect 1869 25925 1903 25959
rect 1903 25925 1912 25959
rect 1860 25916 1912 25925
rect 3148 25916 3200 25968
rect 3976 25916 4028 25968
rect 4436 25916 4488 25968
rect 3700 25891 3752 25900
rect 3700 25857 3709 25891
rect 3709 25857 3743 25891
rect 3743 25857 3752 25891
rect 3700 25848 3752 25857
rect 6276 25916 6328 25968
rect 16764 25984 16816 26036
rect 18880 25984 18932 26036
rect 24216 25984 24268 26036
rect 25596 25984 25648 26036
rect 25780 25984 25832 26036
rect 28264 25984 28316 26036
rect 29368 25984 29420 26036
rect 30840 25984 30892 26036
rect 6368 25891 6420 25900
rect 6368 25857 6377 25891
rect 6377 25857 6411 25891
rect 6411 25857 6420 25891
rect 6368 25848 6420 25857
rect 6552 25891 6604 25900
rect 6552 25857 6559 25891
rect 6559 25857 6604 25891
rect 6552 25848 6604 25857
rect 1584 25823 1636 25832
rect 1584 25789 1593 25823
rect 1593 25789 1627 25823
rect 1627 25789 1636 25823
rect 1584 25780 1636 25789
rect 3976 25823 4028 25832
rect 3976 25789 3985 25823
rect 3985 25789 4019 25823
rect 4019 25789 4028 25823
rect 3976 25780 4028 25789
rect 6552 25712 6604 25764
rect 15384 25916 15436 25968
rect 6828 25848 6880 25900
rect 7012 25848 7064 25900
rect 7196 25891 7248 25900
rect 7196 25857 7206 25891
rect 7206 25857 7240 25891
rect 7240 25857 7248 25891
rect 7196 25848 7248 25857
rect 7472 25891 7524 25900
rect 7472 25857 7481 25891
rect 7481 25857 7515 25891
rect 7515 25857 7524 25891
rect 7472 25848 7524 25857
rect 8484 25848 8536 25900
rect 10048 25891 10100 25900
rect 10048 25857 10057 25891
rect 10057 25857 10091 25891
rect 10091 25857 10100 25891
rect 10048 25848 10100 25857
rect 11704 25891 11756 25900
rect 11704 25857 11713 25891
rect 11713 25857 11747 25891
rect 11747 25857 11756 25891
rect 11704 25848 11756 25857
rect 11888 25891 11940 25900
rect 11888 25857 11897 25891
rect 11897 25857 11931 25891
rect 11931 25857 11940 25891
rect 11888 25848 11940 25857
rect 11980 25848 12032 25900
rect 12440 25891 12492 25900
rect 12440 25857 12449 25891
rect 12449 25857 12483 25891
rect 12483 25857 12492 25891
rect 12440 25848 12492 25857
rect 13084 25848 13136 25900
rect 13360 25891 13412 25900
rect 13360 25857 13369 25891
rect 13369 25857 13403 25891
rect 13403 25857 13412 25891
rect 13360 25848 13412 25857
rect 12532 25780 12584 25832
rect 13636 25891 13688 25900
rect 13636 25857 13645 25891
rect 13645 25857 13679 25891
rect 13679 25857 13688 25891
rect 13636 25848 13688 25857
rect 13820 25891 13872 25900
rect 13820 25857 13829 25891
rect 13829 25857 13863 25891
rect 13863 25857 13872 25891
rect 13820 25848 13872 25857
rect 13912 25891 13964 25900
rect 13912 25857 13921 25891
rect 13921 25857 13955 25891
rect 13955 25857 13964 25891
rect 13912 25848 13964 25857
rect 14004 25891 14056 25900
rect 14004 25857 14013 25891
rect 14013 25857 14047 25891
rect 14047 25857 14056 25891
rect 14004 25848 14056 25857
rect 14096 25848 14148 25900
rect 14556 25891 14608 25900
rect 14556 25857 14565 25891
rect 14565 25857 14599 25891
rect 14599 25857 14608 25891
rect 14556 25848 14608 25857
rect 14924 25848 14976 25900
rect 18236 25848 18288 25900
rect 18328 25848 18380 25900
rect 19064 25891 19116 25900
rect 19064 25857 19073 25891
rect 19073 25857 19107 25891
rect 19107 25857 19116 25891
rect 19064 25848 19116 25857
rect 19340 25916 19392 25968
rect 24676 25848 24728 25900
rect 13728 25712 13780 25764
rect 15108 25780 15160 25832
rect 16028 25780 16080 25832
rect 17684 25780 17736 25832
rect 23204 25780 23256 25832
rect 26056 25848 26108 25900
rect 28540 25916 28592 25968
rect 33968 25984 34020 26036
rect 29276 25891 29328 25900
rect 29276 25857 29285 25891
rect 29285 25857 29319 25891
rect 29319 25857 29328 25891
rect 29276 25848 29328 25857
rect 29368 25891 29420 25900
rect 29368 25857 29377 25891
rect 29377 25857 29411 25891
rect 29411 25857 29420 25891
rect 29368 25848 29420 25857
rect 29552 25848 29604 25900
rect 31116 25916 31168 25968
rect 31300 25916 31352 25968
rect 31392 25916 31444 25968
rect 36084 25984 36136 26036
rect 38016 25984 38068 26036
rect 30932 25891 30984 25900
rect 30932 25857 30941 25891
rect 30941 25857 30975 25891
rect 30975 25857 30984 25891
rect 30932 25848 30984 25857
rect 31576 25848 31628 25900
rect 32496 25891 32548 25900
rect 32496 25857 32505 25891
rect 32505 25857 32539 25891
rect 32539 25857 32548 25891
rect 32496 25848 32548 25857
rect 33876 25891 33928 25900
rect 33876 25857 33885 25891
rect 33885 25857 33919 25891
rect 33919 25857 33928 25891
rect 33876 25848 33928 25857
rect 34336 25848 34388 25900
rect 34428 25891 34480 25900
rect 34428 25857 34437 25891
rect 34437 25857 34471 25891
rect 34471 25857 34480 25891
rect 34428 25848 34480 25857
rect 34520 25848 34572 25900
rect 34888 25891 34940 25900
rect 34888 25857 34897 25891
rect 34897 25857 34931 25891
rect 34931 25857 34940 25891
rect 34888 25848 34940 25857
rect 35348 25916 35400 25968
rect 36176 25916 36228 25968
rect 36728 25916 36780 25968
rect 35072 25891 35124 25900
rect 35072 25857 35081 25891
rect 35081 25857 35115 25891
rect 35115 25857 35124 25891
rect 35072 25848 35124 25857
rect 37648 25848 37700 25900
rect 15200 25712 15252 25764
rect 18144 25712 18196 25764
rect 26148 25712 26200 25764
rect 27988 25712 28040 25764
rect 35164 25780 35216 25832
rect 35992 25780 36044 25832
rect 37004 25780 37056 25832
rect 38476 25891 38528 25900
rect 38476 25857 38485 25891
rect 38485 25857 38519 25891
rect 38519 25857 38528 25891
rect 38476 25848 38528 25857
rect 34428 25755 34480 25764
rect 34428 25721 34437 25755
rect 34437 25721 34471 25755
rect 34471 25721 34480 25755
rect 34428 25712 34480 25721
rect 38752 25780 38804 25832
rect 5540 25687 5592 25696
rect 5540 25653 5549 25687
rect 5549 25653 5583 25687
rect 5583 25653 5592 25687
rect 5540 25644 5592 25653
rect 7012 25687 7064 25696
rect 7012 25653 7021 25687
rect 7021 25653 7055 25687
rect 7055 25653 7064 25687
rect 7012 25644 7064 25653
rect 10324 25687 10376 25696
rect 10324 25653 10333 25687
rect 10333 25653 10367 25687
rect 10367 25653 10376 25687
rect 10324 25644 10376 25653
rect 12164 25644 12216 25696
rect 14464 25644 14516 25696
rect 16856 25644 16908 25696
rect 23572 25644 23624 25696
rect 29000 25687 29052 25696
rect 29000 25653 29009 25687
rect 29009 25653 29043 25687
rect 29043 25653 29052 25687
rect 29000 25644 29052 25653
rect 30748 25687 30800 25696
rect 30748 25653 30757 25687
rect 30757 25653 30791 25687
rect 30791 25653 30800 25687
rect 30748 25644 30800 25653
rect 31944 25644 31996 25696
rect 32128 25644 32180 25696
rect 34704 25644 34756 25696
rect 35808 25644 35860 25696
rect 36360 25644 36412 25696
rect 38016 25644 38068 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 3976 25440 4028 25492
rect 6368 25483 6420 25492
rect 6368 25449 6377 25483
rect 6377 25449 6411 25483
rect 6411 25449 6420 25483
rect 6368 25440 6420 25449
rect 6920 25440 6972 25492
rect 8116 25440 8168 25492
rect 11336 25440 11388 25492
rect 13360 25440 13412 25492
rect 15108 25440 15160 25492
rect 15660 25440 15712 25492
rect 7472 25372 7524 25424
rect 17868 25440 17920 25492
rect 20628 25440 20680 25492
rect 22284 25440 22336 25492
rect 24768 25440 24820 25492
rect 24860 25483 24912 25492
rect 24860 25449 24869 25483
rect 24869 25449 24903 25483
rect 24903 25449 24912 25483
rect 24860 25440 24912 25449
rect 25228 25440 25280 25492
rect 17408 25372 17460 25424
rect 1584 25347 1636 25356
rect 1584 25313 1593 25347
rect 1593 25313 1627 25347
rect 1627 25313 1636 25347
rect 1584 25304 1636 25313
rect 2872 25304 2924 25356
rect 3700 25304 3752 25356
rect 4804 25304 4856 25356
rect 5264 25304 5316 25356
rect 5356 25304 5408 25356
rect 1860 25211 1912 25220
rect 1860 25177 1869 25211
rect 1869 25177 1903 25211
rect 1903 25177 1912 25211
rect 1860 25168 1912 25177
rect 3148 25168 3200 25220
rect 5540 25236 5592 25288
rect 5632 25236 5684 25288
rect 6184 25236 6236 25288
rect 6276 25236 6328 25288
rect 6460 25236 6512 25288
rect 7932 25304 7984 25356
rect 8484 25347 8536 25356
rect 8484 25313 8493 25347
rect 8493 25313 8527 25347
rect 8527 25313 8536 25347
rect 8484 25304 8536 25313
rect 9128 25304 9180 25356
rect 13728 25304 13780 25356
rect 7012 25279 7064 25288
rect 7012 25245 7021 25279
rect 7021 25245 7055 25279
rect 7055 25245 7064 25279
rect 7012 25236 7064 25245
rect 5816 25168 5868 25220
rect 3792 25143 3844 25152
rect 3792 25109 3801 25143
rect 3801 25109 3835 25143
rect 3835 25109 3844 25143
rect 3792 25100 3844 25109
rect 5540 25100 5592 25152
rect 7104 25168 7156 25220
rect 7288 25236 7340 25288
rect 8300 25236 8352 25288
rect 9036 25236 9088 25288
rect 9404 25236 9456 25288
rect 11060 25236 11112 25288
rect 11244 25236 11296 25288
rect 6460 25100 6512 25152
rect 7564 25100 7616 25152
rect 11980 25236 12032 25288
rect 15844 25304 15896 25356
rect 19064 25304 19116 25356
rect 8392 25143 8444 25152
rect 8392 25109 8401 25143
rect 8401 25109 8435 25143
rect 8435 25109 8444 25143
rect 8392 25100 8444 25109
rect 9772 25100 9824 25152
rect 11244 25143 11296 25152
rect 11244 25109 11271 25143
rect 11271 25109 11296 25143
rect 11244 25100 11296 25109
rect 14556 25168 14608 25220
rect 16304 25236 16356 25288
rect 16396 25236 16448 25288
rect 17316 25168 17368 25220
rect 15476 25143 15528 25152
rect 15476 25109 15503 25143
rect 15503 25109 15528 25143
rect 15476 25100 15528 25109
rect 16304 25100 16356 25152
rect 17132 25100 17184 25152
rect 18144 25100 18196 25152
rect 20812 25304 20864 25356
rect 21456 25304 21508 25356
rect 23020 25304 23072 25356
rect 23664 25304 23716 25356
rect 24400 25304 24452 25356
rect 25412 25304 25464 25356
rect 28448 25372 28500 25424
rect 20260 25279 20312 25288
rect 20260 25245 20269 25279
rect 20269 25245 20303 25279
rect 20303 25245 20312 25279
rect 20260 25236 20312 25245
rect 21088 25236 21140 25288
rect 18604 25168 18656 25220
rect 23112 25168 23164 25220
rect 23572 25279 23624 25288
rect 23572 25245 23581 25279
rect 23581 25245 23615 25279
rect 23615 25245 23624 25279
rect 23572 25236 23624 25245
rect 24216 25168 24268 25220
rect 22744 25100 22796 25152
rect 24584 25236 24636 25288
rect 25688 25236 25740 25288
rect 25872 25279 25924 25288
rect 25872 25245 25881 25279
rect 25881 25245 25915 25279
rect 25915 25245 25924 25279
rect 25872 25236 25924 25245
rect 24492 25168 24544 25220
rect 26976 25304 27028 25356
rect 26056 25236 26108 25288
rect 26240 25279 26292 25288
rect 26240 25245 26249 25279
rect 26249 25245 26283 25279
rect 26283 25245 26292 25279
rect 26240 25236 26292 25245
rect 26700 25279 26752 25288
rect 26700 25245 26709 25279
rect 26709 25245 26743 25279
rect 26743 25245 26752 25279
rect 26700 25236 26752 25245
rect 26884 25236 26936 25288
rect 30656 25440 30708 25492
rect 31944 25440 31996 25492
rect 35808 25440 35860 25492
rect 29000 25304 29052 25356
rect 30932 25347 30984 25356
rect 30932 25313 30941 25347
rect 30941 25313 30975 25347
rect 30975 25313 30984 25347
rect 30932 25304 30984 25313
rect 30748 25236 30800 25288
rect 31760 25236 31812 25288
rect 31852 25279 31904 25288
rect 31852 25245 31861 25279
rect 31861 25245 31895 25279
rect 31895 25245 31904 25279
rect 31852 25236 31904 25245
rect 32128 25279 32180 25288
rect 32128 25245 32137 25279
rect 32137 25245 32171 25279
rect 32171 25245 32180 25279
rect 32128 25236 32180 25245
rect 32864 25304 32916 25356
rect 33048 25279 33100 25288
rect 33048 25245 33057 25279
rect 33057 25245 33091 25279
rect 33091 25245 33100 25279
rect 33048 25236 33100 25245
rect 33600 25372 33652 25424
rect 37096 25372 37148 25424
rect 34336 25304 34388 25356
rect 33324 25279 33376 25288
rect 33324 25245 33333 25279
rect 33333 25245 33367 25279
rect 33367 25245 33376 25279
rect 33324 25236 33376 25245
rect 33692 25279 33744 25288
rect 33692 25245 33701 25279
rect 33701 25245 33735 25279
rect 33735 25245 33744 25279
rect 33692 25236 33744 25245
rect 35532 25279 35584 25288
rect 35532 25245 35541 25279
rect 35541 25245 35575 25279
rect 35575 25245 35584 25279
rect 35532 25236 35584 25245
rect 36084 25279 36136 25288
rect 36084 25245 36093 25279
rect 36093 25245 36127 25279
rect 36127 25245 36136 25279
rect 36084 25236 36136 25245
rect 26424 25100 26476 25152
rect 31024 25100 31076 25152
rect 32128 25100 32180 25152
rect 32404 25143 32456 25152
rect 32404 25109 32413 25143
rect 32413 25109 32447 25143
rect 32447 25109 32456 25143
rect 32404 25100 32456 25109
rect 32588 25143 32640 25152
rect 32588 25109 32597 25143
rect 32597 25109 32631 25143
rect 32631 25109 32640 25143
rect 32588 25100 32640 25109
rect 33600 25143 33652 25152
rect 33600 25109 33609 25143
rect 33609 25109 33643 25143
rect 33643 25109 33652 25143
rect 33600 25100 33652 25109
rect 34796 25168 34848 25220
rect 35992 25168 36044 25220
rect 36360 25279 36412 25288
rect 36360 25245 36369 25279
rect 36369 25245 36403 25279
rect 36403 25245 36412 25279
rect 36360 25236 36412 25245
rect 36820 25304 36872 25356
rect 37464 25304 37516 25356
rect 36912 25236 36964 25288
rect 38016 25279 38068 25288
rect 38016 25245 38025 25279
rect 38025 25245 38059 25279
rect 38059 25245 38068 25279
rect 38016 25236 38068 25245
rect 35348 25143 35400 25152
rect 35348 25109 35357 25143
rect 35357 25109 35391 25143
rect 35391 25109 35400 25143
rect 35348 25100 35400 25109
rect 36176 25100 36228 25152
rect 36452 25100 36504 25152
rect 37740 25100 37792 25152
rect 38476 25100 38528 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 1860 24896 1912 24948
rect 3792 24896 3844 24948
rect 5264 24896 5316 24948
rect 8484 24896 8536 24948
rect 3516 24828 3568 24880
rect 4712 24828 4764 24880
rect 7564 24871 7616 24880
rect 7564 24837 7573 24871
rect 7573 24837 7607 24871
rect 7607 24837 7616 24871
rect 7564 24828 7616 24837
rect 9404 24871 9456 24880
rect 9404 24837 9413 24871
rect 9413 24837 9447 24871
rect 9447 24837 9456 24871
rect 9404 24828 9456 24837
rect 10968 24828 11020 24880
rect 5264 24760 5316 24812
rect 5356 24760 5408 24812
rect 5540 24760 5592 24812
rect 5724 24803 5776 24812
rect 5724 24769 5733 24803
rect 5733 24769 5767 24803
rect 5767 24769 5776 24803
rect 5724 24760 5776 24769
rect 6092 24760 6144 24812
rect 9312 24803 9364 24812
rect 3884 24692 3936 24744
rect 9312 24769 9316 24803
rect 9316 24769 9350 24803
rect 9350 24769 9364 24803
rect 9312 24760 9364 24769
rect 9496 24803 9548 24812
rect 9496 24769 9505 24803
rect 9505 24769 9539 24803
rect 9539 24769 9548 24803
rect 9496 24760 9548 24769
rect 9680 24803 9732 24812
rect 9680 24769 9688 24803
rect 9688 24769 9722 24803
rect 9722 24769 9732 24803
rect 9680 24760 9732 24769
rect 9772 24803 9824 24812
rect 9772 24769 9781 24803
rect 9781 24769 9815 24803
rect 9815 24769 9824 24803
rect 9772 24760 9824 24769
rect 10416 24760 10468 24812
rect 10600 24760 10652 24812
rect 10876 24803 10928 24812
rect 10876 24769 10885 24803
rect 10885 24769 10919 24803
rect 10919 24769 10928 24803
rect 10876 24760 10928 24769
rect 11980 24896 12032 24948
rect 3700 24624 3752 24676
rect 9496 24624 9548 24676
rect 2964 24556 3016 24608
rect 5908 24556 5960 24608
rect 6736 24556 6788 24608
rect 7288 24556 7340 24608
rect 7380 24556 7432 24608
rect 8116 24556 8168 24608
rect 9128 24599 9180 24608
rect 9128 24565 9137 24599
rect 9137 24565 9171 24599
rect 9171 24565 9180 24599
rect 9128 24556 9180 24565
rect 10784 24624 10836 24676
rect 11796 24803 11848 24812
rect 11796 24769 11805 24803
rect 11805 24769 11839 24803
rect 11839 24769 11848 24803
rect 11796 24760 11848 24769
rect 11980 24803 12032 24812
rect 11980 24769 11994 24803
rect 11994 24769 12028 24803
rect 12028 24769 12032 24803
rect 12256 24896 12308 24948
rect 15752 24896 15804 24948
rect 11980 24760 12032 24769
rect 14096 24760 14148 24812
rect 14464 24803 14516 24812
rect 14464 24769 14473 24803
rect 14473 24769 14507 24803
rect 14507 24769 14516 24803
rect 14464 24760 14516 24769
rect 14648 24760 14700 24812
rect 14740 24803 14792 24812
rect 14740 24769 14749 24803
rect 14749 24769 14783 24803
rect 14783 24769 14792 24803
rect 14740 24760 14792 24769
rect 15476 24803 15528 24812
rect 15476 24769 15485 24803
rect 15485 24769 15519 24803
rect 15519 24769 15528 24803
rect 15476 24760 15528 24769
rect 16304 24760 16356 24812
rect 17132 24896 17184 24948
rect 18604 24896 18656 24948
rect 20260 24896 20312 24948
rect 21272 24896 21324 24948
rect 22192 24896 22244 24948
rect 22560 24896 22612 24948
rect 23940 24896 23992 24948
rect 17684 24871 17736 24880
rect 17684 24837 17693 24871
rect 17693 24837 17727 24871
rect 17727 24837 17736 24871
rect 17684 24828 17736 24837
rect 15200 24692 15252 24744
rect 15660 24735 15712 24744
rect 15660 24701 15669 24735
rect 15669 24701 15703 24735
rect 15703 24701 15712 24735
rect 15660 24692 15712 24701
rect 17132 24803 17184 24812
rect 17132 24769 17141 24803
rect 17141 24769 17175 24803
rect 17175 24769 17184 24803
rect 17132 24760 17184 24769
rect 17316 24803 17368 24812
rect 17316 24769 17325 24803
rect 17325 24769 17359 24803
rect 17359 24769 17368 24803
rect 17316 24760 17368 24769
rect 17408 24803 17460 24812
rect 17408 24769 17417 24803
rect 17417 24769 17451 24803
rect 17451 24769 17460 24803
rect 17408 24760 17460 24769
rect 15936 24624 15988 24676
rect 18512 24760 18564 24812
rect 19064 24803 19116 24812
rect 19064 24769 19073 24803
rect 19073 24769 19107 24803
rect 19107 24769 19116 24803
rect 19064 24760 19116 24769
rect 18420 24692 18472 24744
rect 18880 24692 18932 24744
rect 12440 24556 12492 24608
rect 12532 24599 12584 24608
rect 12532 24565 12541 24599
rect 12541 24565 12575 24599
rect 12575 24565 12584 24599
rect 12532 24556 12584 24565
rect 12624 24556 12676 24608
rect 14556 24556 14608 24608
rect 16120 24556 16172 24608
rect 19892 24828 19944 24880
rect 20628 24828 20680 24880
rect 20076 24803 20128 24812
rect 20076 24769 20085 24803
rect 20085 24769 20119 24803
rect 20119 24769 20128 24803
rect 20076 24760 20128 24769
rect 19340 24692 19392 24744
rect 20720 24803 20772 24812
rect 20720 24769 20729 24803
rect 20729 24769 20763 24803
rect 20763 24769 20772 24803
rect 20720 24760 20772 24769
rect 21824 24828 21876 24880
rect 24400 24871 24452 24880
rect 24400 24837 24409 24871
rect 24409 24837 24443 24871
rect 24443 24837 24452 24871
rect 24400 24828 24452 24837
rect 21088 24624 21140 24676
rect 21364 24735 21416 24744
rect 21364 24701 21373 24735
rect 21373 24701 21407 24735
rect 21407 24701 21416 24735
rect 21364 24692 21416 24701
rect 21456 24692 21508 24744
rect 21916 24803 21968 24812
rect 21916 24769 21958 24803
rect 21958 24769 21968 24803
rect 21916 24760 21968 24769
rect 22284 24760 22336 24812
rect 23664 24692 23716 24744
rect 22100 24624 22152 24676
rect 21456 24556 21508 24608
rect 21824 24599 21876 24608
rect 21824 24565 21833 24599
rect 21833 24565 21867 24599
rect 21867 24565 21876 24599
rect 21824 24556 21876 24565
rect 22376 24599 22428 24608
rect 22376 24565 22385 24599
rect 22385 24565 22419 24599
rect 22419 24565 22428 24599
rect 22376 24556 22428 24565
rect 24492 24803 24544 24812
rect 24492 24769 24501 24803
rect 24501 24769 24535 24803
rect 24535 24769 24544 24803
rect 24492 24760 24544 24769
rect 25688 24896 25740 24948
rect 25964 24939 26016 24948
rect 25964 24905 25989 24939
rect 25989 24905 26016 24939
rect 25964 24896 26016 24905
rect 24768 24803 24820 24812
rect 24768 24769 24777 24803
rect 24777 24769 24811 24803
rect 24811 24769 24820 24803
rect 24768 24760 24820 24769
rect 24952 24760 25004 24812
rect 25780 24871 25832 24880
rect 25780 24837 25789 24871
rect 25789 24837 25823 24871
rect 25823 24837 25832 24871
rect 25780 24828 25832 24837
rect 26976 24896 27028 24948
rect 25412 24692 25464 24744
rect 26516 24760 26568 24812
rect 24676 24624 24728 24676
rect 26884 24692 26936 24744
rect 27068 24735 27120 24744
rect 27068 24701 27077 24735
rect 27077 24701 27111 24735
rect 27111 24701 27120 24735
rect 27068 24692 27120 24701
rect 27252 24803 27304 24812
rect 27252 24769 27261 24803
rect 27261 24769 27295 24803
rect 27295 24769 27304 24803
rect 27252 24760 27304 24769
rect 27436 24760 27488 24812
rect 26332 24624 26384 24676
rect 25688 24556 25740 24608
rect 25780 24556 25832 24608
rect 26424 24599 26476 24608
rect 26424 24565 26433 24599
rect 26433 24565 26467 24599
rect 26467 24565 26476 24599
rect 26424 24556 26476 24565
rect 27160 24624 27212 24676
rect 28540 24803 28592 24812
rect 28540 24769 28549 24803
rect 28549 24769 28583 24803
rect 28583 24769 28592 24803
rect 28540 24760 28592 24769
rect 30656 24760 30708 24812
rect 30840 24760 30892 24812
rect 33324 24896 33376 24948
rect 36728 24896 36780 24948
rect 40040 24939 40092 24948
rect 40040 24905 40049 24939
rect 40049 24905 40083 24939
rect 40083 24905 40092 24939
rect 40040 24896 40092 24905
rect 28908 24692 28960 24744
rect 30288 24735 30340 24744
rect 30288 24701 30297 24735
rect 30297 24701 30331 24735
rect 30331 24701 30340 24735
rect 30288 24692 30340 24701
rect 34152 24828 34204 24880
rect 38844 24871 38896 24880
rect 38844 24837 38853 24871
rect 38853 24837 38887 24871
rect 38887 24837 38896 24871
rect 38844 24828 38896 24837
rect 31760 24760 31812 24812
rect 31852 24692 31904 24744
rect 32956 24692 33008 24744
rect 35256 24803 35308 24812
rect 35256 24769 35265 24803
rect 35265 24769 35299 24803
rect 35299 24769 35308 24803
rect 35256 24760 35308 24769
rect 35348 24760 35400 24812
rect 37464 24803 37516 24812
rect 37464 24769 37473 24803
rect 37473 24769 37507 24803
rect 37507 24769 37516 24803
rect 37464 24760 37516 24769
rect 37740 24803 37792 24812
rect 37740 24769 37749 24803
rect 37749 24769 37783 24803
rect 37783 24769 37792 24803
rect 37740 24760 37792 24769
rect 38016 24760 38068 24812
rect 38292 24760 38344 24812
rect 36636 24692 36688 24744
rect 36820 24692 36872 24744
rect 37924 24692 37976 24744
rect 38200 24692 38252 24744
rect 38936 24760 38988 24812
rect 40224 24803 40276 24812
rect 40224 24769 40233 24803
rect 40233 24769 40267 24803
rect 40267 24769 40276 24803
rect 40224 24760 40276 24769
rect 31944 24624 31996 24676
rect 35348 24624 35400 24676
rect 37004 24624 37056 24676
rect 27344 24556 27396 24608
rect 27528 24599 27580 24608
rect 27528 24565 27537 24599
rect 27537 24565 27571 24599
rect 27571 24565 27580 24599
rect 27528 24556 27580 24565
rect 27988 24599 28040 24608
rect 27988 24565 27997 24599
rect 27997 24565 28031 24599
rect 28031 24565 28040 24599
rect 27988 24556 28040 24565
rect 28172 24599 28224 24608
rect 28172 24565 28181 24599
rect 28181 24565 28215 24599
rect 28215 24565 28224 24599
rect 28172 24556 28224 24565
rect 28448 24556 28500 24608
rect 33140 24556 33192 24608
rect 37280 24599 37332 24608
rect 37280 24565 37289 24599
rect 37289 24565 37323 24599
rect 37323 24565 37332 24599
rect 37280 24556 37332 24565
rect 39120 24692 39172 24744
rect 39396 24556 39448 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 3884 24352 3936 24404
rect 2872 24216 2924 24268
rect 3700 24216 3752 24268
rect 5724 24216 5776 24268
rect 8024 24352 8076 24404
rect 8116 24352 8168 24404
rect 9680 24352 9732 24404
rect 13636 24352 13688 24404
rect 14464 24352 14516 24404
rect 6368 24284 6420 24336
rect 3148 24148 3200 24200
rect 6276 24148 6328 24200
rect 1676 24123 1728 24132
rect 1676 24089 1685 24123
rect 1685 24089 1719 24123
rect 1719 24089 1728 24123
rect 1676 24080 1728 24089
rect 4068 24123 4120 24132
rect 4068 24089 4077 24123
rect 4077 24089 4111 24123
rect 4111 24089 4120 24123
rect 4068 24080 4120 24089
rect 4620 24080 4672 24132
rect 6000 24080 6052 24132
rect 6552 24191 6604 24200
rect 6552 24157 6561 24191
rect 6561 24157 6595 24191
rect 6595 24157 6604 24191
rect 6552 24148 6604 24157
rect 6828 24284 6880 24336
rect 7656 24284 7708 24336
rect 7840 24284 7892 24336
rect 8300 24284 8352 24336
rect 7840 24148 7892 24200
rect 9036 24284 9088 24336
rect 9312 24284 9364 24336
rect 5632 24055 5684 24064
rect 5632 24021 5641 24055
rect 5641 24021 5675 24055
rect 5675 24021 5684 24055
rect 5632 24012 5684 24021
rect 7380 24080 7432 24132
rect 8392 24123 8444 24132
rect 8392 24089 8401 24123
rect 8401 24089 8435 24123
rect 8435 24089 8444 24123
rect 8392 24080 8444 24089
rect 8576 24012 8628 24064
rect 8668 24055 8720 24064
rect 8668 24021 8677 24055
rect 8677 24021 8711 24055
rect 8711 24021 8720 24055
rect 8668 24012 8720 24021
rect 9220 24191 9272 24200
rect 9220 24157 9229 24191
rect 9229 24157 9263 24191
rect 9263 24157 9272 24191
rect 9220 24148 9272 24157
rect 10876 24216 10928 24268
rect 11336 24259 11388 24268
rect 11336 24225 11345 24259
rect 11345 24225 11379 24259
rect 11379 24225 11388 24259
rect 14924 24284 14976 24336
rect 15660 24352 15712 24404
rect 17316 24352 17368 24404
rect 11336 24216 11388 24225
rect 10416 24148 10468 24200
rect 10600 24148 10652 24200
rect 11244 24148 11296 24200
rect 12624 24148 12676 24200
rect 13912 24148 13964 24200
rect 14740 24216 14792 24268
rect 15476 24284 15528 24336
rect 15752 24327 15804 24336
rect 15752 24293 15761 24327
rect 15761 24293 15795 24327
rect 15795 24293 15804 24327
rect 15752 24284 15804 24293
rect 18972 24284 19024 24336
rect 19892 24284 19944 24336
rect 20904 24284 20956 24336
rect 16304 24216 16356 24268
rect 18604 24216 18656 24268
rect 19524 24216 19576 24268
rect 20076 24216 20128 24268
rect 9312 24123 9364 24132
rect 9312 24089 9321 24123
rect 9321 24089 9355 24123
rect 9355 24089 9364 24123
rect 9312 24080 9364 24089
rect 12256 24080 12308 24132
rect 10876 24012 10928 24064
rect 14556 24191 14608 24200
rect 14556 24157 14565 24191
rect 14565 24157 14599 24191
rect 14599 24157 14608 24191
rect 14556 24148 14608 24157
rect 15292 24148 15344 24200
rect 15476 24148 15528 24200
rect 14924 24080 14976 24132
rect 16396 24191 16448 24200
rect 16396 24157 16405 24191
rect 16405 24157 16439 24191
rect 16439 24157 16448 24191
rect 16396 24148 16448 24157
rect 17960 24191 18012 24200
rect 17960 24157 17969 24191
rect 17969 24157 18003 24191
rect 18003 24157 18012 24191
rect 17960 24148 18012 24157
rect 17040 24080 17092 24132
rect 19156 24148 19208 24200
rect 18420 24080 18472 24132
rect 18512 24080 18564 24132
rect 20628 24148 20680 24200
rect 23020 24191 23072 24200
rect 23020 24157 23029 24191
rect 23029 24157 23063 24191
rect 23063 24157 23072 24191
rect 23020 24148 23072 24157
rect 23848 24395 23900 24404
rect 23848 24361 23857 24395
rect 23857 24361 23891 24395
rect 23891 24361 23900 24395
rect 23848 24352 23900 24361
rect 24124 24395 24176 24404
rect 24124 24361 24133 24395
rect 24133 24361 24167 24395
rect 24167 24361 24176 24395
rect 24124 24352 24176 24361
rect 25596 24352 25648 24404
rect 25872 24352 25924 24404
rect 26700 24352 26752 24404
rect 26976 24352 27028 24404
rect 27344 24352 27396 24404
rect 25136 24284 25188 24336
rect 27528 24284 27580 24336
rect 28356 24352 28408 24404
rect 30932 24352 30984 24404
rect 32496 24352 32548 24404
rect 33508 24352 33560 24404
rect 36084 24352 36136 24404
rect 37924 24395 37976 24404
rect 37924 24361 37933 24395
rect 37933 24361 37967 24395
rect 37967 24361 37976 24395
rect 37924 24352 37976 24361
rect 29644 24284 29696 24336
rect 39488 24352 39540 24404
rect 39672 24352 39724 24404
rect 23480 24191 23532 24200
rect 23480 24157 23494 24191
rect 23494 24157 23528 24191
rect 23528 24157 23532 24191
rect 23480 24148 23532 24157
rect 23664 24148 23716 24200
rect 24400 24216 24452 24268
rect 24768 24216 24820 24268
rect 27252 24216 27304 24268
rect 23848 24148 23900 24200
rect 24676 24148 24728 24200
rect 25136 24148 25188 24200
rect 25872 24191 25924 24200
rect 15936 24012 15988 24064
rect 19984 24055 20036 24064
rect 19984 24021 19993 24055
rect 19993 24021 20027 24055
rect 20027 24021 20036 24055
rect 19984 24012 20036 24021
rect 20076 24012 20128 24064
rect 20904 24080 20956 24132
rect 24216 24080 24268 24132
rect 25872 24157 25881 24191
rect 25881 24157 25915 24191
rect 25915 24157 25924 24191
rect 25872 24148 25924 24157
rect 26700 24148 26752 24200
rect 27988 24216 28040 24268
rect 27528 24191 27580 24200
rect 27528 24157 27537 24191
rect 27537 24157 27571 24191
rect 27571 24157 27580 24191
rect 27528 24148 27580 24157
rect 27712 24191 27764 24200
rect 27712 24157 27721 24191
rect 27721 24157 27755 24191
rect 27755 24157 27764 24191
rect 27712 24148 27764 24157
rect 25780 24080 25832 24132
rect 23480 24012 23532 24064
rect 23664 24012 23716 24064
rect 25872 24012 25924 24064
rect 26424 24123 26476 24132
rect 26424 24089 26433 24123
rect 26433 24089 26467 24123
rect 26467 24089 26476 24123
rect 26424 24080 26476 24089
rect 27436 24012 27488 24064
rect 27528 24012 27580 24064
rect 28080 24191 28132 24200
rect 28080 24157 28089 24191
rect 28089 24157 28123 24191
rect 28123 24157 28132 24191
rect 28080 24148 28132 24157
rect 28724 24216 28776 24268
rect 28448 24191 28500 24200
rect 28448 24157 28457 24191
rect 28457 24157 28491 24191
rect 28491 24157 28500 24191
rect 28448 24148 28500 24157
rect 28540 24191 28592 24200
rect 28540 24157 28554 24191
rect 28554 24157 28588 24191
rect 28588 24157 28592 24191
rect 28540 24148 28592 24157
rect 29000 24191 29052 24200
rect 29000 24157 29009 24191
rect 29009 24157 29043 24191
rect 29043 24157 29052 24191
rect 29000 24148 29052 24157
rect 37832 24216 37884 24268
rect 36544 24148 36596 24200
rect 38568 24284 38620 24336
rect 39396 24148 39448 24200
rect 39672 24191 39724 24200
rect 39672 24157 39681 24191
rect 39681 24157 39715 24191
rect 39715 24157 39724 24191
rect 39672 24148 39724 24157
rect 40132 24148 40184 24200
rect 28632 24080 28684 24132
rect 38200 24123 38252 24132
rect 38200 24089 38209 24123
rect 38209 24089 38243 24123
rect 38243 24089 38252 24123
rect 38200 24080 38252 24089
rect 31116 24012 31168 24064
rect 35348 24012 35400 24064
rect 37096 24012 37148 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 1676 23808 1728 23860
rect 2964 23808 3016 23860
rect 5632 23808 5684 23860
rect 3700 23783 3752 23792
rect 3700 23749 3709 23783
rect 3709 23749 3743 23783
rect 3743 23749 3752 23783
rect 3700 23740 3752 23749
rect 4620 23740 4672 23792
rect 5448 23740 5500 23792
rect 6000 23808 6052 23860
rect 6736 23808 6788 23860
rect 7840 23851 7892 23860
rect 7840 23817 7849 23851
rect 7849 23817 7883 23851
rect 7883 23817 7892 23851
rect 7840 23808 7892 23817
rect 3056 23672 3108 23724
rect 3884 23672 3936 23724
rect 6828 23740 6880 23792
rect 4068 23536 4120 23588
rect 5080 23647 5132 23656
rect 5080 23613 5089 23647
rect 5089 23613 5123 23647
rect 5123 23613 5132 23647
rect 5080 23604 5132 23613
rect 5264 23647 5316 23656
rect 5264 23613 5273 23647
rect 5273 23613 5307 23647
rect 5307 23613 5316 23647
rect 5264 23604 5316 23613
rect 5540 23604 5592 23656
rect 6184 23715 6236 23724
rect 6184 23681 6193 23715
rect 6193 23681 6227 23715
rect 6227 23681 6236 23715
rect 6184 23672 6236 23681
rect 6276 23672 6328 23724
rect 6552 23715 6604 23724
rect 6552 23681 6561 23715
rect 6561 23681 6595 23715
rect 6595 23681 6604 23715
rect 6552 23672 6604 23681
rect 7380 23672 7432 23724
rect 7932 23672 7984 23724
rect 8208 23715 8260 23724
rect 8208 23681 8217 23715
rect 8217 23681 8251 23715
rect 8251 23681 8260 23715
rect 10416 23808 10468 23860
rect 10508 23808 10560 23860
rect 8208 23672 8260 23681
rect 11060 23740 11112 23792
rect 18420 23808 18472 23860
rect 19156 23851 19208 23860
rect 19156 23817 19165 23851
rect 19165 23817 19199 23851
rect 19199 23817 19208 23851
rect 19156 23808 19208 23817
rect 8116 23604 8168 23656
rect 8668 23672 8720 23724
rect 8852 23715 8904 23724
rect 8852 23681 8861 23715
rect 8861 23681 8895 23715
rect 8895 23681 8904 23715
rect 8852 23672 8904 23681
rect 9404 23672 9456 23724
rect 9772 23672 9824 23724
rect 10508 23672 10560 23724
rect 10692 23672 10744 23724
rect 5632 23511 5684 23520
rect 5632 23477 5641 23511
rect 5641 23477 5675 23511
rect 5675 23477 5684 23511
rect 5632 23468 5684 23477
rect 6184 23468 6236 23520
rect 6368 23511 6420 23520
rect 6368 23477 6377 23511
rect 6377 23477 6411 23511
rect 6411 23477 6420 23511
rect 6368 23468 6420 23477
rect 8300 23536 8352 23588
rect 8576 23511 8628 23520
rect 8576 23477 8585 23511
rect 8585 23477 8619 23511
rect 8619 23477 8628 23511
rect 8576 23468 8628 23477
rect 11520 23672 11572 23724
rect 11888 23672 11940 23724
rect 13544 23672 13596 23724
rect 13728 23672 13780 23724
rect 14648 23672 14700 23724
rect 15200 23715 15252 23724
rect 15200 23681 15209 23715
rect 15209 23681 15243 23715
rect 15243 23681 15252 23715
rect 15200 23672 15252 23681
rect 15476 23715 15528 23724
rect 15476 23681 15485 23715
rect 15485 23681 15519 23715
rect 15519 23681 15528 23715
rect 15476 23672 15528 23681
rect 15660 23672 15712 23724
rect 16120 23672 16172 23724
rect 11336 23604 11388 23656
rect 11704 23604 11756 23656
rect 10692 23579 10744 23588
rect 10692 23545 10701 23579
rect 10701 23545 10735 23579
rect 10735 23545 10744 23579
rect 10692 23536 10744 23545
rect 11152 23468 11204 23520
rect 11244 23468 11296 23520
rect 12440 23647 12492 23656
rect 12440 23613 12449 23647
rect 12449 23613 12483 23647
rect 12483 23613 12492 23647
rect 12440 23604 12492 23613
rect 13912 23604 13964 23656
rect 18052 23740 18104 23792
rect 16764 23672 16816 23724
rect 17960 23672 18012 23724
rect 18972 23740 19024 23792
rect 19892 23808 19944 23860
rect 20444 23851 20496 23860
rect 20444 23817 20453 23851
rect 20453 23817 20487 23851
rect 20487 23817 20496 23851
rect 20444 23808 20496 23817
rect 23756 23851 23808 23860
rect 23756 23817 23765 23851
rect 23765 23817 23799 23851
rect 23799 23817 23808 23851
rect 23756 23808 23808 23817
rect 13544 23536 13596 23588
rect 17040 23647 17092 23656
rect 17040 23613 17049 23647
rect 17049 23613 17083 23647
rect 17083 23613 17092 23647
rect 17040 23604 17092 23613
rect 17408 23604 17460 23656
rect 18052 23604 18104 23656
rect 18420 23604 18472 23656
rect 19524 23715 19576 23724
rect 19524 23681 19533 23715
rect 19533 23681 19567 23715
rect 19567 23681 19576 23715
rect 19524 23672 19576 23681
rect 19892 23715 19944 23724
rect 19892 23681 19901 23715
rect 19901 23681 19935 23715
rect 19935 23681 19944 23715
rect 19892 23672 19944 23681
rect 20352 23740 20404 23792
rect 20628 23783 20680 23792
rect 20628 23749 20655 23783
rect 20655 23749 20680 23783
rect 20628 23740 20680 23749
rect 21272 23740 21324 23792
rect 16580 23536 16632 23588
rect 13912 23511 13964 23520
rect 13912 23477 13921 23511
rect 13921 23477 13955 23511
rect 13955 23477 13964 23511
rect 13912 23468 13964 23477
rect 14004 23511 14056 23520
rect 14004 23477 14013 23511
rect 14013 23477 14047 23511
rect 14047 23477 14056 23511
rect 14004 23468 14056 23477
rect 15476 23468 15528 23520
rect 15936 23511 15988 23520
rect 15936 23477 15945 23511
rect 15945 23477 15979 23511
rect 15979 23477 15988 23511
rect 15936 23468 15988 23477
rect 19064 23647 19116 23656
rect 19064 23613 19073 23647
rect 19073 23613 19107 23647
rect 19107 23613 19116 23647
rect 19064 23604 19116 23613
rect 19156 23604 19208 23656
rect 19340 23604 19392 23656
rect 22560 23715 22612 23724
rect 22560 23681 22569 23715
rect 22569 23681 22603 23715
rect 22603 23681 22612 23715
rect 22560 23672 22612 23681
rect 22744 23715 22796 23724
rect 22744 23681 22753 23715
rect 22753 23681 22787 23715
rect 22787 23681 22796 23715
rect 22744 23672 22796 23681
rect 23112 23672 23164 23724
rect 20812 23604 20864 23656
rect 22100 23536 22152 23588
rect 23756 23672 23808 23724
rect 25596 23740 25648 23792
rect 26424 23740 26476 23792
rect 27712 23808 27764 23860
rect 27252 23740 27304 23792
rect 28724 23808 28776 23860
rect 29000 23808 29052 23860
rect 31116 23851 31168 23860
rect 31116 23817 31125 23851
rect 31125 23817 31159 23851
rect 31159 23817 31168 23851
rect 31116 23808 31168 23817
rect 33508 23851 33560 23860
rect 33508 23817 33517 23851
rect 33517 23817 33551 23851
rect 33551 23817 33560 23851
rect 33508 23808 33560 23817
rect 33600 23808 33652 23860
rect 24032 23672 24084 23724
rect 23480 23604 23532 23656
rect 24216 23647 24268 23656
rect 24216 23613 24225 23647
rect 24225 23613 24259 23647
rect 24259 23613 24268 23647
rect 24216 23604 24268 23613
rect 26700 23604 26752 23656
rect 27988 23672 28040 23724
rect 28356 23715 28408 23724
rect 28356 23681 28365 23715
rect 28365 23681 28399 23715
rect 28399 23681 28408 23715
rect 28356 23672 28408 23681
rect 28540 23715 28592 23724
rect 28540 23681 28549 23715
rect 28549 23681 28583 23715
rect 28583 23681 28592 23715
rect 28540 23672 28592 23681
rect 28724 23672 28776 23724
rect 28908 23715 28960 23724
rect 28908 23681 28917 23715
rect 28917 23681 28951 23715
rect 28951 23681 28960 23715
rect 28908 23672 28960 23681
rect 29184 23740 29236 23792
rect 29644 23783 29696 23792
rect 29644 23749 29653 23783
rect 29653 23749 29687 23783
rect 29687 23749 29696 23783
rect 29644 23740 29696 23749
rect 34520 23808 34572 23860
rect 30380 23672 30432 23724
rect 30932 23672 30984 23724
rect 31484 23672 31536 23724
rect 32956 23672 33008 23724
rect 33140 23672 33192 23724
rect 32312 23604 32364 23656
rect 33692 23604 33744 23656
rect 34336 23715 34388 23724
rect 34336 23681 34345 23715
rect 34345 23681 34379 23715
rect 34379 23681 34388 23715
rect 34336 23672 34388 23681
rect 36360 23783 36412 23792
rect 36360 23749 36369 23783
rect 36369 23749 36403 23783
rect 36403 23749 36412 23783
rect 36360 23740 36412 23749
rect 19340 23468 19392 23520
rect 20076 23468 20128 23520
rect 21272 23468 21324 23520
rect 23848 23536 23900 23588
rect 28172 23536 28224 23588
rect 28908 23536 28960 23588
rect 29276 23579 29328 23588
rect 29276 23545 29285 23579
rect 29285 23545 29319 23579
rect 29319 23545 29328 23579
rect 29276 23536 29328 23545
rect 31024 23536 31076 23588
rect 31484 23536 31536 23588
rect 34152 23536 34204 23588
rect 34888 23715 34940 23724
rect 34888 23681 34897 23715
rect 34897 23681 34931 23715
rect 34931 23681 34940 23715
rect 34888 23672 34940 23681
rect 37556 23672 37608 23724
rect 34796 23604 34848 23656
rect 38844 23808 38896 23860
rect 38384 23740 38436 23792
rect 39580 23672 39632 23724
rect 38200 23647 38252 23656
rect 38200 23613 38209 23647
rect 38209 23613 38243 23647
rect 38243 23613 38252 23647
rect 38200 23604 38252 23613
rect 39120 23604 39172 23656
rect 39488 23604 39540 23656
rect 28816 23468 28868 23520
rect 31576 23468 31628 23520
rect 32312 23468 32364 23520
rect 33048 23511 33100 23520
rect 33048 23477 33057 23511
rect 33057 23477 33091 23511
rect 33091 23477 33100 23511
rect 33048 23468 33100 23477
rect 34796 23468 34848 23520
rect 37924 23468 37976 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 4712 23264 4764 23316
rect 9220 23264 9272 23316
rect 9496 23264 9548 23316
rect 10324 23307 10376 23316
rect 10324 23273 10333 23307
rect 10333 23273 10367 23307
rect 10367 23273 10376 23307
rect 10324 23264 10376 23273
rect 11520 23307 11572 23316
rect 11520 23273 11529 23307
rect 11529 23273 11563 23307
rect 11563 23273 11572 23307
rect 11520 23264 11572 23273
rect 5632 23239 5684 23248
rect 5632 23205 5641 23239
rect 5641 23205 5675 23239
rect 5675 23205 5684 23239
rect 5632 23196 5684 23205
rect 3240 23128 3292 23180
rect 2872 23060 2924 23112
rect 3976 23060 4028 23112
rect 5264 23060 5316 23112
rect 6276 23128 6328 23180
rect 8392 23196 8444 23248
rect 8944 23196 8996 23248
rect 11980 23196 12032 23248
rect 12164 23307 12216 23316
rect 12164 23273 12173 23307
rect 12173 23273 12207 23307
rect 12207 23273 12216 23307
rect 12164 23264 12216 23273
rect 12440 23264 12492 23316
rect 16580 23307 16632 23316
rect 16580 23273 16589 23307
rect 16589 23273 16623 23307
rect 16623 23273 16632 23307
rect 16580 23264 16632 23273
rect 16672 23264 16724 23316
rect 18052 23307 18104 23316
rect 18052 23273 18061 23307
rect 18061 23273 18095 23307
rect 18095 23273 18104 23307
rect 18052 23264 18104 23273
rect 18696 23264 18748 23316
rect 19524 23264 19576 23316
rect 23296 23264 23348 23316
rect 24492 23264 24544 23316
rect 29276 23264 29328 23316
rect 34152 23264 34204 23316
rect 37280 23264 37332 23316
rect 38384 23264 38436 23316
rect 9772 23128 9824 23180
rect 10876 23128 10928 23180
rect 11520 23128 11572 23180
rect 12072 23128 12124 23180
rect 2596 22924 2648 22976
rect 5632 22992 5684 23044
rect 6092 23103 6144 23112
rect 6092 23069 6101 23103
rect 6101 23069 6135 23103
rect 6135 23069 6144 23103
rect 6092 23060 6144 23069
rect 6368 23103 6420 23112
rect 6368 23069 6377 23103
rect 6377 23069 6411 23103
rect 6411 23069 6420 23103
rect 6368 23060 6420 23069
rect 6736 23103 6788 23112
rect 6736 23069 6745 23103
rect 6745 23069 6779 23103
rect 6779 23069 6788 23103
rect 6736 23060 6788 23069
rect 7840 23060 7892 23112
rect 8944 23103 8996 23112
rect 8944 23069 8953 23103
rect 8953 23069 8987 23103
rect 8987 23069 8996 23103
rect 8944 23060 8996 23069
rect 10508 23103 10560 23112
rect 10508 23069 10517 23103
rect 10517 23069 10551 23103
rect 10551 23069 10560 23103
rect 10508 23060 10560 23069
rect 6276 22992 6328 23044
rect 7748 22924 7800 22976
rect 9496 22924 9548 22976
rect 9772 23035 9824 23044
rect 9772 23001 9781 23035
rect 9781 23001 9815 23035
rect 9815 23001 9824 23035
rect 9772 22992 9824 23001
rect 10416 22992 10468 23044
rect 9956 22924 10008 22976
rect 11336 23060 11388 23112
rect 11704 23035 11756 23044
rect 11704 23001 11713 23035
rect 11713 23001 11747 23035
rect 11747 23001 11756 23035
rect 11704 22992 11756 23001
rect 10692 22924 10744 22976
rect 10968 22967 11020 22976
rect 10968 22933 10977 22967
rect 10977 22933 11011 22967
rect 11011 22933 11020 22967
rect 10968 22924 11020 22933
rect 11428 22924 11480 22976
rect 11520 22924 11572 22976
rect 14740 23239 14792 23248
rect 14740 23205 14749 23239
rect 14749 23205 14783 23239
rect 14783 23205 14792 23239
rect 14740 23196 14792 23205
rect 13176 23128 13228 23180
rect 13452 23128 13504 23180
rect 19064 23196 19116 23248
rect 19156 23196 19208 23248
rect 25872 23196 25924 23248
rect 27804 23196 27856 23248
rect 28908 23196 28960 23248
rect 30196 23196 30248 23248
rect 18696 23128 18748 23180
rect 24032 23128 24084 23180
rect 34520 23196 34572 23248
rect 32036 23128 32088 23180
rect 33048 23171 33100 23180
rect 33048 23137 33057 23171
rect 33057 23137 33091 23171
rect 33091 23137 33100 23171
rect 33048 23128 33100 23137
rect 33232 23128 33284 23180
rect 33416 23128 33468 23180
rect 33692 23128 33744 23180
rect 37556 23196 37608 23248
rect 38476 23196 38528 23248
rect 39580 23264 39632 23316
rect 14004 23060 14056 23112
rect 14372 23060 14424 23112
rect 12164 22992 12216 23044
rect 13544 22992 13596 23044
rect 13820 23035 13872 23044
rect 13820 23001 13829 23035
rect 13829 23001 13863 23035
rect 13863 23001 13872 23035
rect 13820 22992 13872 23001
rect 16948 23060 17000 23112
rect 18236 23060 18288 23112
rect 18420 23103 18472 23112
rect 18420 23069 18429 23103
rect 18429 23069 18463 23103
rect 18463 23069 18472 23103
rect 18420 23060 18472 23069
rect 18788 23103 18840 23112
rect 18788 23069 18797 23103
rect 18797 23069 18831 23103
rect 18831 23069 18840 23103
rect 18788 23060 18840 23069
rect 19340 23060 19392 23112
rect 14004 22924 14056 22976
rect 19524 22992 19576 23044
rect 20076 23060 20128 23112
rect 20904 23060 20956 23112
rect 21364 23060 21416 23112
rect 22284 23103 22336 23112
rect 22284 23069 22293 23103
rect 22293 23069 22327 23103
rect 22327 23069 22336 23103
rect 22284 23060 22336 23069
rect 22836 23060 22888 23112
rect 23112 23060 23164 23112
rect 29828 23060 29880 23112
rect 21456 22992 21508 23044
rect 29276 23035 29328 23044
rect 29276 23001 29285 23035
rect 29285 23001 29319 23035
rect 29319 23001 29328 23035
rect 29276 22992 29328 23001
rect 31208 23103 31260 23112
rect 31208 23069 31217 23103
rect 31217 23069 31251 23103
rect 31251 23069 31260 23103
rect 31208 23060 31260 23069
rect 31300 23060 31352 23112
rect 31760 23060 31812 23112
rect 14280 22967 14332 22976
rect 14280 22933 14289 22967
rect 14289 22933 14323 22967
rect 14323 22933 14332 22967
rect 14280 22924 14332 22933
rect 17684 22967 17736 22976
rect 17684 22933 17693 22967
rect 17693 22933 17727 22967
rect 17727 22933 17736 22967
rect 17684 22924 17736 22933
rect 17960 22924 18012 22976
rect 18052 22924 18104 22976
rect 18696 22967 18748 22976
rect 18696 22933 18705 22967
rect 18705 22933 18739 22967
rect 18739 22933 18748 22967
rect 18696 22924 18748 22933
rect 19248 22924 19300 22976
rect 19984 22924 20036 22976
rect 21364 22924 21416 22976
rect 27712 22924 27764 22976
rect 28356 22924 28408 22976
rect 31116 22992 31168 23044
rect 33968 23060 34020 23112
rect 31668 22924 31720 22976
rect 33232 22992 33284 23044
rect 33508 22992 33560 23044
rect 34244 22992 34296 23044
rect 35992 22992 36044 23044
rect 32864 22967 32916 22976
rect 32864 22933 32873 22967
rect 32873 22933 32907 22967
rect 32907 22933 32916 22967
rect 32864 22924 32916 22933
rect 33692 22924 33744 22976
rect 35900 22924 35952 22976
rect 36452 23103 36504 23112
rect 36452 23069 36461 23103
rect 36461 23069 36495 23103
rect 36495 23069 36504 23103
rect 36452 23060 36504 23069
rect 36544 23103 36596 23112
rect 39304 23128 39356 23180
rect 39488 23128 39540 23180
rect 36544 23069 36558 23103
rect 36558 23069 36592 23103
rect 36592 23069 36596 23103
rect 36544 23060 36596 23069
rect 38568 23103 38620 23112
rect 38568 23069 38577 23103
rect 38577 23069 38611 23103
rect 38611 23069 38620 23103
rect 38568 23060 38620 23069
rect 39764 23060 39816 23112
rect 37372 22992 37424 23044
rect 38660 22992 38712 23044
rect 38016 22924 38068 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 2596 22763 2648 22772
rect 2596 22729 2605 22763
rect 2605 22729 2639 22763
rect 2639 22729 2648 22763
rect 2596 22720 2648 22729
rect 3056 22720 3108 22772
rect 6736 22720 6788 22772
rect 8116 22720 8168 22772
rect 9312 22720 9364 22772
rect 12348 22720 12400 22772
rect 12624 22720 12676 22772
rect 13636 22720 13688 22772
rect 14280 22720 14332 22772
rect 18052 22720 18104 22772
rect 18236 22720 18288 22772
rect 18604 22720 18656 22772
rect 20352 22720 20404 22772
rect 20628 22720 20680 22772
rect 2872 22584 2924 22636
rect 3332 22559 3384 22568
rect 3332 22525 3341 22559
rect 3341 22525 3375 22559
rect 3375 22525 3384 22559
rect 3332 22516 3384 22525
rect 3792 22516 3844 22568
rect 4712 22652 4764 22704
rect 8024 22652 8076 22704
rect 5724 22584 5776 22636
rect 6184 22584 6236 22636
rect 2872 22448 2924 22500
rect 4712 22448 4764 22500
rect 5264 22448 5316 22500
rect 6736 22516 6788 22568
rect 8576 22584 8628 22636
rect 10508 22652 10560 22704
rect 10232 22584 10284 22636
rect 10876 22627 10928 22636
rect 10876 22593 10885 22627
rect 10885 22593 10919 22627
rect 10919 22593 10928 22627
rect 10876 22584 10928 22593
rect 11336 22652 11388 22704
rect 8576 22491 8628 22500
rect 8576 22457 8585 22491
rect 8585 22457 8619 22491
rect 8619 22457 8628 22491
rect 8576 22448 8628 22457
rect 9496 22559 9548 22568
rect 9496 22525 9505 22559
rect 9505 22525 9539 22559
rect 9539 22525 9548 22559
rect 9496 22516 9548 22525
rect 11612 22516 11664 22568
rect 11980 22627 12032 22636
rect 11980 22593 11989 22627
rect 11989 22593 12023 22627
rect 12023 22593 12032 22627
rect 11980 22584 12032 22593
rect 14188 22695 14240 22704
rect 14188 22661 14197 22695
rect 14197 22661 14231 22695
rect 14231 22661 14240 22695
rect 14188 22652 14240 22661
rect 14004 22627 14056 22636
rect 14004 22593 14013 22627
rect 14013 22593 14047 22627
rect 14047 22593 14056 22627
rect 14004 22584 14056 22593
rect 19340 22584 19392 22636
rect 19892 22584 19944 22636
rect 20352 22627 20404 22636
rect 20352 22593 20361 22627
rect 20361 22593 20395 22627
rect 20395 22593 20404 22627
rect 20352 22584 20404 22593
rect 21456 22695 21508 22704
rect 21456 22661 21465 22695
rect 21465 22661 21499 22695
rect 21499 22661 21508 22695
rect 21456 22652 21508 22661
rect 22192 22720 22244 22772
rect 22928 22720 22980 22772
rect 25412 22763 25464 22772
rect 25412 22729 25421 22763
rect 25421 22729 25455 22763
rect 25455 22729 25464 22763
rect 25412 22720 25464 22729
rect 25688 22763 25740 22772
rect 25688 22729 25697 22763
rect 25697 22729 25731 22763
rect 25731 22729 25740 22763
rect 25688 22720 25740 22729
rect 26424 22720 26476 22772
rect 27528 22763 27580 22772
rect 27528 22729 27537 22763
rect 27537 22729 27571 22763
rect 27571 22729 27580 22763
rect 27528 22720 27580 22729
rect 27620 22720 27672 22772
rect 12164 22516 12216 22568
rect 12992 22516 13044 22568
rect 2228 22423 2280 22432
rect 2228 22389 2237 22423
rect 2237 22389 2271 22423
rect 2271 22389 2280 22423
rect 2228 22380 2280 22389
rect 3884 22380 3936 22432
rect 5632 22380 5684 22432
rect 7840 22380 7892 22432
rect 8944 22423 8996 22432
rect 8944 22389 8953 22423
rect 8953 22389 8987 22423
rect 8987 22389 8996 22423
rect 8944 22380 8996 22389
rect 9036 22380 9088 22432
rect 9588 22380 9640 22432
rect 10048 22423 10100 22432
rect 10048 22389 10057 22423
rect 10057 22389 10091 22423
rect 10091 22389 10100 22423
rect 10048 22380 10100 22389
rect 10232 22448 10284 22500
rect 16948 22448 17000 22500
rect 19984 22448 20036 22500
rect 20168 22516 20220 22568
rect 20444 22448 20496 22500
rect 12164 22380 12216 22432
rect 14556 22380 14608 22432
rect 16488 22380 16540 22432
rect 20812 22584 20864 22636
rect 25320 22652 25372 22704
rect 23756 22584 23808 22636
rect 24032 22627 24084 22636
rect 24032 22593 24041 22627
rect 24041 22593 24075 22627
rect 24075 22593 24084 22627
rect 24032 22584 24084 22593
rect 24124 22627 24176 22636
rect 24124 22593 24133 22627
rect 24133 22593 24167 22627
rect 24167 22593 24176 22627
rect 24124 22584 24176 22593
rect 24308 22627 24360 22636
rect 24308 22593 24317 22627
rect 24317 22593 24351 22627
rect 24351 22593 24360 22627
rect 24308 22584 24360 22593
rect 24492 22584 24544 22636
rect 24952 22584 25004 22636
rect 26332 22584 26384 22636
rect 25872 22516 25924 22568
rect 25964 22516 26016 22568
rect 26516 22516 26568 22568
rect 23296 22448 23348 22500
rect 26792 22584 26844 22636
rect 28448 22627 28500 22636
rect 28448 22593 28457 22627
rect 28457 22593 28491 22627
rect 28491 22593 28500 22627
rect 28448 22584 28500 22593
rect 28632 22584 28684 22636
rect 28908 22627 28960 22636
rect 28908 22593 28912 22627
rect 28912 22593 28946 22627
rect 28946 22593 28960 22627
rect 28908 22584 28960 22593
rect 29000 22627 29052 22636
rect 29000 22593 29009 22627
rect 29009 22593 29043 22627
rect 29043 22593 29052 22627
rect 29000 22584 29052 22593
rect 28724 22559 28776 22568
rect 28724 22525 28733 22559
rect 28733 22525 28767 22559
rect 28767 22525 28776 22559
rect 28724 22516 28776 22525
rect 20904 22423 20956 22432
rect 20904 22389 20913 22423
rect 20913 22389 20947 22423
rect 20947 22389 20956 22423
rect 20904 22380 20956 22389
rect 21088 22423 21140 22432
rect 21088 22389 21097 22423
rect 21097 22389 21131 22423
rect 21131 22389 21140 22423
rect 21088 22380 21140 22389
rect 21272 22423 21324 22432
rect 21272 22389 21281 22423
rect 21281 22389 21315 22423
rect 21315 22389 21324 22423
rect 21272 22380 21324 22389
rect 24676 22380 24728 22432
rect 25688 22380 25740 22432
rect 27068 22448 27120 22500
rect 28172 22448 28224 22500
rect 29644 22763 29696 22772
rect 29644 22729 29653 22763
rect 29653 22729 29687 22763
rect 29687 22729 29696 22763
rect 29644 22720 29696 22729
rect 30196 22720 30248 22772
rect 31852 22720 31904 22772
rect 32036 22720 32088 22772
rect 29460 22584 29512 22636
rect 29920 22627 29972 22636
rect 29920 22593 29929 22627
rect 29929 22593 29963 22627
rect 29963 22593 29972 22627
rect 29920 22584 29972 22593
rect 30380 22627 30432 22636
rect 30380 22593 30389 22627
rect 30389 22593 30423 22627
rect 30423 22593 30432 22627
rect 30380 22584 30432 22593
rect 30564 22516 30616 22568
rect 31392 22627 31444 22636
rect 31392 22593 31401 22627
rect 31401 22593 31435 22627
rect 31435 22593 31444 22627
rect 31392 22584 31444 22593
rect 31668 22627 31720 22636
rect 31668 22593 31677 22627
rect 31677 22593 31711 22627
rect 31711 22593 31720 22627
rect 31668 22584 31720 22593
rect 31760 22627 31812 22636
rect 31760 22593 31769 22627
rect 31769 22593 31803 22627
rect 31803 22593 31812 22627
rect 31760 22584 31812 22593
rect 31852 22584 31904 22636
rect 31576 22516 31628 22568
rect 32404 22627 32456 22636
rect 32404 22593 32413 22627
rect 32413 22593 32447 22627
rect 32447 22593 32456 22627
rect 32404 22584 32456 22593
rect 32864 22627 32916 22636
rect 32864 22593 32873 22627
rect 32873 22593 32907 22627
rect 32907 22593 32916 22627
rect 32864 22584 32916 22593
rect 33048 22627 33100 22636
rect 33048 22593 33057 22627
rect 33057 22593 33091 22627
rect 33091 22593 33100 22627
rect 33048 22584 33100 22593
rect 32680 22516 32732 22568
rect 34428 22652 34480 22704
rect 36268 22720 36320 22772
rect 33416 22584 33468 22636
rect 33876 22584 33928 22636
rect 35440 22584 35492 22636
rect 36176 22627 36228 22636
rect 36176 22593 36185 22627
rect 36185 22593 36219 22627
rect 36219 22593 36228 22627
rect 36176 22584 36228 22593
rect 36544 22584 36596 22636
rect 38016 22627 38068 22636
rect 38016 22593 38025 22627
rect 38025 22593 38059 22627
rect 38059 22593 38068 22627
rect 38016 22584 38068 22593
rect 27344 22380 27396 22432
rect 27620 22380 27672 22432
rect 28080 22423 28132 22432
rect 28080 22389 28089 22423
rect 28089 22389 28123 22423
rect 28123 22389 28132 22423
rect 28080 22380 28132 22389
rect 28448 22380 28500 22432
rect 30288 22448 30340 22500
rect 30012 22380 30064 22432
rect 31300 22380 31352 22432
rect 32128 22448 32180 22500
rect 34796 22516 34848 22568
rect 37924 22516 37976 22568
rect 38384 22516 38436 22568
rect 32864 22448 32916 22500
rect 37464 22448 37516 22500
rect 33048 22380 33100 22432
rect 37924 22380 37976 22432
rect 39764 22380 39816 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 2228 22176 2280 22228
rect 3240 22219 3292 22228
rect 3240 22185 3249 22219
rect 3249 22185 3283 22219
rect 3283 22185 3292 22219
rect 3240 22176 3292 22185
rect 1492 22015 1544 22024
rect 1492 21981 1501 22015
rect 1501 21981 1535 22015
rect 1535 21981 1544 22015
rect 1492 21972 1544 21981
rect 3056 21972 3108 22024
rect 3792 21972 3844 22024
rect 4620 21972 4672 22024
rect 5632 21972 5684 22024
rect 5448 21904 5500 21956
rect 5724 21904 5776 21956
rect 6276 22015 6328 22024
rect 6276 21981 6285 22015
rect 6285 21981 6319 22015
rect 6319 21981 6328 22015
rect 6276 21972 6328 21981
rect 6460 22108 6512 22160
rect 8576 22176 8628 22228
rect 8944 22176 8996 22228
rect 8208 22108 8260 22160
rect 6460 22015 6512 22024
rect 6460 21981 6469 22015
rect 6469 21981 6503 22015
rect 6503 21981 6512 22015
rect 6460 21972 6512 21981
rect 7012 22015 7064 22024
rect 7012 21981 7021 22015
rect 7021 21981 7055 22015
rect 7055 21981 7064 22015
rect 7012 21972 7064 21981
rect 7104 21904 7156 21956
rect 7840 21972 7892 22024
rect 10416 22040 10468 22092
rect 11244 22108 11296 22160
rect 11520 22151 11572 22160
rect 11520 22117 11529 22151
rect 11529 22117 11563 22151
rect 11563 22117 11572 22151
rect 11520 22108 11572 22117
rect 12072 22176 12124 22228
rect 12624 22108 12676 22160
rect 12900 22083 12952 22092
rect 12900 22049 12909 22083
rect 12909 22049 12943 22083
rect 12943 22049 12952 22083
rect 12900 22040 12952 22049
rect 8116 22015 8168 22024
rect 8116 21981 8125 22015
rect 8125 21981 8159 22015
rect 8159 21981 8168 22015
rect 8116 21972 8168 21981
rect 8484 22015 8536 22024
rect 8484 21981 8493 22015
rect 8493 21981 8527 22015
rect 8527 21981 8536 22015
rect 8484 21972 8536 21981
rect 8300 21947 8352 21956
rect 8300 21913 8309 21947
rect 8309 21913 8343 21947
rect 8343 21913 8352 21947
rect 8300 21904 8352 21913
rect 8576 21904 8628 21956
rect 5356 21879 5408 21888
rect 5356 21845 5365 21879
rect 5365 21845 5399 21879
rect 5399 21845 5408 21879
rect 5356 21836 5408 21845
rect 6644 21879 6696 21888
rect 6644 21845 6653 21879
rect 6653 21845 6687 21879
rect 6687 21845 6696 21879
rect 6644 21836 6696 21845
rect 7748 21836 7800 21888
rect 8208 21836 8260 21888
rect 10416 21947 10468 21956
rect 10416 21913 10425 21947
rect 10425 21913 10459 21947
rect 10459 21913 10468 21947
rect 10416 21904 10468 21913
rect 10508 21904 10560 21956
rect 10876 22015 10928 22024
rect 10876 21981 10885 22015
rect 10885 21981 10919 22015
rect 10919 21981 10928 22015
rect 10876 21972 10928 21981
rect 11060 22015 11112 22024
rect 11060 21981 11069 22015
rect 11069 21981 11103 22015
rect 11103 21981 11112 22015
rect 11060 21972 11112 21981
rect 11152 22015 11204 22024
rect 11152 21981 11161 22015
rect 11161 21981 11195 22015
rect 11195 21981 11204 22015
rect 11152 21972 11204 21981
rect 11612 22015 11664 22024
rect 11612 21981 11621 22015
rect 11621 21981 11655 22015
rect 11655 21981 11664 22015
rect 11612 21972 11664 21981
rect 12072 21972 12124 22024
rect 9496 21836 9548 21888
rect 12624 22015 12676 22024
rect 12624 21981 12633 22015
rect 12633 21981 12667 22015
rect 12667 21981 12676 22015
rect 12624 21972 12676 21981
rect 12716 22015 12768 22024
rect 12716 21981 12725 22015
rect 12725 21981 12759 22015
rect 12759 21981 12768 22015
rect 12716 21972 12768 21981
rect 12992 22015 13044 22024
rect 12992 21981 13001 22015
rect 13001 21981 13035 22015
rect 13035 21981 13044 22015
rect 12992 21972 13044 21981
rect 13084 22015 13136 22024
rect 13084 21981 13093 22015
rect 13093 21981 13127 22015
rect 13127 21981 13136 22015
rect 13084 21972 13136 21981
rect 13360 21947 13412 21956
rect 13360 21913 13369 21947
rect 13369 21913 13403 21947
rect 13403 21913 13412 21947
rect 13360 21904 13412 21913
rect 12716 21836 12768 21888
rect 13544 21972 13596 22024
rect 14004 21972 14056 22024
rect 14372 22015 14424 22024
rect 14372 21981 14381 22015
rect 14381 21981 14415 22015
rect 14415 21981 14424 22015
rect 14372 21972 14424 21981
rect 14740 22015 14792 22024
rect 14740 21981 14749 22015
rect 14749 21981 14783 22015
rect 14783 21981 14792 22015
rect 14740 21972 14792 21981
rect 16580 21972 16632 22024
rect 16948 21972 17000 22024
rect 17132 22015 17184 22024
rect 17132 21981 17142 22015
rect 17142 21981 17176 22015
rect 17176 21981 17184 22015
rect 17684 22040 17736 22092
rect 17132 21972 17184 21981
rect 18236 22176 18288 22228
rect 19340 22176 19392 22228
rect 18788 22108 18840 22160
rect 20168 22219 20220 22228
rect 20168 22185 20177 22219
rect 20177 22185 20211 22219
rect 20211 22185 20220 22219
rect 20168 22176 20220 22185
rect 19984 22151 20036 22160
rect 19984 22117 19993 22151
rect 19993 22117 20027 22151
rect 20027 22117 20036 22151
rect 21088 22176 21140 22228
rect 25320 22219 25372 22228
rect 25320 22185 25329 22219
rect 25329 22185 25363 22219
rect 25363 22185 25372 22219
rect 25320 22176 25372 22185
rect 26516 22176 26568 22228
rect 27160 22176 27212 22228
rect 27344 22219 27396 22228
rect 27344 22185 27353 22219
rect 27353 22185 27387 22219
rect 27387 22185 27396 22219
rect 27344 22176 27396 22185
rect 30012 22176 30064 22228
rect 31668 22176 31720 22228
rect 33140 22176 33192 22228
rect 34060 22176 34112 22228
rect 37740 22176 37792 22228
rect 37924 22176 37976 22228
rect 19984 22108 20036 22117
rect 18328 22040 18380 22092
rect 18604 22040 18656 22092
rect 19616 22040 19668 22092
rect 13728 21836 13780 21888
rect 17224 21836 17276 21888
rect 18236 22015 18288 22024
rect 18236 21981 18245 22015
rect 18245 21981 18279 22015
rect 18279 21981 18288 22015
rect 18236 21972 18288 21981
rect 19892 21972 19944 22024
rect 20260 22015 20312 22024
rect 20260 21981 20269 22015
rect 20269 21981 20303 22015
rect 20303 21981 20312 22015
rect 20260 21972 20312 21981
rect 17408 21947 17460 21956
rect 17408 21913 17417 21947
rect 17417 21913 17451 21947
rect 17451 21913 17460 21947
rect 17408 21904 17460 21913
rect 21548 22040 21600 22092
rect 21824 22108 21876 22160
rect 23480 22108 23532 22160
rect 32864 22108 32916 22160
rect 33232 22108 33284 22160
rect 37464 22108 37516 22160
rect 38660 22219 38712 22228
rect 38660 22185 38669 22219
rect 38669 22185 38703 22219
rect 38703 22185 38712 22219
rect 38660 22176 38712 22185
rect 20904 21972 20956 22024
rect 20996 21904 21048 21956
rect 21364 22015 21416 22024
rect 21364 21981 21373 22015
rect 21373 21981 21407 22015
rect 21407 21981 21416 22015
rect 21364 21972 21416 21981
rect 21548 21904 21600 21956
rect 22468 22015 22520 22024
rect 22468 21981 22477 22015
rect 22477 21981 22511 22015
rect 22511 21981 22520 22015
rect 22468 21972 22520 21981
rect 23848 22040 23900 22092
rect 25044 22083 25096 22092
rect 25044 22049 25053 22083
rect 25053 22049 25087 22083
rect 25087 22049 25096 22083
rect 25044 22040 25096 22049
rect 22928 22015 22980 22024
rect 22928 21981 22937 22015
rect 22937 21981 22971 22015
rect 22971 21981 22980 22015
rect 22928 21972 22980 21981
rect 24032 22015 24084 22024
rect 24032 21981 24041 22015
rect 24041 21981 24075 22015
rect 24075 21981 24084 22015
rect 24032 21972 24084 21981
rect 25044 21904 25096 21956
rect 25780 21972 25832 22024
rect 17684 21879 17736 21888
rect 17684 21845 17693 21879
rect 17693 21845 17727 21879
rect 17727 21845 17736 21879
rect 17684 21836 17736 21845
rect 17868 21836 17920 21888
rect 19340 21836 19392 21888
rect 19800 21836 19852 21888
rect 19892 21836 19944 21888
rect 21732 21836 21784 21888
rect 24400 21879 24452 21888
rect 24400 21845 24409 21879
rect 24409 21845 24443 21879
rect 24443 21845 24452 21879
rect 29644 22040 29696 22092
rect 30472 22040 30524 22092
rect 32128 22040 32180 22092
rect 32956 22040 33008 22092
rect 26148 21972 26200 22024
rect 27068 22015 27120 22024
rect 27068 21981 27077 22015
rect 27077 21981 27111 22015
rect 27111 21981 27120 22015
rect 27068 21972 27120 21981
rect 27528 22015 27580 22024
rect 27528 21981 27537 22015
rect 27537 21981 27571 22015
rect 27571 21981 27580 22015
rect 27528 21972 27580 21981
rect 30196 21972 30248 22024
rect 30564 22015 30616 22024
rect 30564 21981 30573 22015
rect 30573 21981 30607 22015
rect 30607 21981 30616 22015
rect 30564 21972 30616 21981
rect 32220 21972 32272 22024
rect 37924 22015 37976 22024
rect 37924 21981 37933 22015
rect 37933 21981 37967 22015
rect 37967 21981 37976 22015
rect 37924 21972 37976 21981
rect 24400 21836 24452 21845
rect 25964 21836 26016 21888
rect 26148 21836 26200 21888
rect 26240 21879 26292 21888
rect 26240 21845 26249 21879
rect 26249 21845 26283 21879
rect 26283 21845 26292 21879
rect 26240 21836 26292 21845
rect 26976 21879 27028 21888
rect 26976 21845 26985 21879
rect 26985 21845 27019 21879
rect 27019 21845 27028 21879
rect 26976 21836 27028 21845
rect 27620 21904 27672 21956
rect 28540 21836 28592 21888
rect 36544 21904 36596 21956
rect 39120 22015 39172 22024
rect 39120 21981 39129 22015
rect 39129 21981 39163 22015
rect 39163 21981 39172 22015
rect 39120 21972 39172 21981
rect 39304 22015 39356 22024
rect 39304 21981 39313 22015
rect 39313 21981 39347 22015
rect 39347 21981 39356 22015
rect 39304 21972 39356 21981
rect 39396 22015 39448 22024
rect 39396 21981 39405 22015
rect 39405 21981 39439 22015
rect 39439 21981 39448 22015
rect 39396 21972 39448 21981
rect 30012 21836 30064 21888
rect 32404 21836 32456 21888
rect 33968 21836 34020 21888
rect 34428 21836 34480 21888
rect 37280 21836 37332 21888
rect 38108 21836 38160 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 3332 21632 3384 21684
rect 4712 21632 4764 21684
rect 5356 21632 5408 21684
rect 5816 21632 5868 21684
rect 6092 21632 6144 21684
rect 3056 21564 3108 21616
rect 8576 21675 8628 21684
rect 8576 21641 8585 21675
rect 8585 21641 8619 21675
rect 8619 21641 8628 21675
rect 8576 21632 8628 21641
rect 10048 21632 10100 21684
rect 10416 21632 10468 21684
rect 11980 21632 12032 21684
rect 13084 21632 13136 21684
rect 17132 21632 17184 21684
rect 17776 21632 17828 21684
rect 20260 21632 20312 21684
rect 20352 21632 20404 21684
rect 3608 21539 3660 21548
rect 3608 21505 3617 21539
rect 3617 21505 3651 21539
rect 3651 21505 3660 21539
rect 3608 21496 3660 21505
rect 3700 21496 3752 21548
rect 3884 21539 3936 21548
rect 3884 21505 3893 21539
rect 3893 21505 3927 21539
rect 3927 21505 3936 21539
rect 3884 21496 3936 21505
rect 4436 21539 4488 21548
rect 4436 21505 4445 21539
rect 4445 21505 4479 21539
rect 4479 21505 4488 21539
rect 4436 21496 4488 21505
rect 5724 21539 5776 21548
rect 5724 21505 5733 21539
rect 5733 21505 5767 21539
rect 5767 21505 5776 21539
rect 5724 21496 5776 21505
rect 5908 21539 5960 21548
rect 5908 21505 5917 21539
rect 5917 21505 5951 21539
rect 5951 21505 5960 21539
rect 5908 21496 5960 21505
rect 11152 21564 11204 21616
rect 8208 21496 8260 21548
rect 8576 21496 8628 21548
rect 1492 21471 1544 21480
rect 1492 21437 1501 21471
rect 1501 21437 1535 21471
rect 1535 21437 1544 21471
rect 1492 21428 1544 21437
rect 5172 21428 5224 21480
rect 5080 21360 5132 21412
rect 5448 21428 5500 21480
rect 6828 21471 6880 21480
rect 6828 21437 6837 21471
rect 6837 21437 6871 21471
rect 6871 21437 6880 21471
rect 6828 21428 6880 21437
rect 7656 21428 7708 21480
rect 8392 21428 8444 21480
rect 10508 21496 10560 21548
rect 9864 21428 9916 21480
rect 5816 21403 5868 21412
rect 5816 21369 5825 21403
rect 5825 21369 5859 21403
rect 5859 21369 5868 21403
rect 5816 21360 5868 21369
rect 5632 21292 5684 21344
rect 6644 21292 6696 21344
rect 11428 21360 11480 21412
rect 8668 21335 8720 21344
rect 8668 21301 8677 21335
rect 8677 21301 8711 21335
rect 8711 21301 8720 21335
rect 8668 21292 8720 21301
rect 12624 21564 12676 21616
rect 12900 21539 12952 21548
rect 12900 21505 12909 21539
rect 12909 21505 12943 21539
rect 12943 21505 12952 21539
rect 12900 21496 12952 21505
rect 12992 21539 13044 21548
rect 12992 21505 13001 21539
rect 13001 21505 13035 21539
rect 13035 21505 13044 21539
rect 12992 21496 13044 21505
rect 13912 21564 13964 21616
rect 13360 21496 13412 21548
rect 14372 21496 14424 21548
rect 14740 21496 14792 21548
rect 20628 21564 20680 21616
rect 21364 21632 21416 21684
rect 22192 21632 22244 21684
rect 24400 21632 24452 21684
rect 25044 21632 25096 21684
rect 25780 21632 25832 21684
rect 26700 21632 26752 21684
rect 23388 21564 23440 21616
rect 25596 21564 25648 21616
rect 27068 21564 27120 21616
rect 33232 21632 33284 21684
rect 33784 21632 33836 21684
rect 27896 21564 27948 21616
rect 29000 21564 29052 21616
rect 31484 21564 31536 21616
rect 34152 21632 34204 21684
rect 34612 21632 34664 21684
rect 34796 21632 34848 21684
rect 13268 21428 13320 21480
rect 12716 21360 12768 21412
rect 16580 21428 16632 21480
rect 15108 21360 15160 21412
rect 17868 21496 17920 21548
rect 18788 21496 18840 21548
rect 20812 21496 20864 21548
rect 17040 21428 17092 21480
rect 18236 21428 18288 21480
rect 19432 21428 19484 21480
rect 17408 21360 17460 21412
rect 20260 21360 20312 21412
rect 21824 21496 21876 21548
rect 23756 21539 23808 21548
rect 23756 21505 23765 21539
rect 23765 21505 23799 21539
rect 23799 21505 23808 21539
rect 23756 21496 23808 21505
rect 24124 21496 24176 21548
rect 24400 21496 24452 21548
rect 24584 21496 24636 21548
rect 24860 21496 24912 21548
rect 25688 21496 25740 21548
rect 27252 21539 27304 21548
rect 27252 21505 27261 21539
rect 27261 21505 27295 21539
rect 27295 21505 27304 21539
rect 27252 21496 27304 21505
rect 27344 21539 27396 21548
rect 27344 21505 27354 21539
rect 27354 21505 27388 21539
rect 27388 21505 27396 21539
rect 27344 21496 27396 21505
rect 27712 21539 27764 21548
rect 27712 21505 27726 21539
rect 27726 21505 27760 21539
rect 27760 21505 27764 21539
rect 27712 21496 27764 21505
rect 27988 21539 28040 21548
rect 27988 21505 27997 21539
rect 27997 21505 28031 21539
rect 28031 21505 28040 21539
rect 27988 21496 28040 21505
rect 29092 21496 29144 21548
rect 31852 21539 31904 21548
rect 31852 21505 31861 21539
rect 31861 21505 31895 21539
rect 31895 21505 31904 21539
rect 31852 21496 31904 21505
rect 33048 21496 33100 21548
rect 35256 21564 35308 21616
rect 36268 21564 36320 21616
rect 22100 21360 22152 21412
rect 22192 21360 22244 21412
rect 24124 21360 24176 21412
rect 12992 21292 13044 21344
rect 14740 21292 14792 21344
rect 15016 21292 15068 21344
rect 17316 21292 17368 21344
rect 20628 21292 20680 21344
rect 21548 21292 21600 21344
rect 26608 21292 26660 21344
rect 32772 21360 32824 21412
rect 34612 21496 34664 21548
rect 33968 21428 34020 21480
rect 34888 21539 34940 21548
rect 34888 21505 34897 21539
rect 34897 21505 34931 21539
rect 34931 21505 34940 21539
rect 34888 21496 34940 21505
rect 35716 21539 35768 21548
rect 35716 21505 35725 21539
rect 35725 21505 35759 21539
rect 35759 21505 35768 21539
rect 35716 21496 35768 21505
rect 35900 21539 35952 21548
rect 35900 21505 35909 21539
rect 35909 21505 35943 21539
rect 35943 21505 35952 21539
rect 35900 21496 35952 21505
rect 35992 21496 36044 21548
rect 36452 21539 36504 21548
rect 36452 21505 36461 21539
rect 36461 21505 36495 21539
rect 36495 21505 36504 21539
rect 36452 21496 36504 21505
rect 36544 21539 36596 21548
rect 36544 21505 36553 21539
rect 36553 21505 36587 21539
rect 36587 21505 36596 21539
rect 36544 21496 36596 21505
rect 34428 21360 34480 21412
rect 38936 21428 38988 21480
rect 27988 21292 28040 21344
rect 28356 21335 28408 21344
rect 28356 21301 28365 21335
rect 28365 21301 28399 21335
rect 28399 21301 28408 21335
rect 28356 21292 28408 21301
rect 29736 21292 29788 21344
rect 30196 21292 30248 21344
rect 30932 21292 30984 21344
rect 31300 21292 31352 21344
rect 31668 21335 31720 21344
rect 31668 21301 31677 21335
rect 31677 21301 31711 21335
rect 31711 21301 31720 21335
rect 31668 21292 31720 21301
rect 32220 21292 32272 21344
rect 33232 21292 33284 21344
rect 35992 21292 36044 21344
rect 36176 21292 36228 21344
rect 37280 21292 37332 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 6276 21088 6328 21140
rect 6736 21088 6788 21140
rect 6184 21020 6236 21072
rect 2872 20952 2924 21004
rect 3332 20952 3384 21004
rect 5080 20995 5132 21004
rect 5080 20961 5089 20995
rect 5089 20961 5123 20995
rect 5123 20961 5132 20995
rect 5080 20952 5132 20961
rect 1584 20884 1636 20936
rect 4896 20927 4948 20936
rect 4896 20893 4905 20927
rect 4905 20893 4939 20927
rect 4939 20893 4948 20927
rect 4896 20884 4948 20893
rect 5448 20884 5500 20936
rect 2136 20859 2188 20868
rect 2136 20825 2145 20859
rect 2145 20825 2179 20859
rect 2179 20825 2188 20859
rect 2136 20816 2188 20825
rect 3792 20816 3844 20868
rect 5356 20816 5408 20868
rect 6000 20927 6052 20936
rect 6000 20893 6009 20927
rect 6009 20893 6043 20927
rect 6043 20893 6052 20927
rect 6000 20884 6052 20893
rect 6184 20927 6236 20936
rect 7012 21020 7064 21072
rect 7656 21131 7708 21140
rect 7656 21097 7665 21131
rect 7665 21097 7699 21131
rect 7699 21097 7708 21131
rect 7656 21088 7708 21097
rect 10232 21088 10284 21140
rect 10508 21088 10560 21140
rect 10876 21131 10928 21140
rect 10876 21097 10885 21131
rect 10885 21097 10919 21131
rect 10919 21097 10928 21131
rect 10876 21088 10928 21097
rect 6184 20893 6212 20927
rect 6212 20893 6236 20927
rect 6184 20884 6236 20893
rect 6736 20884 6788 20936
rect 8484 21020 8536 21072
rect 13268 21088 13320 21140
rect 15476 21088 15528 21140
rect 7472 20952 7524 21004
rect 9864 20952 9916 21004
rect 10140 20952 10192 21004
rect 7196 20927 7248 20936
rect 7196 20893 7205 20927
rect 7205 20893 7239 20927
rect 7239 20893 7248 20927
rect 7196 20884 7248 20893
rect 8668 20884 8720 20936
rect 10232 20927 10284 20936
rect 10232 20893 10241 20927
rect 10241 20893 10275 20927
rect 10275 20893 10284 20927
rect 10232 20884 10284 20893
rect 17132 21020 17184 21072
rect 18420 21020 18472 21072
rect 20812 21020 20864 21072
rect 21916 21020 21968 21072
rect 23204 21020 23256 21072
rect 29000 21088 29052 21140
rect 36452 21088 36504 21140
rect 11244 20952 11296 21004
rect 12900 20952 12952 21004
rect 3608 20791 3660 20800
rect 3608 20757 3617 20791
rect 3617 20757 3651 20791
rect 3651 20757 3660 20791
rect 3608 20748 3660 20757
rect 4436 20791 4488 20800
rect 4436 20757 4445 20791
rect 4445 20757 4479 20791
rect 4479 20757 4488 20791
rect 4436 20748 4488 20757
rect 7012 20859 7064 20868
rect 7012 20825 7021 20859
rect 7021 20825 7055 20859
rect 7055 20825 7064 20859
rect 7012 20816 7064 20825
rect 8576 20816 8628 20868
rect 8208 20748 8260 20800
rect 8300 20748 8352 20800
rect 10048 20748 10100 20800
rect 10600 20859 10652 20868
rect 10600 20825 10609 20859
rect 10609 20825 10643 20859
rect 10643 20825 10652 20859
rect 10600 20816 10652 20825
rect 11520 20816 11572 20868
rect 12256 20816 12308 20868
rect 12900 20816 12952 20868
rect 13820 20927 13872 20936
rect 13820 20893 13829 20927
rect 13829 20893 13863 20927
rect 13863 20893 13872 20927
rect 13820 20884 13872 20893
rect 15476 20952 15528 21004
rect 15660 20884 15712 20936
rect 17040 20927 17092 20936
rect 17040 20893 17049 20927
rect 17049 20893 17083 20927
rect 17083 20893 17092 20927
rect 17040 20884 17092 20893
rect 18236 20884 18288 20936
rect 18972 20952 19024 21004
rect 19800 20995 19852 21004
rect 19800 20961 19809 20995
rect 19809 20961 19843 20995
rect 19843 20961 19852 20995
rect 19800 20952 19852 20961
rect 25044 21020 25096 21072
rect 26240 21020 26292 21072
rect 29644 21020 29696 21072
rect 34796 21020 34848 21072
rect 35716 21020 35768 21072
rect 36084 21020 36136 21072
rect 37004 21131 37056 21140
rect 37004 21097 37013 21131
rect 37013 21097 37047 21131
rect 37047 21097 37056 21131
rect 37004 21088 37056 21097
rect 18512 20927 18564 20936
rect 18512 20893 18521 20927
rect 18521 20893 18555 20927
rect 18555 20893 18564 20927
rect 18512 20884 18564 20893
rect 18604 20816 18656 20868
rect 18788 20816 18840 20868
rect 19616 20884 19668 20936
rect 28356 20952 28408 21004
rect 20444 20927 20496 20936
rect 20444 20893 20453 20927
rect 20453 20893 20487 20927
rect 20487 20893 20496 20927
rect 20444 20884 20496 20893
rect 20628 20884 20680 20936
rect 23572 20927 23624 20936
rect 23572 20893 23581 20927
rect 23581 20893 23615 20927
rect 23615 20893 23624 20927
rect 23572 20884 23624 20893
rect 28908 20927 28960 20936
rect 28908 20893 28917 20927
rect 28917 20893 28951 20927
rect 28951 20893 28960 20927
rect 28908 20884 28960 20893
rect 29092 20884 29144 20936
rect 29920 20927 29972 20936
rect 29920 20893 29929 20927
rect 29929 20893 29963 20927
rect 29963 20893 29972 20927
rect 29920 20884 29972 20893
rect 30012 20884 30064 20936
rect 30472 20884 30524 20936
rect 12808 20791 12860 20800
rect 12808 20757 12817 20791
rect 12817 20757 12851 20791
rect 12851 20757 12860 20791
rect 12808 20748 12860 20757
rect 13912 20748 13964 20800
rect 14372 20748 14424 20800
rect 16120 20748 16172 20800
rect 16856 20748 16908 20800
rect 17408 20748 17460 20800
rect 18696 20748 18748 20800
rect 18972 20748 19024 20800
rect 20812 20859 20864 20868
rect 20812 20825 20821 20859
rect 20821 20825 20855 20859
rect 20855 20825 20864 20859
rect 20812 20816 20864 20825
rect 21732 20816 21784 20868
rect 23940 20816 23992 20868
rect 25964 20816 26016 20868
rect 27620 20816 27672 20868
rect 27712 20816 27764 20868
rect 28356 20816 28408 20868
rect 28724 20816 28776 20868
rect 20904 20748 20956 20800
rect 21548 20748 21600 20800
rect 21824 20748 21876 20800
rect 22008 20748 22060 20800
rect 26608 20791 26660 20800
rect 26608 20757 26617 20791
rect 26617 20757 26651 20791
rect 26651 20757 26660 20791
rect 26608 20748 26660 20757
rect 30288 20816 30340 20868
rect 32496 20995 32548 21004
rect 32496 20961 32505 20995
rect 32505 20961 32539 20995
rect 32539 20961 32548 20995
rect 32496 20952 32548 20961
rect 33048 20952 33100 21004
rect 31852 20884 31904 20936
rect 32220 20927 32272 20936
rect 32220 20893 32229 20927
rect 32229 20893 32263 20927
rect 32263 20893 32272 20927
rect 32220 20884 32272 20893
rect 32864 20884 32916 20936
rect 33784 20927 33836 20936
rect 33784 20893 33793 20927
rect 33793 20893 33827 20927
rect 33827 20893 33836 20927
rect 33784 20884 33836 20893
rect 34428 20884 34480 20936
rect 36176 20952 36228 21004
rect 37004 20952 37056 21004
rect 33876 20859 33928 20868
rect 33876 20825 33885 20859
rect 33885 20825 33919 20859
rect 33919 20825 33928 20859
rect 33876 20816 33928 20825
rect 36360 20884 36412 20936
rect 37280 20884 37332 20936
rect 38108 20884 38160 20936
rect 38476 20884 38528 20936
rect 36268 20816 36320 20868
rect 38292 20816 38344 20868
rect 38844 20816 38896 20868
rect 28816 20748 28868 20800
rect 29000 20748 29052 20800
rect 30472 20748 30524 20800
rect 33508 20791 33560 20800
rect 33508 20757 33517 20791
rect 33517 20757 33551 20791
rect 33551 20757 33560 20791
rect 33508 20748 33560 20757
rect 35256 20748 35308 20800
rect 35900 20791 35952 20800
rect 35900 20757 35909 20791
rect 35909 20757 35943 20791
rect 35943 20757 35952 20791
rect 35900 20748 35952 20757
rect 37280 20748 37332 20800
rect 38384 20748 38436 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 1584 20544 1636 20596
rect 3056 20451 3108 20460
rect 3056 20417 3065 20451
rect 3065 20417 3099 20451
rect 3099 20417 3108 20451
rect 3056 20408 3108 20417
rect 2780 20340 2832 20392
rect 3148 20383 3200 20392
rect 3148 20349 3157 20383
rect 3157 20349 3191 20383
rect 3191 20349 3200 20383
rect 3148 20340 3200 20349
rect 3332 20383 3384 20392
rect 3332 20349 3341 20383
rect 3341 20349 3375 20383
rect 3375 20349 3384 20383
rect 3332 20340 3384 20349
rect 5356 20544 5408 20596
rect 6000 20544 6052 20596
rect 6368 20587 6420 20596
rect 6368 20553 6377 20587
rect 6377 20553 6411 20587
rect 6411 20553 6420 20587
rect 6368 20544 6420 20553
rect 10600 20544 10652 20596
rect 11520 20544 11572 20596
rect 12808 20544 12860 20596
rect 3792 20476 3844 20528
rect 5540 20519 5592 20528
rect 5540 20485 5549 20519
rect 5549 20485 5583 20519
rect 5583 20485 5592 20519
rect 5540 20476 5592 20485
rect 5632 20519 5684 20528
rect 5632 20485 5641 20519
rect 5641 20485 5675 20519
rect 5675 20485 5684 20519
rect 5632 20476 5684 20485
rect 5264 20408 5316 20460
rect 5724 20451 5776 20460
rect 5724 20417 5733 20451
rect 5733 20417 5767 20451
rect 5767 20417 5776 20451
rect 5724 20408 5776 20417
rect 7104 20476 7156 20528
rect 9496 20476 9548 20528
rect 13084 20476 13136 20528
rect 2136 20272 2188 20324
rect 4436 20340 4488 20392
rect 5448 20340 5500 20392
rect 6644 20272 6696 20324
rect 12808 20408 12860 20460
rect 8576 20383 8628 20392
rect 8576 20349 8585 20383
rect 8585 20349 8619 20383
rect 8619 20349 8628 20383
rect 8576 20340 8628 20349
rect 9312 20340 9364 20392
rect 9864 20272 9916 20324
rect 19800 20544 19852 20596
rect 13912 20519 13964 20528
rect 13912 20485 13921 20519
rect 13921 20485 13955 20519
rect 13955 20485 13964 20519
rect 13912 20476 13964 20485
rect 14280 20476 14332 20528
rect 17132 20476 17184 20528
rect 18328 20476 18380 20528
rect 22008 20476 22060 20528
rect 23112 20476 23164 20528
rect 26424 20544 26476 20596
rect 25320 20476 25372 20528
rect 25872 20476 25924 20528
rect 13820 20408 13872 20460
rect 14188 20383 14240 20392
rect 14188 20349 14197 20383
rect 14197 20349 14231 20383
rect 14231 20349 14240 20383
rect 14188 20340 14240 20349
rect 14372 20451 14424 20460
rect 14372 20417 14381 20451
rect 14381 20417 14415 20451
rect 14415 20417 14424 20451
rect 14372 20408 14424 20417
rect 14464 20408 14516 20460
rect 15476 20451 15528 20460
rect 15476 20417 15485 20451
rect 15485 20417 15519 20451
rect 15519 20417 15528 20451
rect 15476 20408 15528 20417
rect 15568 20408 15620 20460
rect 15752 20451 15804 20460
rect 15752 20417 15761 20451
rect 15761 20417 15795 20451
rect 15795 20417 15804 20451
rect 15752 20408 15804 20417
rect 16304 20451 16356 20460
rect 16304 20417 16313 20451
rect 16313 20417 16347 20451
rect 16347 20417 16356 20451
rect 16304 20408 16356 20417
rect 16396 20408 16448 20460
rect 15016 20340 15068 20392
rect 15108 20383 15160 20392
rect 15108 20349 15117 20383
rect 15117 20349 15151 20383
rect 15151 20349 15160 20383
rect 15108 20340 15160 20349
rect 16580 20340 16632 20392
rect 17592 20340 17644 20392
rect 20628 20383 20680 20392
rect 20628 20349 20637 20383
rect 20637 20349 20671 20383
rect 20671 20349 20680 20383
rect 20628 20340 20680 20349
rect 21364 20408 21416 20460
rect 22284 20408 22336 20460
rect 22836 20451 22888 20460
rect 22836 20417 22845 20451
rect 22845 20417 22879 20451
rect 22879 20417 22888 20451
rect 22836 20408 22888 20417
rect 25044 20451 25096 20460
rect 25044 20417 25053 20451
rect 25053 20417 25087 20451
rect 25087 20417 25096 20451
rect 25044 20408 25096 20417
rect 23388 20340 23440 20392
rect 24952 20340 25004 20392
rect 25136 20340 25188 20392
rect 25688 20408 25740 20460
rect 26700 20408 26752 20460
rect 27344 20451 27396 20460
rect 27344 20417 27353 20451
rect 27353 20417 27387 20451
rect 27387 20417 27396 20451
rect 27344 20408 27396 20417
rect 27436 20451 27488 20460
rect 27436 20417 27445 20451
rect 27445 20417 27479 20451
rect 27479 20417 27488 20451
rect 27436 20408 27488 20417
rect 30472 20544 30524 20596
rect 28724 20519 28776 20528
rect 28724 20485 28733 20519
rect 28733 20485 28767 20519
rect 28767 20485 28776 20519
rect 28724 20476 28776 20485
rect 29736 20476 29788 20528
rect 13268 20315 13320 20324
rect 13268 20281 13277 20315
rect 13277 20281 13311 20315
rect 13311 20281 13320 20315
rect 13268 20272 13320 20281
rect 15660 20272 15712 20324
rect 23480 20272 23532 20324
rect 23664 20272 23716 20324
rect 25412 20272 25464 20324
rect 25964 20315 26016 20324
rect 25964 20281 25973 20315
rect 25973 20281 26007 20315
rect 26007 20281 26016 20315
rect 25964 20272 26016 20281
rect 4804 20204 4856 20256
rect 5632 20204 5684 20256
rect 6552 20204 6604 20256
rect 9956 20204 10008 20256
rect 12992 20204 13044 20256
rect 14096 20204 14148 20256
rect 18420 20247 18472 20256
rect 18420 20213 18429 20247
rect 18429 20213 18463 20247
rect 18463 20213 18472 20247
rect 18420 20204 18472 20213
rect 20444 20204 20496 20256
rect 23204 20204 23256 20256
rect 24308 20204 24360 20256
rect 25320 20204 25372 20256
rect 25504 20247 25556 20256
rect 25504 20213 25513 20247
rect 25513 20213 25547 20247
rect 25547 20213 25556 20247
rect 25504 20204 25556 20213
rect 27068 20340 27120 20392
rect 27712 20451 27764 20460
rect 27712 20417 27721 20451
rect 27721 20417 27755 20451
rect 27755 20417 27764 20451
rect 27712 20408 27764 20417
rect 28264 20451 28316 20460
rect 28264 20417 28273 20451
rect 28273 20417 28307 20451
rect 28307 20417 28316 20451
rect 28264 20408 28316 20417
rect 29000 20451 29052 20460
rect 29000 20417 29009 20451
rect 29009 20417 29043 20451
rect 29043 20417 29052 20451
rect 29000 20408 29052 20417
rect 29828 20451 29880 20460
rect 29828 20417 29837 20451
rect 29837 20417 29871 20451
rect 29871 20417 29880 20451
rect 29828 20408 29880 20417
rect 30012 20408 30064 20460
rect 33968 20544 34020 20596
rect 30840 20476 30892 20528
rect 31760 20476 31812 20528
rect 36544 20476 36596 20528
rect 38016 20476 38068 20528
rect 38384 20519 38436 20528
rect 38384 20485 38393 20519
rect 38393 20485 38427 20519
rect 38427 20485 38436 20519
rect 38384 20476 38436 20485
rect 27804 20340 27856 20392
rect 28080 20383 28132 20392
rect 28080 20349 28089 20383
rect 28089 20349 28123 20383
rect 28123 20349 28132 20383
rect 28080 20340 28132 20349
rect 28632 20383 28684 20392
rect 28632 20349 28641 20383
rect 28641 20349 28675 20383
rect 28675 20349 28684 20383
rect 28632 20340 28684 20349
rect 27528 20272 27580 20324
rect 31484 20451 31536 20460
rect 31484 20417 31493 20451
rect 31493 20417 31527 20451
rect 31527 20417 31536 20451
rect 31484 20408 31536 20417
rect 31576 20451 31628 20460
rect 31576 20417 31585 20451
rect 31585 20417 31619 20451
rect 31619 20417 31628 20451
rect 31576 20408 31628 20417
rect 31852 20408 31904 20460
rect 32036 20408 32088 20460
rect 32496 20451 32548 20460
rect 32496 20417 32505 20451
rect 32505 20417 32539 20451
rect 32539 20417 32548 20451
rect 32496 20408 32548 20417
rect 32588 20408 32640 20460
rect 32864 20451 32916 20460
rect 32864 20417 32873 20451
rect 32873 20417 32907 20451
rect 32907 20417 32916 20451
rect 32864 20408 32916 20417
rect 33600 20408 33652 20460
rect 34704 20408 34756 20460
rect 38108 20451 38160 20460
rect 38108 20417 38117 20451
rect 38117 20417 38151 20451
rect 38151 20417 38160 20451
rect 38108 20408 38160 20417
rect 31208 20383 31260 20392
rect 31208 20349 31217 20383
rect 31217 20349 31251 20383
rect 31251 20349 31260 20383
rect 31208 20340 31260 20349
rect 31760 20340 31812 20392
rect 33232 20340 33284 20392
rect 33784 20340 33836 20392
rect 37096 20340 37148 20392
rect 37648 20340 37700 20392
rect 38292 20408 38344 20460
rect 30932 20272 30984 20324
rect 31484 20272 31536 20324
rect 34428 20272 34480 20324
rect 35992 20272 36044 20324
rect 38016 20272 38068 20324
rect 27804 20204 27856 20256
rect 27988 20247 28040 20256
rect 27988 20213 27997 20247
rect 27997 20213 28031 20247
rect 28031 20213 28040 20247
rect 27988 20204 28040 20213
rect 28448 20247 28500 20256
rect 28448 20213 28457 20247
rect 28457 20213 28491 20247
rect 28491 20213 28500 20247
rect 28448 20204 28500 20213
rect 29828 20204 29880 20256
rect 30656 20204 30708 20256
rect 30840 20204 30892 20256
rect 31576 20204 31628 20256
rect 31760 20204 31812 20256
rect 32220 20204 32272 20256
rect 32864 20204 32916 20256
rect 33048 20247 33100 20256
rect 33048 20213 33057 20247
rect 33057 20213 33091 20247
rect 33091 20213 33100 20247
rect 33048 20204 33100 20213
rect 33968 20204 34020 20256
rect 35256 20204 35308 20256
rect 39304 20204 39356 20256
rect 39580 20204 39632 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 3056 20000 3108 20052
rect 5816 20000 5868 20052
rect 6736 20043 6788 20052
rect 6736 20009 6745 20043
rect 6745 20009 6779 20043
rect 6779 20009 6788 20043
rect 6736 20000 6788 20009
rect 7104 20000 7156 20052
rect 7840 20000 7892 20052
rect 8024 20043 8076 20052
rect 8024 20009 8033 20043
rect 8033 20009 8067 20043
rect 8067 20009 8076 20043
rect 8024 20000 8076 20009
rect 9312 20043 9364 20052
rect 9312 20009 9321 20043
rect 9321 20009 9355 20043
rect 9355 20009 9364 20043
rect 9312 20000 9364 20009
rect 10232 20000 10284 20052
rect 13544 20043 13596 20052
rect 13544 20009 13553 20043
rect 13553 20009 13587 20043
rect 13587 20009 13596 20043
rect 13544 20000 13596 20009
rect 13636 20000 13688 20052
rect 14188 20000 14240 20052
rect 14464 20043 14516 20052
rect 14464 20009 14473 20043
rect 14473 20009 14507 20043
rect 14507 20009 14516 20043
rect 14464 20000 14516 20009
rect 5724 19932 5776 19984
rect 6368 19932 6420 19984
rect 6460 19932 6512 19984
rect 3608 19864 3660 19916
rect 3424 19796 3476 19848
rect 5632 19796 5684 19848
rect 5724 19839 5776 19848
rect 5724 19805 5733 19839
rect 5733 19805 5767 19839
rect 5767 19805 5776 19839
rect 5724 19796 5776 19805
rect 6184 19839 6236 19848
rect 6184 19805 6193 19839
rect 6193 19805 6227 19839
rect 6227 19805 6236 19839
rect 6184 19796 6236 19805
rect 6368 19839 6420 19848
rect 6368 19805 6377 19839
rect 6377 19805 6411 19839
rect 6411 19805 6420 19839
rect 6368 19796 6420 19805
rect 6736 19796 6788 19848
rect 7104 19864 7156 19916
rect 3884 19660 3936 19712
rect 5264 19660 5316 19712
rect 6644 19728 6696 19780
rect 7840 19839 7892 19848
rect 7840 19805 7849 19839
rect 7849 19805 7883 19839
rect 7883 19805 7892 19839
rect 7840 19796 7892 19805
rect 8668 19864 8720 19916
rect 9772 19907 9824 19916
rect 9772 19873 9781 19907
rect 9781 19873 9815 19907
rect 9815 19873 9824 19907
rect 9772 19864 9824 19873
rect 9864 19907 9916 19916
rect 9864 19873 9873 19907
rect 9873 19873 9907 19907
rect 9907 19873 9916 19907
rect 9864 19864 9916 19873
rect 10692 19932 10744 19984
rect 10876 19932 10928 19984
rect 13360 19932 13412 19984
rect 15384 20000 15436 20052
rect 20168 20000 20220 20052
rect 12532 19907 12584 19916
rect 9956 19796 10008 19848
rect 12532 19873 12541 19907
rect 12541 19873 12575 19907
rect 12575 19873 12584 19907
rect 12532 19864 12584 19873
rect 12716 19864 12768 19916
rect 10692 19839 10744 19848
rect 10692 19805 10701 19839
rect 10701 19805 10735 19839
rect 10735 19805 10744 19839
rect 10692 19796 10744 19805
rect 12624 19796 12676 19848
rect 12900 19796 12952 19848
rect 12992 19839 13044 19848
rect 12992 19805 13001 19839
rect 13001 19805 13035 19839
rect 13035 19805 13044 19839
rect 12992 19796 13044 19805
rect 15476 19932 15528 19984
rect 17040 19932 17092 19984
rect 14924 19839 14976 19848
rect 14924 19805 14969 19839
rect 14969 19805 14976 19839
rect 14924 19796 14976 19805
rect 15292 19796 15344 19848
rect 15384 19839 15436 19848
rect 15384 19805 15393 19839
rect 15393 19805 15427 19839
rect 15427 19805 15436 19839
rect 15384 19796 15436 19805
rect 19708 19864 19760 19916
rect 21180 19932 21232 19984
rect 21272 19975 21324 19984
rect 21272 19941 21281 19975
rect 21281 19941 21315 19975
rect 21315 19941 21324 19975
rect 21272 19932 21324 19941
rect 21364 19975 21416 19984
rect 21364 19941 21373 19975
rect 21373 19941 21407 19975
rect 21407 19941 21416 19975
rect 21364 19932 21416 19941
rect 22836 20043 22888 20052
rect 22836 20009 22845 20043
rect 22845 20009 22879 20043
rect 22879 20009 22888 20043
rect 22836 20000 22888 20009
rect 23112 20000 23164 20052
rect 22100 19932 22152 19984
rect 23204 19975 23256 19984
rect 23204 19941 23213 19975
rect 23213 19941 23247 19975
rect 23247 19941 23256 19975
rect 23204 19932 23256 19941
rect 25136 20000 25188 20052
rect 25320 20043 25372 20052
rect 25320 20009 25329 20043
rect 25329 20009 25363 20043
rect 25363 20009 25372 20043
rect 25320 20000 25372 20009
rect 25412 20000 25464 20052
rect 26056 20043 26108 20052
rect 26056 20009 26065 20043
rect 26065 20009 26099 20043
rect 26099 20009 26108 20043
rect 26056 20000 26108 20009
rect 26700 20000 26752 20052
rect 27712 20000 27764 20052
rect 22836 19864 22888 19916
rect 23388 19864 23440 19916
rect 10416 19771 10468 19780
rect 10416 19737 10425 19771
rect 10425 19737 10459 19771
rect 10459 19737 10468 19771
rect 10416 19728 10468 19737
rect 7196 19703 7248 19712
rect 7196 19669 7205 19703
rect 7205 19669 7239 19703
rect 7239 19669 7248 19703
rect 7196 19660 7248 19669
rect 8116 19703 8168 19712
rect 8116 19669 8125 19703
rect 8125 19669 8159 19703
rect 8159 19669 8168 19703
rect 8116 19660 8168 19669
rect 10048 19660 10100 19712
rect 13820 19728 13872 19780
rect 13544 19660 13596 19712
rect 14372 19771 14424 19780
rect 14372 19737 14381 19771
rect 14381 19737 14415 19771
rect 14415 19737 14424 19771
rect 14372 19728 14424 19737
rect 14464 19728 14516 19780
rect 15660 19839 15712 19848
rect 15660 19805 15669 19839
rect 15669 19805 15703 19839
rect 15703 19805 15712 19839
rect 15660 19796 15712 19805
rect 14280 19660 14332 19712
rect 15016 19660 15068 19712
rect 15292 19660 15344 19712
rect 18696 19796 18748 19848
rect 19524 19796 19576 19848
rect 20076 19796 20128 19848
rect 17592 19728 17644 19780
rect 19340 19728 19392 19780
rect 19616 19728 19668 19780
rect 20536 19839 20588 19848
rect 20536 19805 20545 19839
rect 20545 19805 20579 19839
rect 20579 19805 20588 19839
rect 20536 19796 20588 19805
rect 20628 19839 20680 19848
rect 20628 19805 20637 19839
rect 20637 19805 20671 19839
rect 20671 19805 20680 19839
rect 20628 19796 20680 19805
rect 20812 19839 20864 19848
rect 20812 19805 20821 19839
rect 20821 19805 20855 19839
rect 20855 19805 20864 19839
rect 20812 19796 20864 19805
rect 21272 19796 21324 19848
rect 21732 19839 21784 19848
rect 21732 19805 21741 19839
rect 21741 19805 21775 19839
rect 21775 19805 21784 19839
rect 21732 19796 21784 19805
rect 21824 19839 21876 19848
rect 21824 19805 21833 19839
rect 21833 19805 21867 19839
rect 21867 19805 21876 19839
rect 21824 19796 21876 19805
rect 22284 19796 22336 19848
rect 22744 19796 22796 19848
rect 23112 19796 23164 19848
rect 23572 19796 23624 19848
rect 25780 19932 25832 19984
rect 26240 19932 26292 19984
rect 28264 19932 28316 19984
rect 29920 19932 29972 19984
rect 30104 19932 30156 19984
rect 33692 19932 33744 19984
rect 34428 19932 34480 19984
rect 24492 19796 24544 19848
rect 25044 19864 25096 19916
rect 22192 19728 22244 19780
rect 25136 19771 25188 19780
rect 25136 19737 25145 19771
rect 25145 19737 25179 19771
rect 25179 19737 25188 19771
rect 25136 19728 25188 19737
rect 25504 19728 25556 19780
rect 17408 19660 17460 19712
rect 18880 19660 18932 19712
rect 22376 19660 22428 19712
rect 23480 19660 23532 19712
rect 23756 19660 23808 19712
rect 24308 19660 24360 19712
rect 24584 19660 24636 19712
rect 28448 19864 28500 19916
rect 26608 19796 26660 19848
rect 27252 19796 27304 19848
rect 27528 19796 27580 19848
rect 26516 19771 26568 19780
rect 26516 19737 26525 19771
rect 26525 19737 26559 19771
rect 26559 19737 26568 19771
rect 26516 19728 26568 19737
rect 27160 19728 27212 19780
rect 27896 19796 27948 19848
rect 28908 19796 28960 19848
rect 31208 19796 31260 19848
rect 31392 19864 31444 19916
rect 33876 19864 33928 19916
rect 35164 19864 35216 19916
rect 35348 19864 35400 19916
rect 37924 19864 37976 19916
rect 31484 19839 31536 19848
rect 31484 19805 31493 19839
rect 31493 19805 31527 19839
rect 31527 19805 31536 19839
rect 31484 19796 31536 19805
rect 31668 19796 31720 19848
rect 33048 19796 33100 19848
rect 36452 19796 36504 19848
rect 36912 19839 36964 19848
rect 36912 19805 36922 19839
rect 36922 19805 36956 19839
rect 36956 19805 36964 19839
rect 36912 19796 36964 19805
rect 37280 19839 37332 19848
rect 37280 19805 37294 19839
rect 37294 19805 37328 19839
rect 37328 19805 37332 19839
rect 37280 19796 37332 19805
rect 38016 19796 38068 19848
rect 27712 19728 27764 19780
rect 27988 19728 28040 19780
rect 30472 19728 30524 19780
rect 33324 19728 33376 19780
rect 36176 19728 36228 19780
rect 36360 19728 36412 19780
rect 37188 19771 37240 19780
rect 37188 19737 37197 19771
rect 37197 19737 37231 19771
rect 37231 19737 37240 19771
rect 37188 19728 37240 19737
rect 38108 19728 38160 19780
rect 39212 19796 39264 19848
rect 39672 19728 39724 19780
rect 28724 19660 28776 19712
rect 31576 19660 31628 19712
rect 32404 19660 32456 19712
rect 33692 19660 33744 19712
rect 33876 19660 33928 19712
rect 37372 19660 37424 19712
rect 37464 19703 37516 19712
rect 37464 19669 37473 19703
rect 37473 19669 37507 19703
rect 37507 19669 37516 19703
rect 37464 19660 37516 19669
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 3424 19499 3476 19508
rect 3424 19465 3433 19499
rect 3433 19465 3467 19499
rect 3467 19465 3476 19499
rect 3424 19456 3476 19465
rect 3884 19499 3936 19508
rect 3884 19465 3893 19499
rect 3893 19465 3927 19499
rect 3927 19465 3936 19499
rect 3884 19456 3936 19465
rect 4804 19456 4856 19508
rect 5172 19456 5224 19508
rect 6828 19456 6880 19508
rect 3516 19388 3568 19440
rect 5724 19388 5776 19440
rect 3056 19320 3108 19372
rect 5540 19320 5592 19372
rect 1584 19252 1636 19304
rect 4068 19295 4120 19304
rect 4068 19261 4077 19295
rect 4077 19261 4111 19295
rect 4111 19261 4120 19295
rect 4068 19252 4120 19261
rect 4620 19252 4672 19304
rect 4896 19295 4948 19304
rect 4896 19261 4905 19295
rect 4905 19261 4939 19295
rect 4939 19261 4948 19295
rect 4896 19252 4948 19261
rect 5448 19252 5500 19304
rect 5908 19252 5960 19304
rect 6644 19320 6696 19372
rect 8576 19456 8628 19508
rect 8668 19499 8720 19508
rect 8668 19465 8677 19499
rect 8677 19465 8711 19499
rect 8711 19465 8720 19499
rect 8668 19456 8720 19465
rect 10416 19456 10468 19508
rect 7472 19388 7524 19440
rect 9496 19388 9548 19440
rect 8576 19320 8628 19372
rect 12532 19456 12584 19508
rect 14280 19499 14332 19508
rect 14280 19465 14289 19499
rect 14289 19465 14323 19499
rect 14323 19465 14332 19499
rect 14280 19456 14332 19465
rect 15016 19456 15068 19508
rect 15292 19456 15344 19508
rect 15568 19456 15620 19508
rect 17132 19499 17184 19508
rect 17132 19465 17141 19499
rect 17141 19465 17175 19499
rect 17175 19465 17184 19499
rect 17132 19456 17184 19465
rect 17408 19456 17460 19508
rect 6736 19252 6788 19304
rect 7656 19252 7708 19304
rect 9496 19252 9548 19304
rect 14096 19320 14148 19372
rect 14372 19320 14424 19372
rect 15752 19388 15804 19440
rect 15292 19320 15344 19372
rect 15844 19320 15896 19372
rect 16212 19363 16264 19372
rect 16212 19329 16221 19363
rect 16221 19329 16255 19363
rect 16255 19329 16264 19363
rect 16212 19320 16264 19329
rect 16396 19363 16448 19372
rect 16396 19329 16405 19363
rect 16405 19329 16439 19363
rect 16439 19329 16448 19363
rect 16396 19320 16448 19329
rect 18052 19388 18104 19440
rect 18696 19388 18748 19440
rect 17592 19363 17644 19372
rect 17592 19329 17596 19363
rect 17596 19329 17630 19363
rect 17630 19329 17644 19363
rect 16764 19252 16816 19304
rect 17592 19320 17644 19329
rect 17776 19363 17828 19372
rect 17776 19329 17785 19363
rect 17785 19329 17819 19363
rect 17819 19329 17828 19363
rect 17776 19320 17828 19329
rect 18328 19320 18380 19372
rect 18512 19363 18564 19372
rect 18512 19329 18521 19363
rect 18521 19329 18555 19363
rect 18555 19329 18564 19363
rect 18512 19320 18564 19329
rect 20812 19456 20864 19508
rect 21364 19456 21416 19508
rect 21640 19456 21692 19508
rect 21824 19456 21876 19508
rect 21916 19456 21968 19508
rect 22376 19456 22428 19508
rect 23296 19456 23348 19508
rect 19248 19320 19300 19372
rect 21272 19320 21324 19372
rect 4988 19184 5040 19236
rect 14188 19184 14240 19236
rect 14740 19184 14792 19236
rect 4620 19116 4672 19168
rect 4712 19116 4764 19168
rect 10600 19159 10652 19168
rect 10600 19125 10609 19159
rect 10609 19125 10643 19159
rect 10643 19125 10652 19159
rect 10600 19116 10652 19125
rect 15936 19116 15988 19168
rect 16856 19227 16908 19236
rect 16856 19193 16865 19227
rect 16865 19193 16899 19227
rect 16899 19193 16908 19227
rect 16856 19184 16908 19193
rect 21640 19252 21692 19304
rect 22928 19388 22980 19440
rect 23480 19388 23532 19440
rect 22192 19320 22244 19372
rect 22836 19320 22888 19372
rect 23388 19320 23440 19372
rect 23572 19363 23624 19372
rect 23572 19329 23581 19363
rect 23581 19329 23615 19363
rect 23615 19329 23624 19363
rect 23572 19320 23624 19329
rect 23756 19295 23808 19304
rect 23756 19261 23765 19295
rect 23765 19261 23799 19295
rect 23799 19261 23808 19295
rect 25504 19456 25556 19508
rect 27252 19456 27304 19508
rect 27344 19456 27396 19508
rect 24492 19388 24544 19440
rect 29000 19456 29052 19508
rect 30288 19499 30340 19508
rect 30288 19465 30297 19499
rect 30297 19465 30331 19499
rect 30331 19465 30340 19499
rect 30288 19456 30340 19465
rect 31024 19456 31076 19508
rect 27620 19431 27672 19440
rect 27620 19397 27647 19431
rect 27647 19397 27672 19431
rect 27620 19388 27672 19397
rect 27804 19431 27856 19440
rect 27804 19397 27813 19431
rect 27813 19397 27847 19431
rect 27847 19397 27856 19431
rect 31668 19456 31720 19508
rect 27804 19388 27856 19397
rect 25136 19320 25188 19372
rect 25412 19320 25464 19372
rect 26332 19320 26384 19372
rect 28724 19363 28776 19372
rect 28724 19329 28733 19363
rect 28733 19329 28767 19363
rect 28767 19329 28776 19363
rect 28724 19320 28776 19329
rect 29368 19320 29420 19372
rect 29460 19320 29512 19372
rect 29920 19363 29972 19372
rect 29920 19329 29929 19363
rect 29929 19329 29963 19363
rect 29963 19329 29972 19363
rect 29920 19320 29972 19329
rect 30012 19320 30064 19372
rect 23756 19252 23808 19261
rect 29092 19295 29144 19304
rect 29092 19261 29101 19295
rect 29101 19261 29135 19295
rect 29135 19261 29144 19295
rect 29092 19252 29144 19261
rect 30104 19295 30156 19304
rect 30104 19261 30113 19295
rect 30113 19261 30147 19295
rect 30147 19261 30156 19295
rect 30104 19252 30156 19261
rect 30196 19295 30248 19304
rect 30196 19261 30205 19295
rect 30205 19261 30239 19295
rect 30239 19261 30248 19295
rect 30196 19252 30248 19261
rect 30840 19320 30892 19372
rect 31024 19320 31076 19372
rect 32588 19388 32640 19440
rect 33324 19388 33376 19440
rect 33968 19431 34020 19440
rect 33968 19397 33985 19431
rect 33985 19397 34020 19431
rect 33968 19388 34020 19397
rect 34152 19431 34204 19440
rect 34152 19397 34161 19431
rect 34161 19397 34195 19431
rect 34195 19397 34204 19431
rect 34152 19388 34204 19397
rect 34612 19388 34664 19440
rect 21824 19227 21876 19236
rect 21824 19193 21833 19227
rect 21833 19193 21867 19227
rect 21867 19193 21876 19227
rect 21824 19184 21876 19193
rect 27712 19184 27764 19236
rect 18328 19116 18380 19168
rect 27252 19116 27304 19168
rect 28264 19116 28316 19168
rect 29276 19184 29328 19236
rect 29644 19184 29696 19236
rect 34060 19363 34112 19372
rect 34060 19329 34069 19363
rect 34069 19329 34103 19363
rect 34103 19329 34112 19363
rect 34060 19320 34112 19329
rect 34244 19363 34296 19372
rect 34244 19329 34253 19363
rect 34253 19329 34287 19363
rect 34287 19329 34296 19363
rect 34244 19320 34296 19329
rect 34796 19456 34848 19508
rect 35532 19456 35584 19508
rect 35808 19456 35860 19508
rect 36360 19388 36412 19440
rect 34980 19363 35032 19372
rect 34980 19329 34989 19363
rect 34989 19329 35023 19363
rect 35023 19329 35032 19363
rect 34980 19320 35032 19329
rect 35164 19320 35216 19372
rect 34888 19295 34940 19304
rect 34888 19261 34897 19295
rect 34897 19261 34931 19295
rect 34931 19261 34940 19295
rect 34888 19252 34940 19261
rect 35440 19320 35492 19372
rect 35808 19363 35860 19372
rect 35808 19329 35817 19363
rect 35817 19329 35851 19363
rect 35851 19329 35860 19363
rect 35808 19320 35860 19329
rect 36176 19320 36228 19372
rect 36452 19363 36504 19372
rect 36452 19329 36461 19363
rect 36461 19329 36495 19363
rect 36495 19329 36504 19363
rect 36452 19320 36504 19329
rect 37188 19456 37240 19508
rect 38108 19456 38160 19508
rect 39028 19456 39080 19508
rect 39488 19456 39540 19508
rect 30840 19184 30892 19236
rect 29920 19116 29972 19168
rect 30104 19116 30156 19168
rect 31208 19159 31260 19168
rect 31208 19125 31217 19159
rect 31217 19125 31251 19159
rect 31251 19125 31260 19159
rect 31208 19116 31260 19125
rect 34060 19184 34112 19236
rect 34428 19184 34480 19236
rect 36176 19184 36228 19236
rect 39212 19252 39264 19304
rect 33968 19116 34020 19168
rect 35808 19116 35860 19168
rect 35900 19116 35952 19168
rect 36544 19116 36596 19168
rect 36820 19116 36872 19168
rect 38752 19116 38804 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 4896 18912 4948 18964
rect 5080 18912 5132 18964
rect 3792 18844 3844 18896
rect 1584 18819 1636 18828
rect 1584 18785 1593 18819
rect 1593 18785 1627 18819
rect 1627 18785 1636 18819
rect 1584 18776 1636 18785
rect 3056 18776 3108 18828
rect 4068 18776 4120 18828
rect 4436 18776 4488 18828
rect 5080 18776 5132 18828
rect 5172 18819 5224 18828
rect 5172 18785 5181 18819
rect 5181 18785 5215 18819
rect 5215 18785 5224 18819
rect 5172 18776 5224 18785
rect 7656 18955 7708 18964
rect 7656 18921 7665 18955
rect 7665 18921 7699 18955
rect 7699 18921 7708 18955
rect 7656 18912 7708 18921
rect 9496 18955 9548 18964
rect 9496 18921 9505 18955
rect 9505 18921 9539 18955
rect 9539 18921 9548 18955
rect 9496 18912 9548 18921
rect 12624 18955 12676 18964
rect 12624 18921 12633 18955
rect 12633 18921 12667 18955
rect 12667 18921 12676 18955
rect 12624 18912 12676 18921
rect 15844 18955 15896 18964
rect 15844 18921 15853 18955
rect 15853 18921 15887 18955
rect 15887 18921 15896 18955
rect 15844 18912 15896 18921
rect 20628 18912 20680 18964
rect 21640 18955 21692 18964
rect 21640 18921 21649 18955
rect 21649 18921 21683 18955
rect 21683 18921 21692 18955
rect 21640 18912 21692 18921
rect 23388 18912 23440 18964
rect 20260 18844 20312 18896
rect 1860 18683 1912 18692
rect 1860 18649 1869 18683
rect 1869 18649 1903 18683
rect 1903 18649 1912 18683
rect 1860 18640 1912 18649
rect 4712 18751 4764 18760
rect 4712 18717 4721 18751
rect 4721 18717 4755 18751
rect 4755 18717 4764 18751
rect 4712 18708 4764 18717
rect 4988 18708 5040 18760
rect 7012 18776 7064 18828
rect 11152 18776 11204 18828
rect 11244 18776 11296 18828
rect 8116 18708 8168 18760
rect 8760 18708 8812 18760
rect 9404 18751 9456 18760
rect 9404 18717 9413 18751
rect 9413 18717 9447 18751
rect 9447 18717 9456 18751
rect 9404 18708 9456 18717
rect 10600 18708 10652 18760
rect 3240 18640 3292 18692
rect 3792 18572 3844 18624
rect 4068 18572 4120 18624
rect 5448 18683 5500 18692
rect 5448 18649 5457 18683
rect 5457 18649 5491 18683
rect 5491 18649 5500 18683
rect 5448 18640 5500 18649
rect 12256 18708 12308 18760
rect 11152 18683 11204 18692
rect 11152 18649 11161 18683
rect 11161 18649 11195 18683
rect 11195 18649 11204 18683
rect 11152 18640 11204 18649
rect 12624 18708 12676 18760
rect 15936 18751 15988 18760
rect 15936 18717 15945 18751
rect 15945 18717 15979 18751
rect 15979 18717 15988 18751
rect 15936 18708 15988 18717
rect 14096 18640 14148 18692
rect 20352 18751 20404 18760
rect 20352 18717 20361 18751
rect 20361 18717 20395 18751
rect 20395 18717 20404 18751
rect 20352 18708 20404 18717
rect 23112 18844 23164 18896
rect 23756 18844 23808 18896
rect 24952 18912 25004 18964
rect 26516 18912 26568 18964
rect 26792 18912 26844 18964
rect 25228 18844 25280 18896
rect 26240 18844 26292 18896
rect 27436 18955 27488 18964
rect 27436 18921 27445 18955
rect 27445 18921 27479 18955
rect 27479 18921 27488 18955
rect 27436 18912 27488 18921
rect 27620 18955 27672 18964
rect 27620 18921 27629 18955
rect 27629 18921 27663 18955
rect 27663 18921 27672 18955
rect 27620 18912 27672 18921
rect 28724 18912 28776 18964
rect 30564 18912 30616 18964
rect 32772 18912 32824 18964
rect 35532 18912 35584 18964
rect 36544 18912 36596 18964
rect 27804 18844 27856 18896
rect 28172 18887 28224 18896
rect 28172 18853 28181 18887
rect 28181 18853 28215 18887
rect 28215 18853 28224 18887
rect 28172 18844 28224 18853
rect 29276 18887 29328 18896
rect 29276 18853 29285 18887
rect 29285 18853 29319 18887
rect 29319 18853 29328 18887
rect 29276 18844 29328 18853
rect 31024 18844 31076 18896
rect 31668 18844 31720 18896
rect 34612 18844 34664 18896
rect 35992 18844 36044 18896
rect 21272 18776 21324 18828
rect 24584 18776 24636 18828
rect 20720 18708 20772 18760
rect 21640 18708 21692 18760
rect 21824 18708 21876 18760
rect 22008 18751 22060 18760
rect 22008 18717 22017 18751
rect 22017 18717 22051 18751
rect 22051 18717 22060 18751
rect 22008 18708 22060 18717
rect 19708 18640 19760 18692
rect 7196 18572 7248 18624
rect 7748 18572 7800 18624
rect 8116 18615 8168 18624
rect 8116 18581 8125 18615
rect 8125 18581 8159 18615
rect 8159 18581 8168 18615
rect 8116 18572 8168 18581
rect 9864 18572 9916 18624
rect 9956 18615 10008 18624
rect 9956 18581 9965 18615
rect 9965 18581 9999 18615
rect 9999 18581 10008 18615
rect 9956 18572 10008 18581
rect 10048 18572 10100 18624
rect 12624 18572 12676 18624
rect 12716 18615 12768 18624
rect 12716 18581 12725 18615
rect 12725 18581 12759 18615
rect 12759 18581 12768 18615
rect 12716 18572 12768 18581
rect 17960 18572 18012 18624
rect 21640 18572 21692 18624
rect 23204 18708 23256 18760
rect 24400 18708 24452 18760
rect 24952 18708 25004 18760
rect 25780 18751 25832 18760
rect 25780 18717 25789 18751
rect 25789 18717 25823 18751
rect 25823 18717 25832 18751
rect 25780 18708 25832 18717
rect 22192 18572 22244 18624
rect 24584 18572 24636 18624
rect 25136 18615 25188 18624
rect 25136 18581 25163 18615
rect 25163 18581 25188 18615
rect 25136 18572 25188 18581
rect 25412 18640 25464 18692
rect 25964 18751 26016 18760
rect 25964 18717 25973 18751
rect 25973 18717 26007 18751
rect 26007 18717 26016 18751
rect 25964 18708 26016 18717
rect 27620 18708 27672 18760
rect 30932 18776 30984 18828
rect 27896 18708 27948 18760
rect 28724 18708 28776 18760
rect 29000 18708 29052 18760
rect 29368 18751 29420 18760
rect 29368 18717 29377 18751
rect 29377 18717 29411 18751
rect 29411 18717 29420 18751
rect 29368 18708 29420 18717
rect 28356 18683 28408 18692
rect 28356 18649 28365 18683
rect 28365 18649 28399 18683
rect 28399 18649 28408 18683
rect 28356 18640 28408 18649
rect 28632 18640 28684 18692
rect 29920 18708 29972 18760
rect 30288 18751 30340 18760
rect 30288 18717 30297 18751
rect 30297 18717 30331 18751
rect 30331 18717 30340 18751
rect 30288 18708 30340 18717
rect 34428 18776 34480 18828
rect 31208 18751 31260 18760
rect 31208 18717 31217 18751
rect 31217 18717 31251 18751
rect 31251 18717 31260 18751
rect 31208 18708 31260 18717
rect 31484 18708 31536 18760
rect 31760 18708 31812 18760
rect 34704 18708 34756 18760
rect 35348 18708 35400 18760
rect 30932 18640 30984 18692
rect 31852 18683 31904 18692
rect 25688 18572 25740 18624
rect 25964 18572 26016 18624
rect 27436 18572 27488 18624
rect 27988 18572 28040 18624
rect 28816 18572 28868 18624
rect 29276 18572 29328 18624
rect 29920 18572 29972 18624
rect 30196 18572 30248 18624
rect 31852 18649 31861 18683
rect 31861 18649 31895 18683
rect 31895 18649 31904 18683
rect 31852 18640 31904 18649
rect 32864 18640 32916 18692
rect 35808 18751 35860 18760
rect 35808 18717 35817 18751
rect 35817 18717 35851 18751
rect 35851 18717 35860 18751
rect 35808 18708 35860 18717
rect 35900 18751 35952 18760
rect 35900 18717 35909 18751
rect 35909 18717 35943 18751
rect 35943 18717 35952 18751
rect 35900 18708 35952 18717
rect 38936 18776 38988 18828
rect 39120 18708 39172 18760
rect 39212 18751 39264 18760
rect 39212 18717 39221 18751
rect 39221 18717 39255 18751
rect 39255 18717 39264 18751
rect 39212 18708 39264 18717
rect 32220 18572 32272 18624
rect 34612 18572 34664 18624
rect 36176 18615 36228 18624
rect 36176 18581 36185 18615
rect 36185 18581 36219 18615
rect 36219 18581 36228 18615
rect 36176 18572 36228 18581
rect 38568 18572 38620 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 1860 18368 1912 18420
rect 3332 18368 3384 18420
rect 3700 18368 3752 18420
rect 2504 18300 2556 18352
rect 4804 18368 4856 18420
rect 5448 18368 5500 18420
rect 8116 18368 8168 18420
rect 10048 18368 10100 18420
rect 11152 18368 11204 18420
rect 12716 18368 12768 18420
rect 14188 18368 14240 18420
rect 16028 18368 16080 18420
rect 16764 18411 16816 18420
rect 16764 18377 16773 18411
rect 16773 18377 16807 18411
rect 16807 18377 16816 18411
rect 16764 18368 16816 18377
rect 20260 18368 20312 18420
rect 4068 18343 4120 18352
rect 4068 18309 4077 18343
rect 4077 18309 4111 18343
rect 4111 18309 4120 18343
rect 4068 18300 4120 18309
rect 4160 18300 4212 18352
rect 5356 18300 5408 18352
rect 7840 18300 7892 18352
rect 12808 18300 12860 18352
rect 14096 18300 14148 18352
rect 16304 18300 16356 18352
rect 7748 18275 7800 18284
rect 7748 18241 7757 18275
rect 7757 18241 7791 18275
rect 7791 18241 7800 18275
rect 7748 18232 7800 18241
rect 15568 18275 15620 18284
rect 15568 18241 15577 18275
rect 15577 18241 15611 18275
rect 15611 18241 15620 18275
rect 15568 18232 15620 18241
rect 15936 18232 15988 18284
rect 21824 18232 21876 18284
rect 22284 18300 22336 18352
rect 22192 18275 22244 18284
rect 22192 18241 22201 18275
rect 22201 18241 22235 18275
rect 22235 18241 22244 18275
rect 22192 18232 22244 18241
rect 22376 18275 22428 18284
rect 22376 18241 22385 18275
rect 22385 18241 22419 18275
rect 22419 18241 22428 18275
rect 22376 18232 22428 18241
rect 4620 18164 4672 18216
rect 5540 18207 5592 18216
rect 5540 18173 5549 18207
rect 5549 18173 5583 18207
rect 5583 18173 5592 18207
rect 5540 18164 5592 18173
rect 7012 18207 7064 18216
rect 7012 18173 7021 18207
rect 7021 18173 7055 18207
rect 7055 18173 7064 18207
rect 7012 18164 7064 18173
rect 11060 18164 11112 18216
rect 12256 18207 12308 18216
rect 12256 18173 12265 18207
rect 12265 18173 12299 18207
rect 12299 18173 12308 18207
rect 12256 18164 12308 18173
rect 5448 18096 5500 18148
rect 7472 18096 7524 18148
rect 7564 18096 7616 18148
rect 12440 18096 12492 18148
rect 4436 18028 4488 18080
rect 4712 18028 4764 18080
rect 9220 18028 9272 18080
rect 12808 18207 12860 18216
rect 12808 18173 12817 18207
rect 12817 18173 12851 18207
rect 12851 18173 12860 18207
rect 12808 18164 12860 18173
rect 13268 18164 13320 18216
rect 18144 18164 18196 18216
rect 15476 18096 15528 18148
rect 16580 18096 16632 18148
rect 15752 18071 15804 18080
rect 15752 18037 15761 18071
rect 15761 18037 15795 18071
rect 15795 18037 15804 18071
rect 15752 18028 15804 18037
rect 18604 18028 18656 18080
rect 23940 18232 23992 18284
rect 24676 18275 24728 18284
rect 24676 18241 24685 18275
rect 24685 18241 24719 18275
rect 24719 18241 24728 18275
rect 24676 18232 24728 18241
rect 24124 18164 24176 18216
rect 24768 18164 24820 18216
rect 27160 18368 27212 18420
rect 27436 18368 27488 18420
rect 31576 18368 31628 18420
rect 25780 18300 25832 18352
rect 26056 18232 26108 18284
rect 28172 18300 28224 18352
rect 26516 18275 26568 18284
rect 26516 18241 26525 18275
rect 26525 18241 26559 18275
rect 26559 18241 26568 18275
rect 26516 18232 26568 18241
rect 27068 18232 27120 18284
rect 27712 18232 27764 18284
rect 27988 18232 28040 18284
rect 26240 18096 26292 18148
rect 26792 18164 26844 18216
rect 27252 18164 27304 18216
rect 31852 18300 31904 18352
rect 33600 18300 33652 18352
rect 34428 18300 34480 18352
rect 30012 18164 30064 18216
rect 32404 18232 32456 18284
rect 33784 18232 33836 18284
rect 35440 18232 35492 18284
rect 36452 18232 36504 18284
rect 38016 18232 38068 18284
rect 38292 18232 38344 18284
rect 38568 18275 38620 18284
rect 38568 18241 38577 18275
rect 38577 18241 38611 18275
rect 38611 18241 38620 18275
rect 38568 18232 38620 18241
rect 34520 18164 34572 18216
rect 36176 18164 36228 18216
rect 39396 18207 39448 18216
rect 39396 18173 39405 18207
rect 39405 18173 39439 18207
rect 39439 18173 39448 18207
rect 39396 18164 39448 18173
rect 39672 18207 39724 18216
rect 39672 18173 39681 18207
rect 39681 18173 39715 18207
rect 39715 18173 39724 18207
rect 39672 18164 39724 18173
rect 29368 18096 29420 18148
rect 33140 18096 33192 18148
rect 22376 18028 22428 18080
rect 23848 18028 23900 18080
rect 26424 18028 26476 18080
rect 26976 18071 27028 18080
rect 26976 18037 26985 18071
rect 26985 18037 27019 18071
rect 27019 18037 27028 18071
rect 26976 18028 27028 18037
rect 27620 18028 27672 18080
rect 27988 18028 28040 18080
rect 31484 18028 31536 18080
rect 32128 18028 32180 18080
rect 34060 18096 34112 18148
rect 37464 18096 37516 18148
rect 38568 18096 38620 18148
rect 38752 18028 38804 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 12808 17867 12860 17876
rect 12808 17833 12817 17867
rect 12817 17833 12851 17867
rect 12851 17833 12860 17867
rect 12808 17824 12860 17833
rect 13452 17824 13504 17876
rect 9588 17756 9640 17808
rect 16580 17867 16632 17876
rect 16580 17833 16589 17867
rect 16589 17833 16623 17867
rect 16623 17833 16632 17867
rect 16580 17824 16632 17833
rect 17040 17867 17092 17876
rect 17040 17833 17049 17867
rect 17049 17833 17083 17867
rect 17083 17833 17092 17867
rect 17040 17824 17092 17833
rect 18052 17824 18104 17876
rect 4620 17688 4672 17740
rect 5264 17731 5316 17740
rect 5264 17697 5273 17731
rect 5273 17697 5307 17731
rect 5307 17697 5316 17731
rect 5264 17688 5316 17697
rect 8024 17688 8076 17740
rect 7288 17620 7340 17672
rect 3148 17552 3200 17604
rect 2780 17484 2832 17536
rect 7472 17552 7524 17604
rect 8760 17663 8812 17672
rect 8760 17629 8769 17663
rect 8769 17629 8803 17663
rect 8803 17629 8812 17663
rect 8760 17620 8812 17629
rect 9220 17663 9272 17672
rect 9220 17629 9229 17663
rect 9229 17629 9263 17663
rect 9263 17629 9272 17663
rect 9220 17620 9272 17629
rect 9680 17663 9732 17672
rect 9680 17629 9689 17663
rect 9689 17629 9723 17663
rect 9723 17629 9732 17663
rect 9680 17620 9732 17629
rect 10876 17688 10928 17740
rect 12808 17688 12860 17740
rect 18972 17756 19024 17808
rect 19800 17756 19852 17808
rect 19340 17688 19392 17740
rect 23480 17824 23532 17876
rect 23756 17824 23808 17876
rect 26424 17824 26476 17876
rect 26608 17824 26660 17876
rect 22192 17756 22244 17808
rect 28540 17824 28592 17876
rect 28816 17824 28868 17876
rect 32772 17824 32824 17876
rect 9956 17620 10008 17672
rect 13268 17620 13320 17672
rect 12900 17552 12952 17604
rect 5356 17484 5408 17536
rect 7288 17484 7340 17536
rect 8668 17527 8720 17536
rect 8668 17493 8677 17527
rect 8677 17493 8711 17527
rect 8711 17493 8720 17527
rect 8668 17484 8720 17493
rect 8852 17484 8904 17536
rect 9404 17484 9456 17536
rect 10048 17484 10100 17536
rect 11152 17527 11204 17536
rect 11152 17493 11161 17527
rect 11161 17493 11195 17527
rect 11195 17493 11204 17527
rect 11152 17484 11204 17493
rect 14188 17484 14240 17536
rect 16948 17620 17000 17672
rect 18236 17663 18288 17672
rect 18236 17629 18245 17663
rect 18245 17629 18279 17663
rect 18279 17629 18288 17663
rect 18236 17620 18288 17629
rect 20812 17620 20864 17672
rect 21824 17620 21876 17672
rect 22376 17663 22428 17672
rect 22376 17629 22385 17663
rect 22385 17629 22419 17663
rect 22419 17629 22428 17663
rect 22376 17620 22428 17629
rect 22652 17663 22704 17672
rect 22652 17629 22661 17663
rect 22661 17629 22695 17663
rect 22695 17629 22704 17663
rect 22652 17620 22704 17629
rect 24308 17688 24360 17740
rect 30932 17756 30984 17808
rect 31300 17756 31352 17808
rect 34060 17867 34112 17876
rect 34060 17833 34069 17867
rect 34069 17833 34103 17867
rect 34103 17833 34112 17867
rect 34060 17824 34112 17833
rect 39856 17824 39908 17876
rect 33508 17756 33560 17808
rect 23388 17620 23440 17672
rect 23756 17620 23808 17672
rect 24216 17620 24268 17672
rect 26884 17620 26936 17672
rect 28540 17663 28592 17672
rect 28540 17629 28549 17663
rect 28549 17629 28583 17663
rect 28583 17629 28592 17663
rect 28540 17620 28592 17629
rect 28724 17620 28776 17672
rect 28816 17663 28868 17672
rect 28816 17629 28825 17663
rect 28825 17629 28859 17663
rect 28859 17629 28868 17663
rect 28816 17620 28868 17629
rect 29276 17620 29328 17672
rect 31024 17620 31076 17672
rect 31484 17663 31536 17672
rect 31484 17629 31493 17663
rect 31493 17629 31527 17663
rect 31527 17629 31536 17663
rect 31484 17620 31536 17629
rect 17040 17595 17092 17604
rect 17040 17561 17049 17595
rect 17049 17561 17083 17595
rect 17083 17561 17092 17595
rect 17040 17552 17092 17561
rect 18604 17552 18656 17604
rect 19248 17552 19300 17604
rect 18052 17527 18104 17536
rect 18052 17493 18061 17527
rect 18061 17493 18095 17527
rect 18095 17493 18104 17527
rect 18052 17484 18104 17493
rect 18420 17484 18472 17536
rect 19156 17484 19208 17536
rect 23664 17552 23716 17604
rect 24400 17552 24452 17604
rect 27712 17552 27764 17604
rect 28448 17552 28500 17604
rect 29092 17552 29144 17604
rect 31300 17595 31352 17604
rect 31300 17561 31309 17595
rect 31309 17561 31343 17595
rect 31343 17561 31352 17595
rect 31300 17552 31352 17561
rect 31852 17663 31904 17672
rect 31852 17629 31861 17663
rect 31861 17629 31895 17663
rect 31895 17629 31904 17663
rect 31852 17620 31904 17629
rect 32128 17620 32180 17672
rect 32680 17620 32732 17672
rect 33048 17688 33100 17740
rect 36544 17756 36596 17808
rect 38292 17756 38344 17808
rect 32956 17663 33008 17672
rect 32956 17629 32965 17663
rect 32965 17629 32999 17663
rect 32999 17629 33008 17663
rect 32956 17620 33008 17629
rect 33324 17663 33376 17672
rect 33324 17629 33333 17663
rect 33333 17629 33367 17663
rect 33367 17629 33376 17663
rect 33324 17620 33376 17629
rect 33784 17620 33836 17672
rect 34152 17663 34204 17672
rect 34152 17629 34161 17663
rect 34161 17629 34195 17663
rect 34195 17629 34204 17663
rect 34152 17620 34204 17629
rect 34428 17620 34480 17672
rect 23480 17484 23532 17536
rect 24216 17484 24268 17536
rect 27160 17484 27212 17536
rect 27252 17484 27304 17536
rect 33508 17595 33560 17604
rect 33508 17561 33517 17595
rect 33517 17561 33551 17595
rect 33551 17561 33560 17595
rect 33508 17552 33560 17561
rect 33600 17595 33652 17604
rect 33600 17561 33609 17595
rect 33609 17561 33643 17595
rect 33643 17561 33652 17595
rect 33600 17552 33652 17561
rect 36084 17663 36136 17672
rect 36084 17629 36093 17663
rect 36093 17629 36127 17663
rect 36127 17629 36136 17663
rect 36084 17620 36136 17629
rect 36176 17663 36228 17672
rect 36176 17629 36186 17663
rect 36186 17629 36220 17663
rect 36220 17629 36228 17663
rect 37096 17688 37148 17740
rect 38568 17731 38620 17740
rect 38568 17697 38577 17731
rect 38577 17697 38611 17731
rect 38611 17697 38620 17731
rect 38568 17688 38620 17697
rect 36176 17620 36228 17629
rect 36544 17663 36596 17672
rect 36544 17629 36558 17663
rect 36558 17629 36592 17663
rect 36592 17629 36596 17663
rect 36544 17620 36596 17629
rect 32956 17484 33008 17536
rect 34152 17484 34204 17536
rect 34428 17527 34480 17536
rect 34428 17493 34437 17527
rect 34437 17493 34471 17527
rect 34471 17493 34480 17527
rect 34428 17484 34480 17493
rect 34888 17484 34940 17536
rect 38476 17620 38528 17672
rect 37372 17552 37424 17604
rect 38108 17484 38160 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 5264 17280 5316 17332
rect 5356 17280 5408 17332
rect 2780 17255 2832 17264
rect 2780 17221 2789 17255
rect 2789 17221 2823 17255
rect 2823 17221 2832 17255
rect 2780 17212 2832 17221
rect 3792 17212 3844 17264
rect 6552 17212 6604 17264
rect 7380 17212 7432 17264
rect 2504 17187 2556 17196
rect 2504 17153 2513 17187
rect 2513 17153 2547 17187
rect 2547 17153 2556 17187
rect 2504 17144 2556 17153
rect 6920 17144 6972 17196
rect 7472 17144 7524 17196
rect 7840 17212 7892 17264
rect 8024 17144 8076 17196
rect 11244 17280 11296 17332
rect 17408 17280 17460 17332
rect 18420 17323 18472 17332
rect 18420 17289 18429 17323
rect 18429 17289 18463 17323
rect 18463 17289 18472 17323
rect 18420 17280 18472 17289
rect 18512 17280 18564 17332
rect 20628 17280 20680 17332
rect 24400 17323 24452 17332
rect 24400 17289 24409 17323
rect 24409 17289 24443 17323
rect 24443 17289 24452 17323
rect 24400 17280 24452 17289
rect 9404 17212 9456 17264
rect 8668 17144 8720 17196
rect 11060 17212 11112 17264
rect 14648 17212 14700 17264
rect 5448 17076 5500 17128
rect 6000 17076 6052 17128
rect 7656 17076 7708 17128
rect 12532 17144 12584 17196
rect 10876 17008 10928 17060
rect 11888 17076 11940 17128
rect 16856 17144 16908 17196
rect 17776 17212 17828 17264
rect 18604 17255 18656 17264
rect 18604 17221 18613 17255
rect 18613 17221 18647 17255
rect 18647 17221 18656 17255
rect 18604 17212 18656 17221
rect 18696 17212 18748 17264
rect 19248 17255 19300 17264
rect 19248 17221 19257 17255
rect 19257 17221 19291 17255
rect 19291 17221 19300 17255
rect 19248 17212 19300 17221
rect 19616 17255 19668 17264
rect 19616 17221 19625 17255
rect 19625 17221 19659 17255
rect 19659 17221 19668 17255
rect 19616 17212 19668 17221
rect 17040 17187 17092 17196
rect 17040 17153 17049 17187
rect 17049 17153 17083 17187
rect 17083 17153 17092 17187
rect 17040 17144 17092 17153
rect 18236 17144 18288 17196
rect 19432 17187 19484 17196
rect 19432 17153 19441 17187
rect 19441 17153 19475 17187
rect 19475 17153 19484 17187
rect 19432 17144 19484 17153
rect 19800 17187 19852 17196
rect 19800 17153 19809 17187
rect 19809 17153 19843 17187
rect 19843 17153 19852 17187
rect 19800 17144 19852 17153
rect 7380 16983 7432 16992
rect 7380 16949 7389 16983
rect 7389 16949 7423 16983
rect 7423 16949 7432 16983
rect 7380 16940 7432 16949
rect 7564 16940 7616 16992
rect 8116 16940 8168 16992
rect 9588 16940 9640 16992
rect 11980 16940 12032 16992
rect 13636 16983 13688 16992
rect 13636 16949 13645 16983
rect 13645 16949 13679 16983
rect 13679 16949 13688 16983
rect 13636 16940 13688 16949
rect 16948 16940 17000 16992
rect 20168 17076 20220 17128
rect 22928 17076 22980 17128
rect 23296 17076 23348 17128
rect 24216 17187 24268 17196
rect 24216 17153 24225 17187
rect 24225 17153 24259 17187
rect 24259 17153 24268 17187
rect 24216 17144 24268 17153
rect 27252 17280 27304 17332
rect 27344 17280 27396 17332
rect 25136 17212 25188 17264
rect 28816 17280 28868 17332
rect 33508 17280 33560 17332
rect 38384 17323 38436 17332
rect 38384 17289 38393 17323
rect 38393 17289 38427 17323
rect 38427 17289 38436 17323
rect 38384 17280 38436 17289
rect 24676 17187 24728 17196
rect 24676 17153 24685 17187
rect 24685 17153 24719 17187
rect 24719 17153 24728 17187
rect 24676 17144 24728 17153
rect 25596 17144 25648 17196
rect 20628 17008 20680 17060
rect 25044 17076 25096 17128
rect 27160 17187 27212 17196
rect 27160 17153 27169 17187
rect 27169 17153 27203 17187
rect 27203 17153 27212 17187
rect 27160 17144 27212 17153
rect 28172 17144 28224 17196
rect 32680 17212 32732 17264
rect 19156 16940 19208 16992
rect 19984 16983 20036 16992
rect 19984 16949 19993 16983
rect 19993 16949 20027 16983
rect 20027 16949 20036 16983
rect 19984 16940 20036 16949
rect 22836 16940 22888 16992
rect 24860 16983 24912 16992
rect 24860 16949 24869 16983
rect 24869 16949 24903 16983
rect 24903 16949 24912 16983
rect 25228 17008 25280 17060
rect 27804 17008 27856 17060
rect 28724 17076 28776 17128
rect 29000 17008 29052 17060
rect 31944 17144 31996 17196
rect 32588 17144 32640 17196
rect 33600 17144 33652 17196
rect 34428 17212 34480 17264
rect 30380 17119 30432 17128
rect 30380 17085 30389 17119
rect 30389 17085 30423 17119
rect 30423 17085 30432 17119
rect 30380 17076 30432 17085
rect 34796 17144 34848 17196
rect 35256 17187 35308 17196
rect 35256 17153 35263 17187
rect 35263 17153 35308 17187
rect 35256 17144 35308 17153
rect 35348 17187 35400 17196
rect 35348 17153 35357 17187
rect 35357 17153 35391 17187
rect 35391 17153 35400 17187
rect 35348 17144 35400 17153
rect 33600 17008 33652 17060
rect 35348 17008 35400 17060
rect 35992 17144 36044 17196
rect 38108 17187 38160 17196
rect 38108 17153 38117 17187
rect 38117 17153 38151 17187
rect 38151 17153 38160 17187
rect 38108 17144 38160 17153
rect 36452 17076 36504 17128
rect 37096 17076 37148 17128
rect 24860 16940 24912 16949
rect 28356 16940 28408 16992
rect 29276 16940 29328 16992
rect 35440 16940 35492 16992
rect 37924 16983 37976 16992
rect 37924 16949 37933 16983
rect 37933 16949 37967 16983
rect 37967 16949 37976 16983
rect 37924 16940 37976 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 6552 16779 6604 16788
rect 6552 16745 6561 16779
rect 6561 16745 6595 16779
rect 6595 16745 6604 16779
rect 6552 16736 6604 16745
rect 6920 16736 6972 16788
rect 7288 16779 7340 16788
rect 7288 16745 7297 16779
rect 7297 16745 7331 16779
rect 7331 16745 7340 16779
rect 7288 16736 7340 16745
rect 7656 16736 7708 16788
rect 7012 16711 7064 16720
rect 7012 16677 7021 16711
rect 7021 16677 7055 16711
rect 7055 16677 7064 16711
rect 7012 16668 7064 16677
rect 4804 16643 4856 16652
rect 4804 16609 4813 16643
rect 4813 16609 4847 16643
rect 4847 16609 4856 16643
rect 4804 16600 4856 16609
rect 6092 16600 6144 16652
rect 6828 16600 6880 16652
rect 7564 16600 7616 16652
rect 8208 16779 8260 16788
rect 8208 16745 8217 16779
rect 8217 16745 8251 16779
rect 8251 16745 8260 16779
rect 8208 16736 8260 16745
rect 12348 16736 12400 16788
rect 16396 16736 16448 16788
rect 19064 16736 19116 16788
rect 7932 16668 7984 16720
rect 7288 16532 7340 16584
rect 8116 16643 8168 16652
rect 8116 16609 8125 16643
rect 8125 16609 8159 16643
rect 8159 16609 8168 16643
rect 8116 16600 8168 16609
rect 9496 16643 9548 16652
rect 9496 16609 9505 16643
rect 9505 16609 9539 16643
rect 9539 16609 9548 16643
rect 9496 16600 9548 16609
rect 10508 16643 10560 16652
rect 10508 16609 10517 16643
rect 10517 16609 10551 16643
rect 10551 16609 10560 16643
rect 10508 16600 10560 16609
rect 12164 16668 12216 16720
rect 11704 16643 11756 16652
rect 11704 16609 11713 16643
rect 11713 16609 11747 16643
rect 11747 16609 11756 16643
rect 11704 16600 11756 16609
rect 3792 16464 3844 16516
rect 6920 16464 6972 16516
rect 7380 16464 7432 16516
rect 11244 16532 11296 16584
rect 12992 16600 13044 16652
rect 8208 16464 8260 16516
rect 7288 16439 7340 16448
rect 7288 16405 7315 16439
rect 7315 16405 7340 16439
rect 7288 16396 7340 16405
rect 7656 16439 7708 16448
rect 7656 16405 7665 16439
rect 7665 16405 7699 16439
rect 7699 16405 7708 16439
rect 7656 16396 7708 16405
rect 8392 16439 8444 16448
rect 8392 16405 8401 16439
rect 8401 16405 8435 16439
rect 8435 16405 8444 16439
rect 8392 16396 8444 16405
rect 8944 16439 8996 16448
rect 8944 16405 8953 16439
rect 8953 16405 8987 16439
rect 8987 16405 8996 16439
rect 8944 16396 8996 16405
rect 11060 16507 11112 16516
rect 11060 16473 11069 16507
rect 11069 16473 11103 16507
rect 11103 16473 11112 16507
rect 11060 16464 11112 16473
rect 12164 16464 12216 16516
rect 10692 16439 10744 16448
rect 10692 16405 10701 16439
rect 10701 16405 10735 16439
rect 10735 16405 10744 16439
rect 10692 16396 10744 16405
rect 11704 16396 11756 16448
rect 12532 16439 12584 16448
rect 12532 16405 12541 16439
rect 12541 16405 12575 16439
rect 12575 16405 12584 16439
rect 12532 16396 12584 16405
rect 13820 16600 13872 16652
rect 14004 16600 14056 16652
rect 14372 16643 14424 16652
rect 14372 16609 14381 16643
rect 14381 16609 14415 16643
rect 14415 16609 14424 16643
rect 14372 16600 14424 16609
rect 14096 16575 14148 16584
rect 14096 16541 14105 16575
rect 14105 16541 14139 16575
rect 14139 16541 14148 16575
rect 14096 16532 14148 16541
rect 14464 16532 14516 16584
rect 14556 16575 14608 16584
rect 14556 16541 14565 16575
rect 14565 16541 14599 16575
rect 14599 16541 14608 16575
rect 14556 16532 14608 16541
rect 15016 16643 15068 16652
rect 15016 16609 15025 16643
rect 15025 16609 15059 16643
rect 15059 16609 15068 16643
rect 15016 16600 15068 16609
rect 17408 16668 17460 16720
rect 18052 16668 18104 16720
rect 22652 16668 22704 16720
rect 19432 16600 19484 16652
rect 19800 16600 19852 16652
rect 20444 16600 20496 16652
rect 20628 16600 20680 16652
rect 22192 16600 22244 16652
rect 13728 16396 13780 16448
rect 13820 16396 13872 16448
rect 14188 16439 14240 16448
rect 14188 16405 14197 16439
rect 14197 16405 14231 16439
rect 14231 16405 14240 16439
rect 14188 16396 14240 16405
rect 16672 16396 16724 16448
rect 17224 16532 17276 16584
rect 18144 16532 18196 16584
rect 21180 16532 21232 16584
rect 20720 16507 20772 16516
rect 20720 16473 20737 16507
rect 20737 16473 20772 16507
rect 20720 16464 20772 16473
rect 20812 16507 20864 16516
rect 20812 16473 20821 16507
rect 20821 16473 20855 16507
rect 20855 16473 20864 16507
rect 20812 16464 20864 16473
rect 20904 16507 20956 16516
rect 20904 16473 20913 16507
rect 20913 16473 20947 16507
rect 20947 16473 20956 16507
rect 20904 16464 20956 16473
rect 19616 16396 19668 16448
rect 19984 16396 20036 16448
rect 21824 16532 21876 16584
rect 22284 16507 22336 16516
rect 22284 16473 22293 16507
rect 22293 16473 22327 16507
rect 22327 16473 22336 16507
rect 22284 16464 22336 16473
rect 22652 16532 22704 16584
rect 22928 16779 22980 16788
rect 22928 16745 22937 16779
rect 22937 16745 22971 16779
rect 22971 16745 22980 16779
rect 22928 16736 22980 16745
rect 26700 16736 26752 16788
rect 28080 16736 28132 16788
rect 28264 16736 28316 16788
rect 28632 16668 28684 16720
rect 29092 16736 29144 16788
rect 35348 16736 35400 16788
rect 36452 16736 36504 16788
rect 36820 16736 36872 16788
rect 38292 16736 38344 16788
rect 22928 16643 22980 16652
rect 22928 16609 22937 16643
rect 22937 16609 22971 16643
rect 22971 16609 22980 16643
rect 22928 16600 22980 16609
rect 25688 16643 25740 16652
rect 25688 16609 25697 16643
rect 25697 16609 25731 16643
rect 25731 16609 25740 16643
rect 25688 16600 25740 16609
rect 25780 16600 25832 16652
rect 28172 16600 28224 16652
rect 32956 16668 33008 16720
rect 36912 16668 36964 16720
rect 37372 16668 37424 16720
rect 24492 16532 24544 16584
rect 24768 16507 24820 16516
rect 24768 16473 24777 16507
rect 24777 16473 24811 16507
rect 24811 16473 24820 16507
rect 24768 16464 24820 16473
rect 25504 16575 25556 16584
rect 25504 16541 25513 16575
rect 25513 16541 25547 16575
rect 25547 16541 25556 16575
rect 25504 16532 25556 16541
rect 26056 16575 26108 16584
rect 26056 16541 26065 16575
rect 26065 16541 26099 16575
rect 26099 16541 26108 16575
rect 26056 16532 26108 16541
rect 25596 16464 25648 16516
rect 26424 16575 26476 16584
rect 26424 16541 26433 16575
rect 26433 16541 26467 16575
rect 26467 16541 26476 16575
rect 26424 16532 26476 16541
rect 28080 16532 28132 16584
rect 28632 16575 28684 16584
rect 28632 16541 28677 16575
rect 28677 16541 28684 16575
rect 28632 16532 28684 16541
rect 31392 16532 31444 16584
rect 27988 16464 28040 16516
rect 28448 16507 28500 16516
rect 28448 16473 28457 16507
rect 28457 16473 28491 16507
rect 28491 16473 28500 16507
rect 28448 16464 28500 16473
rect 30012 16464 30064 16516
rect 22560 16396 22612 16448
rect 23388 16396 23440 16448
rect 24492 16396 24544 16448
rect 27436 16396 27488 16448
rect 33600 16464 33652 16516
rect 34060 16464 34112 16516
rect 30748 16396 30800 16448
rect 31944 16396 31996 16448
rect 34980 16396 35032 16448
rect 36360 16532 36412 16584
rect 36636 16575 36688 16584
rect 36636 16541 36643 16575
rect 36643 16541 36688 16575
rect 36636 16532 36688 16541
rect 36820 16600 36872 16652
rect 38476 16643 38528 16652
rect 38476 16609 38485 16643
rect 38485 16609 38519 16643
rect 38519 16609 38528 16643
rect 38476 16600 38528 16609
rect 37464 16532 37516 16584
rect 38016 16532 38068 16584
rect 37004 16396 37056 16448
rect 39488 16396 39540 16448
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 7104 16192 7156 16244
rect 7288 16192 7340 16244
rect 8208 16192 8260 16244
rect 9496 16235 9548 16244
rect 9496 16201 9505 16235
rect 9505 16201 9539 16235
rect 9539 16201 9548 16235
rect 9496 16192 9548 16201
rect 3240 16124 3292 16176
rect 3792 16124 3844 16176
rect 5448 16056 5500 16108
rect 5816 15988 5868 16040
rect 10692 16124 10744 16176
rect 9404 16099 9456 16108
rect 9404 16065 9413 16099
rect 9413 16065 9447 16099
rect 9447 16065 9456 16099
rect 9404 16056 9456 16065
rect 11060 16192 11112 16244
rect 11704 16192 11756 16244
rect 12256 16192 12308 16244
rect 24768 16192 24820 16244
rect 25872 16192 25924 16244
rect 26332 16192 26384 16244
rect 26424 16192 26476 16244
rect 11244 16124 11296 16176
rect 12992 16124 13044 16176
rect 14096 16124 14148 16176
rect 11980 16099 12032 16108
rect 11980 16065 11989 16099
rect 11989 16065 12023 16099
rect 12023 16065 12032 16099
rect 11980 16056 12032 16065
rect 12808 16056 12860 16108
rect 13636 16099 13688 16108
rect 13636 16065 13645 16099
rect 13645 16065 13679 16099
rect 13679 16065 13688 16099
rect 13636 16056 13688 16065
rect 13820 16056 13872 16108
rect 14464 16124 14516 16176
rect 14556 16124 14608 16176
rect 15108 16056 15160 16108
rect 16488 16124 16540 16176
rect 22284 16124 22336 16176
rect 16120 16099 16172 16108
rect 16120 16065 16129 16099
rect 16129 16065 16163 16099
rect 16163 16065 16172 16099
rect 16120 16056 16172 16065
rect 10876 15920 10928 15972
rect 14372 15988 14424 16040
rect 16396 16099 16448 16108
rect 16396 16065 16405 16099
rect 16405 16065 16439 16099
rect 16439 16065 16448 16099
rect 16396 16056 16448 16065
rect 25688 16124 25740 16176
rect 24492 16099 24544 16108
rect 24492 16065 24501 16099
rect 24501 16065 24535 16099
rect 24535 16065 24544 16099
rect 24492 16056 24544 16065
rect 24676 16056 24728 16108
rect 25228 16056 25280 16108
rect 28080 16192 28132 16244
rect 29552 16192 29604 16244
rect 30012 16235 30064 16244
rect 30012 16201 30021 16235
rect 30021 16201 30055 16235
rect 30055 16201 30064 16235
rect 30012 16192 30064 16201
rect 27528 16124 27580 16176
rect 27436 16099 27488 16108
rect 27436 16065 27445 16099
rect 27445 16065 27479 16099
rect 27479 16065 27488 16099
rect 27436 16056 27488 16065
rect 27712 16056 27764 16108
rect 27988 16056 28040 16108
rect 28264 16056 28316 16108
rect 28356 16099 28408 16108
rect 28356 16065 28365 16099
rect 28365 16065 28399 16099
rect 28399 16065 28408 16099
rect 28356 16056 28408 16065
rect 30472 16192 30524 16244
rect 30380 16167 30432 16176
rect 30380 16133 30389 16167
rect 30389 16133 30423 16167
rect 30423 16133 30432 16167
rect 30380 16124 30432 16133
rect 31300 16167 31352 16176
rect 31300 16133 31309 16167
rect 31309 16133 31343 16167
rect 31343 16133 31352 16167
rect 31300 16124 31352 16133
rect 33324 16124 33376 16176
rect 34060 16124 34112 16176
rect 34244 16124 34296 16176
rect 34428 16167 34480 16176
rect 34428 16133 34437 16167
rect 34437 16133 34471 16167
rect 34471 16133 34480 16167
rect 34428 16124 34480 16133
rect 17408 15988 17460 16040
rect 29276 15988 29328 16040
rect 12164 15920 12216 15972
rect 11428 15852 11480 15904
rect 11796 15852 11848 15904
rect 13268 15852 13320 15904
rect 15844 15920 15896 15972
rect 16120 15920 16172 15972
rect 20720 15920 20772 15972
rect 27252 15920 27304 15972
rect 28448 15920 28500 15972
rect 30564 16099 30616 16108
rect 30564 16065 30573 16099
rect 30573 16065 30607 16099
rect 30607 16065 30616 16099
rect 30564 16056 30616 16065
rect 30748 16056 30800 16108
rect 31392 16099 31444 16108
rect 31392 16065 31401 16099
rect 31401 16065 31435 16099
rect 31435 16065 31444 16099
rect 31392 16056 31444 16065
rect 31484 16099 31536 16108
rect 31484 16065 31493 16099
rect 31493 16065 31527 16099
rect 31527 16065 31536 16099
rect 31484 16056 31536 16065
rect 33232 16056 33284 16108
rect 33876 16056 33928 16108
rect 34520 16099 34572 16108
rect 34520 16065 34529 16099
rect 34529 16065 34563 16099
rect 34563 16065 34572 16099
rect 34520 16056 34572 16065
rect 35164 16167 35216 16176
rect 35164 16133 35173 16167
rect 35173 16133 35207 16167
rect 35207 16133 35216 16167
rect 35164 16124 35216 16133
rect 36820 16167 36872 16176
rect 36820 16133 36829 16167
rect 36829 16133 36863 16167
rect 36863 16133 36872 16167
rect 36820 16124 36872 16133
rect 34888 16099 34940 16108
rect 34888 16065 34897 16099
rect 34897 16065 34931 16099
rect 34931 16065 34940 16099
rect 34888 16056 34940 16065
rect 36544 16099 36596 16108
rect 36544 16065 36553 16099
rect 36553 16065 36587 16099
rect 36587 16065 36596 16099
rect 36544 16056 36596 16065
rect 31024 16031 31076 16040
rect 31024 15997 31033 16031
rect 31033 15997 31067 16031
rect 31067 15997 31076 16031
rect 31024 15988 31076 15997
rect 31576 15988 31628 16040
rect 34244 15988 34296 16040
rect 34796 16031 34848 16040
rect 34796 15997 34805 16031
rect 34805 15997 34839 16031
rect 34839 15997 34848 16031
rect 34796 15988 34848 15997
rect 34980 15988 35032 16040
rect 37464 16056 37516 16108
rect 31300 15920 31352 15972
rect 38292 15920 38344 15972
rect 14188 15852 14240 15904
rect 18420 15852 18472 15904
rect 27528 15852 27580 15904
rect 27896 15895 27948 15904
rect 27896 15861 27905 15895
rect 27905 15861 27939 15895
rect 27939 15861 27948 15895
rect 27896 15852 27948 15861
rect 27988 15895 28040 15904
rect 27988 15861 27997 15895
rect 27997 15861 28031 15895
rect 28031 15861 28040 15895
rect 27988 15852 28040 15861
rect 28080 15852 28132 15904
rect 28356 15852 28408 15904
rect 28908 15852 28960 15904
rect 30288 15852 30340 15904
rect 30840 15852 30892 15904
rect 32772 15852 32824 15904
rect 33784 15852 33836 15904
rect 34888 15852 34940 15904
rect 37096 15895 37148 15904
rect 37096 15861 37105 15895
rect 37105 15861 37139 15895
rect 37139 15861 37148 15895
rect 37096 15852 37148 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 5448 15691 5500 15700
rect 5448 15657 5457 15691
rect 5457 15657 5491 15691
rect 5491 15657 5500 15691
rect 5448 15648 5500 15657
rect 6092 15648 6144 15700
rect 9864 15648 9916 15700
rect 6000 15580 6052 15632
rect 5264 15512 5316 15564
rect 5540 15487 5592 15496
rect 5540 15453 5549 15487
rect 5549 15453 5583 15487
rect 5583 15453 5592 15487
rect 5540 15444 5592 15453
rect 5816 15512 5868 15564
rect 5908 15512 5960 15564
rect 6184 15444 6236 15496
rect 6552 15444 6604 15496
rect 6828 15487 6880 15496
rect 6828 15453 6837 15487
rect 6837 15453 6871 15487
rect 6871 15453 6880 15487
rect 6828 15444 6880 15453
rect 7012 15487 7064 15496
rect 7012 15453 7021 15487
rect 7021 15453 7055 15487
rect 7055 15453 7064 15487
rect 7012 15444 7064 15453
rect 8024 15487 8076 15496
rect 8024 15453 8033 15487
rect 8033 15453 8067 15487
rect 8067 15453 8076 15487
rect 8024 15444 8076 15453
rect 10048 15487 10100 15496
rect 10048 15453 10057 15487
rect 10057 15453 10091 15487
rect 10091 15453 10100 15487
rect 10048 15444 10100 15453
rect 16396 15691 16448 15700
rect 16396 15657 16405 15691
rect 16405 15657 16439 15691
rect 16439 15657 16448 15691
rect 16396 15648 16448 15657
rect 16764 15648 16816 15700
rect 17040 15691 17092 15700
rect 17040 15657 17049 15691
rect 17049 15657 17083 15691
rect 17083 15657 17092 15691
rect 17040 15648 17092 15657
rect 17408 15691 17460 15700
rect 17408 15657 17417 15691
rect 17417 15657 17451 15691
rect 17451 15657 17460 15691
rect 17408 15648 17460 15657
rect 19432 15648 19484 15700
rect 21548 15648 21600 15700
rect 22008 15691 22060 15700
rect 22008 15657 22017 15691
rect 22017 15657 22051 15691
rect 22051 15657 22060 15691
rect 22008 15648 22060 15657
rect 22192 15648 22244 15700
rect 24676 15648 24728 15700
rect 27252 15648 27304 15700
rect 28724 15648 28776 15700
rect 31852 15648 31904 15700
rect 33048 15691 33100 15700
rect 33048 15657 33057 15691
rect 33057 15657 33091 15691
rect 33091 15657 33100 15691
rect 33048 15648 33100 15657
rect 34336 15648 34388 15700
rect 34704 15648 34756 15700
rect 34980 15691 35032 15700
rect 34980 15657 34989 15691
rect 34989 15657 35023 15691
rect 35023 15657 35032 15691
rect 34980 15648 35032 15657
rect 37924 15648 37976 15700
rect 38292 15691 38344 15700
rect 38292 15657 38301 15691
rect 38301 15657 38335 15691
rect 38335 15657 38344 15691
rect 38292 15648 38344 15657
rect 17592 15512 17644 15564
rect 18512 15512 18564 15564
rect 19340 15580 19392 15632
rect 22008 15512 22060 15564
rect 22100 15512 22152 15564
rect 22836 15512 22888 15564
rect 30012 15580 30064 15632
rect 11060 15444 11112 15496
rect 5816 15419 5868 15428
rect 5816 15385 5825 15419
rect 5825 15385 5859 15419
rect 5859 15385 5868 15419
rect 5816 15376 5868 15385
rect 10508 15376 10560 15428
rect 11796 15487 11848 15496
rect 11796 15453 11805 15487
rect 11805 15453 11839 15487
rect 11839 15453 11848 15487
rect 11796 15444 11848 15453
rect 11888 15444 11940 15496
rect 12532 15444 12584 15496
rect 13176 15487 13228 15496
rect 13176 15453 13185 15487
rect 13185 15453 13219 15487
rect 13219 15453 13228 15487
rect 13176 15444 13228 15453
rect 12164 15376 12216 15428
rect 16672 15487 16724 15496
rect 16672 15453 16681 15487
rect 16681 15453 16715 15487
rect 16715 15453 16724 15487
rect 16672 15444 16724 15453
rect 16764 15444 16816 15496
rect 16948 15487 17000 15496
rect 16948 15453 16957 15487
rect 16957 15453 16991 15487
rect 16991 15453 17000 15487
rect 16948 15444 17000 15453
rect 17960 15444 18012 15496
rect 18052 15444 18104 15496
rect 18236 15444 18288 15496
rect 18420 15487 18472 15496
rect 18420 15453 18429 15487
rect 18429 15453 18463 15487
rect 18463 15453 18472 15487
rect 18420 15444 18472 15453
rect 20536 15444 20588 15496
rect 17776 15376 17828 15428
rect 22192 15487 22244 15496
rect 22192 15453 22201 15487
rect 22201 15453 22235 15487
rect 22235 15453 22244 15487
rect 22192 15444 22244 15453
rect 22468 15487 22520 15496
rect 22468 15453 22477 15487
rect 22477 15453 22511 15487
rect 22511 15453 22520 15487
rect 22468 15444 22520 15453
rect 23664 15444 23716 15496
rect 24400 15487 24452 15496
rect 24400 15453 24409 15487
rect 24409 15453 24443 15487
rect 24443 15453 24452 15487
rect 24400 15444 24452 15453
rect 24676 15444 24728 15496
rect 29920 15555 29972 15564
rect 25596 15444 25648 15496
rect 26240 15444 26292 15496
rect 28908 15487 28960 15496
rect 28908 15453 28917 15487
rect 28917 15453 28951 15487
rect 28951 15453 28960 15487
rect 28908 15444 28960 15453
rect 29092 15444 29144 15496
rect 29920 15521 29929 15555
rect 29929 15521 29963 15555
rect 29963 15521 29972 15555
rect 29920 15512 29972 15521
rect 24032 15419 24084 15428
rect 24032 15385 24041 15419
rect 24041 15385 24075 15419
rect 24075 15385 24084 15419
rect 24032 15376 24084 15385
rect 24124 15376 24176 15428
rect 26424 15376 26476 15428
rect 29828 15487 29880 15496
rect 29828 15453 29837 15487
rect 29837 15453 29871 15487
rect 29871 15453 29880 15487
rect 29828 15444 29880 15453
rect 29644 15376 29696 15428
rect 30196 15444 30248 15496
rect 30840 15487 30892 15496
rect 30840 15453 30849 15487
rect 30849 15453 30883 15487
rect 30883 15453 30892 15487
rect 30840 15444 30892 15453
rect 31024 15487 31076 15496
rect 31024 15453 31033 15487
rect 31033 15453 31067 15487
rect 31067 15453 31076 15487
rect 31024 15444 31076 15453
rect 31208 15487 31260 15496
rect 31208 15453 31217 15487
rect 31217 15453 31251 15487
rect 31251 15453 31260 15487
rect 31208 15444 31260 15453
rect 30748 15376 30800 15428
rect 31576 15487 31628 15496
rect 31576 15453 31586 15487
rect 31586 15453 31620 15487
rect 31620 15453 31628 15487
rect 31576 15444 31628 15453
rect 32496 15580 32548 15632
rect 32772 15512 32824 15564
rect 36544 15580 36596 15632
rect 36636 15580 36688 15632
rect 39212 15623 39264 15632
rect 39212 15589 39221 15623
rect 39221 15589 39255 15623
rect 39255 15589 39264 15623
rect 39212 15580 39264 15589
rect 34520 15512 34572 15564
rect 4620 15308 4672 15360
rect 6276 15308 6328 15360
rect 6552 15308 6604 15360
rect 7932 15351 7984 15360
rect 7932 15317 7941 15351
rect 7941 15317 7975 15351
rect 7975 15317 7984 15351
rect 7932 15308 7984 15317
rect 10048 15308 10100 15360
rect 10416 15351 10468 15360
rect 10416 15317 10425 15351
rect 10425 15317 10459 15351
rect 10459 15317 10468 15351
rect 10416 15308 10468 15317
rect 13360 15351 13412 15360
rect 13360 15317 13369 15351
rect 13369 15317 13403 15351
rect 13403 15317 13412 15351
rect 13360 15308 13412 15317
rect 17960 15351 18012 15360
rect 17960 15317 17969 15351
rect 17969 15317 18003 15351
rect 18003 15317 18012 15351
rect 17960 15308 18012 15317
rect 20536 15351 20588 15360
rect 20536 15317 20545 15351
rect 20545 15317 20579 15351
rect 20579 15317 20588 15351
rect 20536 15308 20588 15317
rect 21732 15308 21784 15360
rect 22652 15308 22704 15360
rect 28908 15308 28960 15360
rect 29276 15308 29328 15360
rect 30196 15308 30248 15360
rect 30288 15351 30340 15360
rect 30288 15317 30297 15351
rect 30297 15317 30331 15351
rect 30331 15317 30340 15351
rect 30288 15308 30340 15317
rect 30380 15308 30432 15360
rect 31760 15419 31812 15428
rect 31760 15385 31769 15419
rect 31769 15385 31803 15419
rect 31803 15385 31812 15419
rect 31760 15376 31812 15385
rect 31852 15419 31904 15428
rect 31852 15385 31861 15419
rect 31861 15385 31895 15419
rect 31895 15385 31904 15419
rect 31852 15376 31904 15385
rect 34796 15444 34848 15496
rect 36912 15444 36964 15496
rect 38568 15487 38620 15496
rect 38568 15453 38577 15487
rect 38577 15453 38611 15487
rect 38611 15453 38620 15487
rect 38568 15444 38620 15453
rect 31484 15308 31536 15360
rect 32128 15351 32180 15360
rect 32128 15317 32137 15351
rect 32137 15317 32171 15351
rect 32171 15317 32180 15351
rect 32128 15308 32180 15317
rect 33232 15376 33284 15428
rect 37464 15376 37516 15428
rect 39120 15444 39172 15496
rect 39396 15444 39448 15496
rect 33048 15308 33100 15360
rect 33876 15308 33928 15360
rect 36084 15308 36136 15360
rect 38660 15308 38712 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 4620 15147 4672 15156
rect 4620 15113 4629 15147
rect 4629 15113 4663 15147
rect 4663 15113 4672 15147
rect 4620 15104 4672 15113
rect 5540 15104 5592 15156
rect 5724 15104 5776 15156
rect 5264 14968 5316 15020
rect 4620 14900 4672 14952
rect 5908 14968 5960 15020
rect 6000 15011 6052 15020
rect 6000 14977 6009 15011
rect 6009 14977 6043 15011
rect 6043 14977 6052 15011
rect 6000 14968 6052 14977
rect 6828 15036 6880 15088
rect 7012 15036 7064 15088
rect 6460 14764 6512 14816
rect 6920 14900 6972 14952
rect 7840 15104 7892 15156
rect 8484 15104 8536 15156
rect 8944 15104 8996 15156
rect 7564 14968 7616 15020
rect 7932 14968 7984 15020
rect 8024 14968 8076 15020
rect 8576 14968 8628 15020
rect 10232 15104 10284 15156
rect 9220 15036 9272 15088
rect 9404 15011 9456 15020
rect 9404 14977 9413 15011
rect 9413 14977 9447 15011
rect 9447 14977 9456 15011
rect 9404 14968 9456 14977
rect 9864 14968 9916 15020
rect 7012 14875 7064 14884
rect 7012 14841 7021 14875
rect 7021 14841 7055 14875
rect 7055 14841 7064 14875
rect 7012 14832 7064 14841
rect 7196 14807 7248 14816
rect 7196 14773 7205 14807
rect 7205 14773 7239 14807
rect 7239 14773 7248 14807
rect 7196 14764 7248 14773
rect 7288 14807 7340 14816
rect 7288 14773 7297 14807
rect 7297 14773 7331 14807
rect 7331 14773 7340 14807
rect 7288 14764 7340 14773
rect 7472 14807 7524 14816
rect 7472 14773 7481 14807
rect 7481 14773 7515 14807
rect 7515 14773 7524 14807
rect 7472 14764 7524 14773
rect 8116 14764 8168 14816
rect 9496 14900 9548 14952
rect 10232 14943 10284 14952
rect 10232 14909 10241 14943
rect 10241 14909 10275 14943
rect 10275 14909 10284 14943
rect 10232 14900 10284 14909
rect 10324 14943 10376 14952
rect 10324 14909 10333 14943
rect 10333 14909 10367 14943
rect 10367 14909 10376 14943
rect 10324 14900 10376 14909
rect 10784 15011 10836 15020
rect 10784 14977 10793 15011
rect 10793 14977 10827 15011
rect 10827 14977 10836 15011
rect 10784 14968 10836 14977
rect 11612 14900 11664 14952
rect 12532 15036 12584 15088
rect 13360 15104 13412 15156
rect 12440 15011 12492 15020
rect 12440 14977 12449 15011
rect 12449 14977 12483 15011
rect 12483 14977 12492 15011
rect 12440 14968 12492 14977
rect 13452 15036 13504 15088
rect 16764 15036 16816 15088
rect 17500 15036 17552 15088
rect 17868 15079 17920 15088
rect 17868 15045 17877 15079
rect 17877 15045 17911 15079
rect 17911 15045 17920 15079
rect 17868 15036 17920 15045
rect 18144 15036 18196 15088
rect 12716 15011 12768 15020
rect 12716 14977 12725 15011
rect 12725 14977 12759 15011
rect 12759 14977 12768 15011
rect 12716 14968 12768 14977
rect 12900 14968 12952 15020
rect 13176 15011 13228 15020
rect 13176 14977 13185 15011
rect 13185 14977 13219 15011
rect 13219 14977 13228 15011
rect 13176 14968 13228 14977
rect 13268 14968 13320 15020
rect 12072 14943 12124 14952
rect 12072 14909 12081 14943
rect 12081 14909 12115 14943
rect 12115 14909 12124 14943
rect 12072 14900 12124 14909
rect 15108 15011 15160 15020
rect 15108 14977 15117 15011
rect 15117 14977 15151 15011
rect 15151 14977 15160 15011
rect 15108 14968 15160 14977
rect 15844 15011 15896 15020
rect 15844 14977 15853 15011
rect 15853 14977 15887 15011
rect 15887 14977 15896 15011
rect 15844 14968 15896 14977
rect 16488 14968 16540 15020
rect 16856 15011 16908 15020
rect 16856 14977 16865 15011
rect 16865 14977 16899 15011
rect 16899 14977 16908 15011
rect 16856 14968 16908 14977
rect 19340 14968 19392 15020
rect 19616 14968 19668 15020
rect 19800 15011 19852 15020
rect 19800 14977 19809 15011
rect 19809 14977 19843 15011
rect 19843 14977 19852 15011
rect 19800 14968 19852 14977
rect 19984 15011 20036 15020
rect 19984 14977 19993 15011
rect 19993 14977 20027 15011
rect 20027 14977 20036 15011
rect 19984 14968 20036 14977
rect 20168 15079 20220 15088
rect 20168 15045 20177 15079
rect 20177 15045 20211 15079
rect 20211 15045 20220 15079
rect 20168 15036 20220 15045
rect 20628 15104 20680 15156
rect 22652 15104 22704 15156
rect 23112 15104 23164 15156
rect 24676 15104 24728 15156
rect 21272 15036 21324 15088
rect 21548 15036 21600 15088
rect 10140 14764 10192 14816
rect 11704 14764 11756 14816
rect 12900 14807 12952 14816
rect 12900 14773 12909 14807
rect 12909 14773 12943 14807
rect 12943 14773 12952 14807
rect 12900 14764 12952 14773
rect 13636 14807 13688 14816
rect 13636 14773 13645 14807
rect 13645 14773 13679 14807
rect 13679 14773 13688 14807
rect 13636 14764 13688 14773
rect 14832 14832 14884 14884
rect 17040 14943 17092 14952
rect 17040 14909 17049 14943
rect 17049 14909 17083 14943
rect 17083 14909 17092 14943
rect 17040 14900 17092 14909
rect 17960 14900 18012 14952
rect 20444 14900 20496 14952
rect 21272 14900 21324 14952
rect 18696 14832 18748 14884
rect 21180 14832 21232 14884
rect 22284 14968 22336 15020
rect 22836 15011 22888 15020
rect 22836 14977 22845 15011
rect 22845 14977 22879 15011
rect 22879 14977 22888 15011
rect 22836 14968 22888 14977
rect 24216 14968 24268 15020
rect 24676 14968 24728 15020
rect 25136 15036 25188 15088
rect 31024 15104 31076 15156
rect 31760 15104 31812 15156
rect 33968 15104 34020 15156
rect 34980 15104 35032 15156
rect 30288 15036 30340 15088
rect 33140 15036 33192 15088
rect 35440 15036 35492 15088
rect 38476 15104 38528 15156
rect 39028 15104 39080 15156
rect 22652 14900 22704 14952
rect 24400 14900 24452 14952
rect 24492 14900 24544 14952
rect 29000 14968 29052 15020
rect 31484 14900 31536 14952
rect 33968 14968 34020 15020
rect 35348 14968 35400 15020
rect 38660 15011 38712 15020
rect 38660 14977 38669 15011
rect 38669 14977 38703 15011
rect 38703 14977 38712 15011
rect 38660 14968 38712 14977
rect 38844 15011 38896 15020
rect 38844 14977 38853 15011
rect 38853 14977 38887 15011
rect 38887 14977 38896 15011
rect 38844 14968 38896 14977
rect 34612 14900 34664 14952
rect 24676 14832 24728 14884
rect 27712 14832 27764 14884
rect 33324 14832 33376 14884
rect 37556 14832 37608 14884
rect 14740 14807 14792 14816
rect 14740 14773 14749 14807
rect 14749 14773 14783 14807
rect 14783 14773 14792 14807
rect 14740 14764 14792 14773
rect 16488 14764 16540 14816
rect 17776 14807 17828 14816
rect 17776 14773 17785 14807
rect 17785 14773 17819 14807
rect 17819 14773 17828 14807
rect 17776 14764 17828 14773
rect 19524 14807 19576 14816
rect 19524 14773 19533 14807
rect 19533 14773 19567 14807
rect 19567 14773 19576 14807
rect 19524 14764 19576 14773
rect 20720 14764 20772 14816
rect 20812 14764 20864 14816
rect 22928 14764 22980 14816
rect 24400 14764 24452 14816
rect 34060 14764 34112 14816
rect 34428 14764 34480 14816
rect 38660 14807 38712 14816
rect 38660 14773 38669 14807
rect 38669 14773 38703 14807
rect 38703 14773 38712 14807
rect 38660 14764 38712 14773
rect 39028 14807 39080 14816
rect 39028 14773 39037 14807
rect 39037 14773 39071 14807
rect 39071 14773 39080 14807
rect 39028 14764 39080 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 5816 14560 5868 14612
rect 6276 14603 6328 14612
rect 6276 14569 6285 14603
rect 6285 14569 6319 14603
rect 6319 14569 6328 14603
rect 6276 14560 6328 14569
rect 7012 14560 7064 14612
rect 4620 14535 4672 14544
rect 4620 14501 4629 14535
rect 4629 14501 4663 14535
rect 4663 14501 4672 14535
rect 4620 14492 4672 14501
rect 4252 14467 4304 14476
rect 4252 14433 4261 14467
rect 4261 14433 4295 14467
rect 4295 14433 4304 14467
rect 4252 14424 4304 14433
rect 4344 14356 4396 14408
rect 4712 14356 4764 14408
rect 5908 14399 5960 14408
rect 5908 14365 5917 14399
rect 5917 14365 5951 14399
rect 5951 14365 5960 14399
rect 5908 14356 5960 14365
rect 6000 14263 6052 14272
rect 6000 14229 6009 14263
rect 6009 14229 6043 14263
rect 6043 14229 6052 14263
rect 6000 14220 6052 14229
rect 6460 14467 6512 14476
rect 6460 14433 6469 14467
rect 6469 14433 6503 14467
rect 6503 14433 6512 14467
rect 6460 14424 6512 14433
rect 6552 14467 6604 14476
rect 6552 14433 6561 14467
rect 6561 14433 6595 14467
rect 6595 14433 6604 14467
rect 6552 14424 6604 14433
rect 6828 14424 6880 14476
rect 7104 14356 7156 14408
rect 7196 14399 7248 14408
rect 7196 14365 7205 14399
rect 7205 14365 7239 14399
rect 7239 14365 7248 14399
rect 7196 14356 7248 14365
rect 7564 14424 7616 14476
rect 9128 14492 9180 14544
rect 9404 14560 9456 14612
rect 9496 14560 9548 14612
rect 9956 14560 10008 14612
rect 10140 14560 10192 14612
rect 10324 14560 10376 14612
rect 10784 14560 10836 14612
rect 14740 14560 14792 14612
rect 15660 14603 15712 14612
rect 15660 14569 15669 14603
rect 15669 14569 15703 14603
rect 15703 14569 15712 14603
rect 15660 14560 15712 14569
rect 15844 14603 15896 14612
rect 15844 14569 15853 14603
rect 15853 14569 15887 14603
rect 15887 14569 15896 14603
rect 15844 14560 15896 14569
rect 16028 14603 16080 14612
rect 16028 14569 16037 14603
rect 16037 14569 16071 14603
rect 16071 14569 16080 14603
rect 16028 14560 16080 14569
rect 17960 14560 18012 14612
rect 18236 14560 18288 14612
rect 18880 14560 18932 14612
rect 19524 14603 19576 14612
rect 19524 14569 19533 14603
rect 19533 14569 19567 14603
rect 19567 14569 19576 14603
rect 19524 14560 19576 14569
rect 19800 14603 19852 14612
rect 19800 14569 19809 14603
rect 19809 14569 19843 14603
rect 19843 14569 19852 14603
rect 19800 14560 19852 14569
rect 20628 14560 20680 14612
rect 8760 14424 8812 14476
rect 6828 14288 6880 14340
rect 7564 14331 7616 14340
rect 7564 14297 7573 14331
rect 7573 14297 7607 14331
rect 7607 14297 7616 14331
rect 7564 14288 7616 14297
rect 8484 14399 8536 14408
rect 8484 14365 8493 14399
rect 8493 14365 8527 14399
rect 8527 14365 8536 14399
rect 8484 14356 8536 14365
rect 8576 14399 8628 14408
rect 8576 14365 8585 14399
rect 8585 14365 8619 14399
rect 8619 14365 8628 14399
rect 8576 14356 8628 14365
rect 8668 14399 8720 14408
rect 8668 14365 8677 14399
rect 8677 14365 8711 14399
rect 8711 14365 8720 14399
rect 8668 14356 8720 14365
rect 9496 14399 9548 14408
rect 9496 14365 9500 14399
rect 9500 14365 9534 14399
rect 9534 14365 9548 14399
rect 9496 14356 9548 14365
rect 9680 14399 9732 14408
rect 9680 14365 9689 14399
rect 9689 14365 9723 14399
rect 9723 14365 9732 14399
rect 9680 14356 9732 14365
rect 10140 14424 10192 14476
rect 9956 14399 10008 14408
rect 9956 14365 9965 14399
rect 9965 14365 9999 14399
rect 9999 14365 10008 14399
rect 9956 14356 10008 14365
rect 10048 14399 10100 14408
rect 10048 14365 10057 14399
rect 10057 14365 10091 14399
rect 10091 14365 10100 14399
rect 10048 14356 10100 14365
rect 15752 14492 15804 14544
rect 15936 14492 15988 14544
rect 10416 14356 10468 14408
rect 11612 14356 11664 14408
rect 16856 14424 16908 14476
rect 17592 14424 17644 14476
rect 18696 14467 18748 14476
rect 18696 14433 18705 14467
rect 18705 14433 18739 14467
rect 18739 14433 18748 14467
rect 18696 14424 18748 14433
rect 18880 14467 18932 14476
rect 18880 14433 18889 14467
rect 18889 14433 18923 14467
rect 18923 14433 18932 14467
rect 18880 14424 18932 14433
rect 20168 14492 20220 14544
rect 19800 14424 19852 14476
rect 21180 14424 21232 14476
rect 7380 14220 7432 14272
rect 8208 14263 8260 14272
rect 8208 14229 8217 14263
rect 8217 14229 8251 14263
rect 8251 14229 8260 14263
rect 8208 14220 8260 14229
rect 8668 14220 8720 14272
rect 9404 14220 9456 14272
rect 12992 14288 13044 14340
rect 10416 14263 10468 14272
rect 10416 14229 10425 14263
rect 10425 14229 10459 14263
rect 10459 14229 10468 14263
rect 10416 14220 10468 14229
rect 11888 14220 11940 14272
rect 12072 14220 12124 14272
rect 13176 14220 13228 14272
rect 15292 14288 15344 14340
rect 15568 14399 15620 14408
rect 15568 14365 15577 14399
rect 15577 14365 15611 14399
rect 15611 14365 15620 14399
rect 15568 14356 15620 14365
rect 15936 14356 15988 14408
rect 16764 14356 16816 14408
rect 17316 14356 17368 14408
rect 19616 14399 19668 14408
rect 19616 14365 19625 14399
rect 19625 14365 19659 14399
rect 19659 14365 19668 14399
rect 19616 14356 19668 14365
rect 20168 14356 20220 14408
rect 20536 14399 20588 14408
rect 20536 14365 20545 14399
rect 20545 14365 20579 14399
rect 20579 14365 20588 14399
rect 20536 14356 20588 14365
rect 21732 14492 21784 14544
rect 22192 14603 22244 14612
rect 22192 14569 22201 14603
rect 22201 14569 22235 14603
rect 22235 14569 22244 14603
rect 22192 14560 22244 14569
rect 22652 14603 22704 14612
rect 22652 14569 22661 14603
rect 22661 14569 22695 14603
rect 22695 14569 22704 14603
rect 22652 14560 22704 14569
rect 24952 14560 25004 14612
rect 25504 14560 25556 14612
rect 27804 14560 27856 14612
rect 28540 14603 28592 14612
rect 28540 14569 28549 14603
rect 28549 14569 28583 14603
rect 28583 14569 28592 14603
rect 28540 14560 28592 14569
rect 22836 14492 22888 14544
rect 24032 14492 24084 14544
rect 27252 14492 27304 14544
rect 13452 14220 13504 14272
rect 16764 14220 16816 14272
rect 18972 14288 19024 14340
rect 20352 14288 20404 14340
rect 21272 14288 21324 14340
rect 21732 14399 21784 14408
rect 21732 14365 21741 14399
rect 21741 14365 21775 14399
rect 21775 14365 21784 14399
rect 21732 14356 21784 14365
rect 22100 14356 22152 14408
rect 22744 14399 22796 14408
rect 22744 14365 22753 14399
rect 22753 14365 22787 14399
rect 22787 14365 22796 14399
rect 22744 14356 22796 14365
rect 23572 14424 23624 14476
rect 24308 14424 24360 14476
rect 24952 14424 25004 14476
rect 25320 14424 25372 14476
rect 22468 14331 22520 14340
rect 22468 14297 22477 14331
rect 22477 14297 22511 14331
rect 22511 14297 22520 14331
rect 23112 14399 23164 14408
rect 23112 14365 23121 14399
rect 23121 14365 23155 14399
rect 23155 14365 23164 14399
rect 23112 14356 23164 14365
rect 24584 14356 24636 14408
rect 24676 14356 24728 14408
rect 25044 14399 25096 14408
rect 25044 14365 25053 14399
rect 25053 14365 25087 14399
rect 25087 14365 25096 14399
rect 25044 14356 25096 14365
rect 25872 14356 25924 14408
rect 25964 14399 26016 14408
rect 25964 14365 25973 14399
rect 25973 14365 26007 14399
rect 26007 14365 26016 14399
rect 25964 14356 26016 14365
rect 27436 14356 27488 14408
rect 22468 14288 22520 14297
rect 17408 14220 17460 14272
rect 17868 14220 17920 14272
rect 20536 14220 20588 14272
rect 23756 14220 23808 14272
rect 23940 14220 23992 14272
rect 26424 14263 26476 14272
rect 26424 14229 26433 14263
rect 26433 14229 26467 14263
rect 26467 14229 26476 14263
rect 26424 14220 26476 14229
rect 26608 14220 26660 14272
rect 28080 14399 28132 14408
rect 28080 14365 28089 14399
rect 28089 14365 28123 14399
rect 28123 14365 28132 14399
rect 28080 14356 28132 14365
rect 27712 14288 27764 14340
rect 28264 14399 28316 14408
rect 28264 14365 28273 14399
rect 28273 14365 28307 14399
rect 28307 14365 28316 14399
rect 28264 14356 28316 14365
rect 29000 14560 29052 14612
rect 35900 14560 35952 14612
rect 36084 14560 36136 14612
rect 36452 14560 36504 14612
rect 37464 14560 37516 14612
rect 28908 14535 28960 14544
rect 28908 14501 28917 14535
rect 28917 14501 28951 14535
rect 28951 14501 28960 14535
rect 28908 14492 28960 14501
rect 29644 14492 29696 14544
rect 28540 14288 28592 14340
rect 28908 14356 28960 14408
rect 29000 14399 29052 14408
rect 29000 14365 29009 14399
rect 29009 14365 29043 14399
rect 29043 14365 29052 14399
rect 29000 14356 29052 14365
rect 31024 14424 31076 14476
rect 33600 14424 33652 14476
rect 30472 14356 30524 14408
rect 35900 14356 35952 14408
rect 32956 14288 33008 14340
rect 36636 14356 36688 14408
rect 36820 14356 36872 14408
rect 30380 14220 30432 14272
rect 30564 14220 30616 14272
rect 35348 14220 35400 14272
rect 37280 14263 37332 14272
rect 37280 14229 37289 14263
rect 37289 14229 37323 14263
rect 37323 14229 37332 14263
rect 37280 14220 37332 14229
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 4252 14016 4304 14068
rect 6000 14016 6052 14068
rect 7564 14016 7616 14068
rect 4160 13880 4212 13932
rect 4528 13880 4580 13932
rect 5908 13948 5960 14000
rect 7104 13948 7156 14000
rect 8668 13948 8720 14000
rect 4712 13923 4764 13932
rect 4712 13889 4721 13923
rect 4721 13889 4755 13923
rect 4755 13889 4764 13923
rect 4712 13880 4764 13889
rect 10140 14016 10192 14068
rect 9956 13948 10008 14000
rect 9772 13880 9824 13932
rect 10416 13880 10468 13932
rect 10508 13923 10560 13932
rect 10508 13889 10517 13923
rect 10517 13889 10551 13923
rect 10551 13889 10560 13923
rect 10508 13880 10560 13889
rect 13176 14016 13228 14068
rect 16672 14016 16724 14068
rect 16764 14016 16816 14068
rect 20076 14016 20128 14068
rect 21732 14016 21784 14068
rect 12532 13948 12584 14000
rect 16212 13991 16264 14000
rect 16212 13957 16221 13991
rect 16221 13957 16255 13991
rect 16255 13957 16264 13991
rect 16212 13948 16264 13957
rect 17224 13948 17276 14000
rect 17868 13948 17920 14000
rect 18972 13948 19024 14000
rect 7288 13812 7340 13864
rect 11060 13923 11112 13932
rect 11060 13889 11069 13923
rect 11069 13889 11103 13923
rect 11103 13889 11112 13923
rect 11060 13880 11112 13889
rect 11520 13880 11572 13932
rect 4344 13744 4396 13796
rect 5172 13744 5224 13796
rect 5724 13744 5776 13796
rect 9864 13744 9916 13796
rect 10968 13812 11020 13864
rect 12348 13880 12400 13932
rect 12624 13923 12676 13932
rect 12624 13889 12633 13923
rect 12633 13889 12667 13923
rect 12667 13889 12676 13923
rect 12624 13880 12676 13889
rect 12808 13923 12860 13932
rect 12808 13889 12817 13923
rect 12817 13889 12851 13923
rect 12851 13889 12860 13923
rect 12808 13880 12860 13889
rect 12992 13880 13044 13932
rect 13268 13880 13320 13932
rect 13360 13923 13412 13932
rect 13360 13889 13369 13923
rect 13369 13889 13403 13923
rect 13403 13889 13412 13923
rect 13360 13880 13412 13889
rect 12440 13812 12492 13864
rect 11060 13744 11112 13796
rect 12716 13744 12768 13796
rect 13636 13812 13688 13864
rect 14464 13880 14516 13932
rect 9220 13719 9272 13728
rect 9220 13685 9229 13719
rect 9229 13685 9263 13719
rect 9263 13685 9272 13719
rect 9220 13676 9272 13685
rect 10232 13719 10284 13728
rect 10232 13685 10241 13719
rect 10241 13685 10275 13719
rect 10275 13685 10284 13719
rect 10232 13676 10284 13685
rect 11796 13676 11848 13728
rect 12440 13719 12492 13728
rect 12440 13685 12449 13719
rect 12449 13685 12483 13719
rect 12483 13685 12492 13719
rect 12440 13676 12492 13685
rect 12808 13676 12860 13728
rect 13084 13676 13136 13728
rect 14096 13719 14148 13728
rect 14096 13685 14105 13719
rect 14105 13685 14139 13719
rect 14139 13685 14148 13719
rect 14096 13676 14148 13685
rect 15200 13744 15252 13796
rect 15568 13744 15620 13796
rect 19248 13880 19300 13932
rect 19892 13880 19944 13932
rect 20352 13948 20404 14000
rect 22284 14016 22336 14068
rect 23756 14016 23808 14068
rect 23940 14016 23992 14068
rect 24216 14016 24268 14068
rect 24308 14059 24360 14068
rect 24308 14025 24317 14059
rect 24317 14025 24351 14059
rect 24351 14025 24360 14059
rect 24308 14016 24360 14025
rect 24492 14059 24544 14068
rect 24492 14025 24519 14059
rect 24519 14025 24544 14059
rect 24492 14016 24544 14025
rect 25964 14016 26016 14068
rect 22008 13948 22060 14000
rect 24124 13948 24176 14000
rect 24676 13991 24728 14000
rect 24676 13957 24685 13991
rect 24685 13957 24719 13991
rect 24719 13957 24728 13991
rect 24676 13948 24728 13957
rect 20720 13880 20772 13932
rect 23020 13880 23072 13932
rect 20168 13812 20220 13864
rect 18604 13744 18656 13796
rect 19892 13744 19944 13796
rect 20260 13744 20312 13796
rect 22100 13812 22152 13864
rect 23112 13812 23164 13864
rect 25044 13880 25096 13932
rect 26240 13948 26292 14000
rect 26700 14016 26752 14068
rect 27068 14059 27120 14068
rect 27068 14025 27077 14059
rect 27077 14025 27111 14059
rect 27111 14025 27120 14059
rect 27068 14016 27120 14025
rect 28264 14016 28316 14068
rect 27252 13948 27304 14000
rect 32956 14016 33008 14068
rect 28448 13991 28500 14000
rect 28448 13957 28457 13991
rect 28457 13957 28491 13991
rect 28491 13957 28500 13991
rect 28448 13948 28500 13957
rect 28540 13948 28592 14000
rect 28724 13948 28776 14000
rect 32036 13948 32088 14000
rect 32220 13948 32272 14000
rect 37004 14016 37056 14068
rect 39212 14016 39264 14068
rect 21272 13744 21324 13796
rect 22836 13744 22888 13796
rect 24124 13812 24176 13864
rect 24492 13812 24544 13864
rect 26056 13812 26108 13864
rect 26516 13855 26568 13864
rect 26516 13821 26525 13855
rect 26525 13821 26559 13855
rect 26559 13821 26568 13855
rect 26516 13812 26568 13821
rect 26700 13855 26752 13864
rect 26700 13821 26709 13855
rect 26709 13821 26743 13855
rect 26743 13821 26752 13855
rect 26700 13812 26752 13821
rect 27436 13880 27488 13932
rect 28080 13880 28132 13932
rect 27252 13812 27304 13864
rect 27620 13812 27672 13864
rect 28816 13880 28868 13932
rect 29552 13880 29604 13932
rect 30564 13923 30616 13932
rect 30564 13889 30573 13923
rect 30573 13889 30607 13923
rect 30607 13889 30616 13923
rect 30564 13880 30616 13889
rect 31392 13880 31444 13932
rect 31576 13880 31628 13932
rect 30288 13812 30340 13864
rect 30748 13812 30800 13864
rect 32772 13923 32824 13932
rect 32772 13889 32781 13923
rect 32781 13889 32815 13923
rect 32815 13889 32824 13923
rect 32772 13880 32824 13889
rect 34704 13948 34756 14000
rect 36084 13948 36136 14000
rect 36820 13948 36872 14000
rect 37188 13948 37240 14000
rect 36728 13923 36780 13932
rect 36728 13889 36737 13923
rect 36737 13889 36771 13923
rect 36771 13889 36780 13923
rect 36728 13880 36780 13889
rect 36912 13923 36964 13932
rect 36912 13889 36921 13923
rect 36921 13889 36955 13923
rect 36955 13889 36964 13923
rect 36912 13880 36964 13889
rect 18236 13676 18288 13728
rect 19524 13676 19576 13728
rect 23940 13676 23992 13728
rect 24492 13719 24544 13728
rect 24492 13685 24501 13719
rect 24501 13685 24535 13719
rect 24535 13685 24544 13719
rect 24492 13676 24544 13685
rect 27160 13744 27212 13796
rect 27804 13744 27856 13796
rect 28080 13676 28132 13728
rect 29000 13744 29052 13796
rect 32956 13812 33008 13864
rect 33232 13744 33284 13796
rect 33600 13812 33652 13864
rect 39396 13948 39448 14000
rect 37464 13923 37516 13932
rect 37464 13889 37473 13923
rect 37473 13889 37507 13923
rect 37507 13889 37516 13923
rect 37464 13880 37516 13889
rect 37556 13923 37608 13932
rect 37556 13889 37565 13923
rect 37565 13889 37599 13923
rect 37599 13889 37608 13923
rect 37556 13880 37608 13889
rect 38384 13923 38436 13932
rect 38384 13889 38393 13923
rect 38393 13889 38427 13923
rect 38427 13889 38436 13923
rect 38384 13880 38436 13889
rect 37648 13812 37700 13864
rect 36820 13744 36872 13796
rect 29184 13676 29236 13728
rect 30748 13676 30800 13728
rect 32128 13676 32180 13728
rect 32588 13719 32640 13728
rect 32588 13685 32597 13719
rect 32597 13685 32631 13719
rect 32631 13685 32640 13719
rect 32588 13676 32640 13685
rect 38108 13744 38160 13796
rect 39764 13880 39816 13932
rect 38844 13744 38896 13796
rect 39488 13744 39540 13796
rect 37280 13719 37332 13728
rect 37280 13685 37289 13719
rect 37289 13685 37323 13719
rect 37323 13685 37332 13719
rect 37280 13676 37332 13685
rect 38568 13719 38620 13728
rect 38568 13685 38577 13719
rect 38577 13685 38611 13719
rect 38611 13685 38620 13719
rect 38568 13676 38620 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 4068 13472 4120 13524
rect 4620 13472 4672 13524
rect 4160 13404 4212 13456
rect 5356 13472 5408 13524
rect 5908 13472 5960 13524
rect 9220 13472 9272 13524
rect 16028 13472 16080 13524
rect 16672 13472 16724 13524
rect 16856 13515 16908 13524
rect 16856 13481 16865 13515
rect 16865 13481 16899 13515
rect 16899 13481 16908 13515
rect 16856 13472 16908 13481
rect 17040 13515 17092 13524
rect 17040 13481 17049 13515
rect 17049 13481 17083 13515
rect 17083 13481 17092 13515
rect 17040 13472 17092 13481
rect 17224 13515 17276 13524
rect 17224 13481 17233 13515
rect 17233 13481 17267 13515
rect 17267 13481 17276 13515
rect 17224 13472 17276 13481
rect 17960 13515 18012 13524
rect 17960 13481 17969 13515
rect 17969 13481 18003 13515
rect 18003 13481 18012 13515
rect 17960 13472 18012 13481
rect 8116 13404 8168 13456
rect 3976 13268 4028 13320
rect 3792 13243 3844 13252
rect 3792 13209 3801 13243
rect 3801 13209 3835 13243
rect 3835 13209 3844 13243
rect 3792 13200 3844 13209
rect 4160 13243 4212 13252
rect 4160 13209 4169 13243
rect 4169 13209 4203 13243
rect 4203 13209 4212 13243
rect 4160 13200 4212 13209
rect 4620 13268 4672 13320
rect 4804 13311 4856 13320
rect 4804 13277 4813 13311
rect 4813 13277 4847 13311
rect 4847 13277 4856 13311
rect 4804 13268 4856 13277
rect 7472 13336 7524 13388
rect 5172 13311 5224 13320
rect 5172 13277 5181 13311
rect 5181 13277 5215 13311
rect 5215 13277 5224 13311
rect 5172 13268 5224 13277
rect 5816 13268 5868 13320
rect 6644 13268 6696 13320
rect 7104 13311 7156 13320
rect 7104 13277 7113 13311
rect 7113 13277 7147 13311
rect 7147 13277 7156 13311
rect 7104 13268 7156 13277
rect 7748 13268 7800 13320
rect 8208 13336 8260 13388
rect 9864 13404 9916 13456
rect 11060 13404 11112 13456
rect 9772 13379 9824 13388
rect 9772 13345 9781 13379
rect 9781 13345 9815 13379
rect 9815 13345 9824 13379
rect 9772 13336 9824 13345
rect 11520 13336 11572 13388
rect 12256 13336 12308 13388
rect 7472 13200 7524 13252
rect 8024 13268 8076 13320
rect 8760 13268 8812 13320
rect 9956 13311 10008 13320
rect 9956 13277 9965 13311
rect 9965 13277 9999 13311
rect 9999 13277 10008 13311
rect 9956 13268 10008 13277
rect 8208 13243 8260 13252
rect 8208 13209 8217 13243
rect 8217 13209 8251 13243
rect 8251 13209 8260 13243
rect 8208 13200 8260 13209
rect 11336 13200 11388 13252
rect 11520 13243 11572 13252
rect 11520 13209 11529 13243
rect 11529 13209 11563 13243
rect 11563 13209 11572 13243
rect 11520 13200 11572 13209
rect 4804 13132 4856 13184
rect 5540 13132 5592 13184
rect 6460 13132 6512 13184
rect 7748 13175 7800 13184
rect 7748 13141 7757 13175
rect 7757 13141 7791 13175
rect 7791 13141 7800 13175
rect 7748 13132 7800 13141
rect 8300 13132 8352 13184
rect 8668 13132 8720 13184
rect 12348 13268 12400 13320
rect 12716 13268 12768 13320
rect 12808 13311 12860 13320
rect 12808 13277 12817 13311
rect 12817 13277 12851 13311
rect 12851 13277 12860 13311
rect 12808 13268 12860 13277
rect 13176 13379 13228 13388
rect 13176 13345 13185 13379
rect 13185 13345 13219 13379
rect 13219 13345 13228 13379
rect 13176 13336 13228 13345
rect 14740 13336 14792 13388
rect 21732 13472 21784 13524
rect 13084 13311 13136 13320
rect 13084 13277 13093 13311
rect 13093 13277 13127 13311
rect 13127 13277 13136 13311
rect 13084 13268 13136 13277
rect 13176 13200 13228 13252
rect 14372 13311 14424 13320
rect 14372 13277 14381 13311
rect 14381 13277 14415 13311
rect 14415 13277 14424 13311
rect 14372 13268 14424 13277
rect 15200 13311 15252 13320
rect 15200 13277 15209 13311
rect 15209 13277 15243 13311
rect 15243 13277 15252 13311
rect 15200 13268 15252 13277
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 16672 13311 16724 13320
rect 16672 13277 16681 13311
rect 16681 13277 16715 13311
rect 16715 13277 16724 13311
rect 16672 13268 16724 13277
rect 16764 13268 16816 13320
rect 17224 13311 17276 13320
rect 17224 13277 17233 13311
rect 17233 13277 17267 13311
rect 17267 13277 17276 13311
rect 17224 13268 17276 13277
rect 12440 13132 12492 13184
rect 12992 13132 13044 13184
rect 13728 13132 13780 13184
rect 13820 13132 13872 13184
rect 15660 13132 15712 13184
rect 17132 13200 17184 13252
rect 17408 13268 17460 13320
rect 17500 13243 17552 13252
rect 17500 13209 17509 13243
rect 17509 13209 17543 13243
rect 17543 13209 17552 13243
rect 17500 13200 17552 13209
rect 17592 13132 17644 13184
rect 17868 13311 17920 13320
rect 17868 13277 17877 13311
rect 17877 13277 17911 13311
rect 17911 13277 17920 13311
rect 17868 13268 17920 13277
rect 17960 13268 18012 13320
rect 18512 13268 18564 13320
rect 18604 13268 18656 13320
rect 18972 13200 19024 13252
rect 19340 13311 19392 13320
rect 19340 13277 19349 13311
rect 19349 13277 19383 13311
rect 19383 13277 19392 13311
rect 19340 13268 19392 13277
rect 20720 13336 20772 13388
rect 21732 13336 21784 13388
rect 22100 13336 22152 13388
rect 18512 13132 18564 13184
rect 18880 13132 18932 13184
rect 19984 13268 20036 13320
rect 20076 13311 20128 13320
rect 20076 13277 20085 13311
rect 20085 13277 20119 13311
rect 20119 13277 20128 13311
rect 20076 13268 20128 13277
rect 20352 13311 20404 13320
rect 20352 13277 20361 13311
rect 20361 13277 20395 13311
rect 20395 13277 20404 13311
rect 20352 13268 20404 13277
rect 20904 13311 20956 13320
rect 20904 13277 20913 13311
rect 20913 13277 20947 13311
rect 20947 13277 20956 13311
rect 20904 13268 20956 13277
rect 19800 13243 19852 13252
rect 19800 13209 19809 13243
rect 19809 13209 19843 13243
rect 19843 13209 19852 13243
rect 19800 13200 19852 13209
rect 20628 13200 20680 13252
rect 21180 13311 21232 13320
rect 21180 13277 21189 13311
rect 21189 13277 21223 13311
rect 21223 13277 21232 13311
rect 21180 13268 21232 13277
rect 21548 13268 21600 13320
rect 22376 13404 22428 13456
rect 22376 13311 22428 13320
rect 22376 13277 22385 13311
rect 22385 13277 22419 13311
rect 22419 13277 22428 13311
rect 22376 13268 22428 13277
rect 23020 13515 23072 13524
rect 23020 13481 23029 13515
rect 23029 13481 23063 13515
rect 23063 13481 23072 13515
rect 23020 13472 23072 13481
rect 23756 13472 23808 13524
rect 26332 13472 26384 13524
rect 30472 13472 30524 13524
rect 22744 13404 22796 13456
rect 27528 13404 27580 13456
rect 28264 13404 28316 13456
rect 31760 13472 31812 13524
rect 32128 13472 32180 13524
rect 32404 13472 32456 13524
rect 34152 13472 34204 13524
rect 36728 13472 36780 13524
rect 36820 13472 36872 13524
rect 22928 13336 22980 13388
rect 31852 13404 31904 13456
rect 32772 13404 32824 13456
rect 32864 13404 32916 13456
rect 33232 13404 33284 13456
rect 38936 13515 38988 13524
rect 38936 13481 38945 13515
rect 38945 13481 38979 13515
rect 38979 13481 38988 13515
rect 38936 13472 38988 13481
rect 21548 13175 21600 13184
rect 21548 13141 21557 13175
rect 21557 13141 21591 13175
rect 21591 13141 21600 13175
rect 21548 13132 21600 13141
rect 22836 13268 22888 13320
rect 26148 13311 26200 13320
rect 26148 13277 26157 13311
rect 26157 13277 26191 13311
rect 26191 13277 26200 13311
rect 26148 13268 26200 13277
rect 26240 13311 26292 13320
rect 26240 13277 26249 13311
rect 26249 13277 26283 13311
rect 26283 13277 26292 13311
rect 26240 13268 26292 13277
rect 26608 13311 26660 13320
rect 26608 13277 26617 13311
rect 26617 13277 26651 13311
rect 26651 13277 26660 13311
rect 26608 13268 26660 13277
rect 27160 13311 27212 13320
rect 27160 13277 27169 13311
rect 27169 13277 27203 13311
rect 27203 13277 27212 13311
rect 27160 13268 27212 13277
rect 23388 13200 23440 13252
rect 24860 13200 24912 13252
rect 25596 13200 25648 13252
rect 27988 13268 28040 13320
rect 22836 13132 22888 13184
rect 23020 13175 23072 13184
rect 23020 13141 23047 13175
rect 23047 13141 23072 13175
rect 23020 13132 23072 13141
rect 23112 13132 23164 13184
rect 24216 13132 24268 13184
rect 25872 13132 25924 13184
rect 27804 13200 27856 13252
rect 29276 13200 29328 13252
rect 30196 13268 30248 13320
rect 30288 13311 30340 13320
rect 30288 13277 30297 13311
rect 30297 13277 30331 13311
rect 30331 13277 30340 13311
rect 30288 13268 30340 13277
rect 31484 13268 31536 13320
rect 31852 13268 31904 13320
rect 31392 13200 31444 13252
rect 31944 13243 31996 13252
rect 31944 13209 31953 13243
rect 31953 13209 31987 13243
rect 31987 13209 31996 13243
rect 31944 13200 31996 13209
rect 27712 13132 27764 13184
rect 28356 13132 28408 13184
rect 29184 13132 29236 13184
rect 30932 13132 30984 13184
rect 31484 13132 31536 13184
rect 32496 13268 32548 13320
rect 32772 13311 32824 13320
rect 32772 13277 32781 13311
rect 32781 13277 32815 13311
rect 32815 13277 32824 13311
rect 32772 13268 32824 13277
rect 35440 13336 35492 13388
rect 38568 13336 38620 13388
rect 33232 13268 33284 13320
rect 33048 13243 33100 13252
rect 33048 13209 33057 13243
rect 33057 13209 33091 13243
rect 33091 13209 33100 13243
rect 33048 13200 33100 13209
rect 33968 13200 34020 13252
rect 32496 13175 32548 13184
rect 32496 13141 32505 13175
rect 32505 13141 32539 13175
rect 32539 13141 32548 13175
rect 32496 13132 32548 13141
rect 34704 13311 34756 13320
rect 34704 13277 34713 13311
rect 34713 13277 34747 13311
rect 34747 13277 34756 13311
rect 34704 13268 34756 13277
rect 38108 13268 38160 13320
rect 34796 13200 34848 13252
rect 35348 13132 35400 13184
rect 38108 13132 38160 13184
rect 38752 13132 38804 13184
rect 39856 13268 39908 13320
rect 39304 13132 39356 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 3240 12928 3292 12980
rect 4620 12928 4672 12980
rect 4712 12928 4764 12980
rect 6920 12928 6972 12980
rect 7748 12928 7800 12980
rect 3792 12860 3844 12912
rect 4344 12835 4396 12844
rect 4344 12801 4353 12835
rect 4353 12801 4387 12835
rect 4387 12801 4396 12835
rect 4344 12792 4396 12801
rect 4436 12835 4488 12844
rect 4436 12801 4445 12835
rect 4445 12801 4479 12835
rect 4479 12801 4488 12835
rect 4436 12792 4488 12801
rect 4620 12835 4672 12844
rect 4620 12801 4629 12835
rect 4629 12801 4663 12835
rect 4663 12801 4672 12835
rect 4620 12792 4672 12801
rect 4896 12792 4948 12844
rect 5540 12835 5592 12844
rect 5540 12801 5549 12835
rect 5549 12801 5583 12835
rect 5583 12801 5592 12835
rect 5540 12792 5592 12801
rect 7472 12860 7524 12912
rect 12440 12928 12492 12980
rect 12532 12971 12584 12980
rect 12532 12937 12541 12971
rect 12541 12937 12575 12971
rect 12575 12937 12584 12971
rect 12532 12928 12584 12937
rect 13176 12971 13228 12980
rect 13176 12937 13185 12971
rect 13185 12937 13219 12971
rect 13219 12937 13228 12971
rect 13176 12928 13228 12937
rect 5908 12792 5960 12844
rect 6920 12792 6972 12844
rect 4436 12656 4488 12708
rect 5264 12656 5316 12708
rect 5724 12767 5776 12776
rect 5724 12733 5733 12767
rect 5733 12733 5767 12767
rect 5767 12733 5776 12767
rect 5724 12724 5776 12733
rect 6736 12767 6788 12776
rect 6736 12733 6745 12767
rect 6745 12733 6779 12767
rect 6779 12733 6788 12767
rect 6736 12724 6788 12733
rect 7104 12835 7156 12844
rect 7104 12801 7113 12835
rect 7113 12801 7147 12835
rect 7147 12801 7156 12835
rect 7104 12792 7156 12801
rect 7288 12792 7340 12844
rect 11520 12860 11572 12912
rect 7840 12835 7892 12844
rect 7840 12801 7849 12835
rect 7849 12801 7883 12835
rect 7883 12801 7892 12835
rect 7840 12792 7892 12801
rect 8024 12835 8076 12844
rect 8024 12801 8033 12835
rect 8033 12801 8067 12835
rect 8067 12801 8076 12835
rect 8024 12792 8076 12801
rect 8300 12835 8352 12844
rect 8300 12801 8309 12835
rect 8309 12801 8343 12835
rect 8343 12801 8352 12835
rect 8300 12792 8352 12801
rect 8576 12835 8628 12844
rect 8576 12801 8585 12835
rect 8585 12801 8619 12835
rect 8619 12801 8628 12835
rect 8576 12792 8628 12801
rect 10232 12792 10284 12844
rect 10968 12792 11020 12844
rect 11796 12792 11848 12844
rect 9680 12724 9732 12776
rect 11060 12724 11112 12776
rect 12992 12792 13044 12844
rect 5448 12588 5500 12640
rect 5816 12631 5868 12640
rect 5816 12597 5825 12631
rect 5825 12597 5859 12631
rect 5859 12597 5868 12631
rect 7564 12656 7616 12708
rect 8668 12656 8720 12708
rect 8944 12656 8996 12708
rect 12348 12724 12400 12776
rect 11336 12656 11388 12708
rect 13360 12656 13412 12708
rect 13728 12835 13780 12844
rect 13728 12801 13737 12835
rect 13737 12801 13771 12835
rect 13771 12801 13780 12835
rect 13728 12792 13780 12801
rect 14372 12792 14424 12844
rect 14556 12835 14608 12844
rect 14556 12801 14565 12835
rect 14565 12801 14599 12835
rect 14599 12801 14608 12835
rect 14556 12792 14608 12801
rect 15384 12928 15436 12980
rect 16672 12860 16724 12912
rect 17500 12971 17552 12980
rect 17500 12937 17509 12971
rect 17509 12937 17543 12971
rect 17543 12937 17552 12971
rect 17500 12928 17552 12937
rect 17592 12928 17644 12980
rect 18604 12928 18656 12980
rect 18972 12928 19024 12980
rect 19708 12928 19760 12980
rect 20168 12928 20220 12980
rect 20812 12928 20864 12980
rect 20996 12971 21048 12980
rect 20996 12937 21005 12971
rect 21005 12937 21039 12971
rect 21039 12937 21048 12971
rect 20996 12928 21048 12937
rect 21088 12928 21140 12980
rect 21640 12928 21692 12980
rect 15292 12792 15344 12844
rect 17040 12724 17092 12776
rect 17316 12724 17368 12776
rect 17684 12835 17736 12844
rect 17684 12801 17693 12835
rect 17693 12801 17727 12835
rect 17727 12801 17736 12835
rect 17684 12792 17736 12801
rect 17776 12835 17828 12844
rect 17776 12801 17785 12835
rect 17785 12801 17819 12835
rect 17819 12801 17828 12835
rect 17776 12792 17828 12801
rect 17960 12835 18012 12844
rect 17960 12801 17969 12835
rect 17969 12801 18003 12835
rect 18003 12801 18012 12835
rect 17960 12792 18012 12801
rect 18052 12835 18104 12844
rect 18052 12801 18061 12835
rect 18061 12801 18095 12835
rect 18095 12801 18104 12835
rect 18052 12792 18104 12801
rect 18512 12835 18564 12844
rect 18512 12801 18521 12835
rect 18521 12801 18555 12835
rect 18555 12801 18564 12835
rect 18512 12792 18564 12801
rect 18696 12767 18748 12776
rect 18696 12733 18705 12767
rect 18705 12733 18739 12767
rect 18739 12733 18748 12767
rect 18696 12724 18748 12733
rect 18880 12860 18932 12912
rect 18972 12835 19024 12844
rect 18972 12801 18981 12835
rect 18981 12801 19015 12835
rect 19015 12801 19024 12835
rect 18972 12792 19024 12801
rect 20076 12792 20128 12844
rect 21364 12792 21416 12844
rect 22100 12835 22152 12844
rect 22100 12801 22109 12835
rect 22109 12801 22143 12835
rect 22143 12801 22152 12835
rect 22100 12792 22152 12801
rect 22928 12928 22980 12980
rect 23204 12928 23256 12980
rect 22376 12835 22428 12844
rect 22376 12801 22385 12835
rect 22385 12801 22419 12835
rect 22419 12801 22428 12835
rect 22376 12792 22428 12801
rect 22744 12792 22796 12844
rect 22928 12792 22980 12844
rect 23480 12792 23532 12844
rect 23848 12835 23900 12844
rect 23848 12801 23857 12835
rect 23857 12801 23891 12835
rect 23891 12801 23900 12835
rect 23848 12792 23900 12801
rect 23940 12835 23992 12844
rect 23940 12801 23949 12835
rect 23949 12801 23983 12835
rect 23983 12801 23992 12835
rect 23940 12792 23992 12801
rect 28908 12971 28960 12980
rect 28908 12937 28917 12971
rect 28917 12937 28951 12971
rect 28951 12937 28960 12971
rect 28908 12928 28960 12937
rect 29092 12971 29144 12980
rect 29092 12937 29101 12971
rect 29101 12937 29135 12971
rect 29135 12937 29144 12971
rect 29092 12928 29144 12937
rect 29736 12928 29788 12980
rect 30104 12928 30156 12980
rect 32956 12928 33008 12980
rect 38384 12928 38436 12980
rect 38660 12928 38712 12980
rect 24584 12835 24636 12844
rect 24584 12801 24593 12835
rect 24593 12801 24627 12835
rect 24627 12801 24636 12835
rect 24584 12792 24636 12801
rect 24860 12792 24912 12844
rect 25964 12860 26016 12912
rect 26516 12860 26568 12912
rect 26792 12860 26844 12912
rect 25596 12835 25648 12844
rect 25596 12801 25605 12835
rect 25605 12801 25639 12835
rect 25639 12801 25648 12835
rect 25596 12792 25648 12801
rect 22192 12724 22244 12776
rect 25228 12724 25280 12776
rect 27252 12835 27304 12844
rect 27252 12801 27261 12835
rect 27261 12801 27295 12835
rect 27295 12801 27304 12835
rect 27252 12792 27304 12801
rect 27528 12835 27580 12844
rect 27528 12801 27537 12835
rect 27537 12801 27571 12835
rect 27571 12801 27580 12835
rect 27528 12792 27580 12801
rect 27712 12792 27764 12844
rect 27896 12724 27948 12776
rect 5816 12588 5868 12597
rect 6184 12588 6236 12640
rect 6368 12588 6420 12640
rect 8024 12588 8076 12640
rect 8116 12631 8168 12640
rect 8116 12597 8125 12631
rect 8125 12597 8159 12631
rect 8159 12597 8168 12631
rect 8116 12588 8168 12597
rect 11612 12588 11664 12640
rect 12348 12588 12400 12640
rect 13268 12588 13320 12640
rect 14096 12631 14148 12640
rect 14096 12597 14105 12631
rect 14105 12597 14139 12631
rect 14139 12597 14148 12631
rect 14096 12588 14148 12597
rect 15200 12656 15252 12708
rect 16672 12631 16724 12640
rect 16672 12597 16681 12631
rect 16681 12597 16715 12631
rect 16715 12597 16724 12631
rect 16672 12588 16724 12597
rect 17408 12656 17460 12708
rect 17960 12656 18012 12708
rect 17224 12631 17276 12640
rect 17224 12597 17233 12631
rect 17233 12597 17267 12631
rect 17267 12597 17276 12631
rect 17224 12588 17276 12597
rect 18328 12631 18380 12640
rect 18328 12597 18337 12631
rect 18337 12597 18371 12631
rect 18371 12597 18380 12631
rect 18328 12588 18380 12597
rect 19800 12588 19852 12640
rect 21548 12588 21600 12640
rect 21732 12588 21784 12640
rect 23388 12656 23440 12708
rect 23848 12588 23900 12640
rect 27528 12656 27580 12708
rect 29276 12860 29328 12912
rect 28080 12835 28132 12844
rect 28080 12801 28089 12835
rect 28089 12801 28123 12835
rect 28123 12801 28132 12835
rect 28080 12792 28132 12801
rect 28080 12656 28132 12708
rect 28264 12792 28316 12844
rect 28356 12835 28408 12844
rect 28356 12801 28365 12835
rect 28365 12801 28399 12835
rect 28399 12801 28408 12835
rect 28356 12792 28408 12801
rect 28724 12835 28776 12844
rect 28724 12801 28733 12835
rect 28733 12801 28767 12835
rect 28767 12801 28776 12835
rect 28724 12792 28776 12801
rect 28816 12792 28868 12844
rect 29184 12835 29236 12844
rect 29184 12801 29193 12835
rect 29193 12801 29227 12835
rect 29227 12801 29236 12835
rect 29184 12792 29236 12801
rect 29920 12860 29972 12912
rect 30104 12792 30156 12844
rect 30472 12835 30524 12844
rect 30472 12801 30481 12835
rect 30481 12801 30515 12835
rect 30515 12801 30524 12835
rect 30472 12792 30524 12801
rect 30932 12860 30984 12912
rect 29736 12767 29788 12776
rect 29736 12733 29745 12767
rect 29745 12733 29779 12767
rect 29779 12733 29788 12767
rect 29736 12724 29788 12733
rect 30288 12724 30340 12776
rect 30840 12835 30892 12844
rect 30840 12801 30849 12835
rect 30849 12801 30883 12835
rect 30883 12801 30892 12835
rect 30840 12792 30892 12801
rect 31392 12860 31444 12912
rect 35348 12860 35400 12912
rect 35532 12860 35584 12912
rect 31760 12792 31812 12844
rect 31852 12792 31904 12844
rect 32220 12792 32272 12844
rect 28264 12699 28316 12708
rect 28264 12665 28273 12699
rect 28273 12665 28307 12699
rect 28307 12665 28316 12699
rect 28264 12656 28316 12665
rect 28356 12656 28408 12708
rect 24492 12588 24544 12640
rect 24860 12631 24912 12640
rect 24860 12597 24869 12631
rect 24869 12597 24903 12631
rect 24903 12597 24912 12631
rect 24860 12588 24912 12597
rect 25320 12588 25372 12640
rect 25872 12588 25924 12640
rect 27804 12588 27856 12640
rect 27988 12588 28040 12640
rect 28816 12588 28868 12640
rect 30012 12656 30064 12708
rect 31208 12656 31260 12708
rect 32496 12835 32548 12844
rect 32496 12801 32505 12835
rect 32505 12801 32539 12835
rect 32539 12801 32548 12835
rect 32496 12792 32548 12801
rect 32956 12792 33008 12844
rect 33232 12792 33284 12844
rect 34796 12835 34848 12844
rect 34796 12801 34805 12835
rect 34805 12801 34839 12835
rect 34839 12801 34848 12835
rect 34796 12792 34848 12801
rect 33508 12724 33560 12776
rect 34612 12724 34664 12776
rect 38660 12835 38712 12844
rect 38660 12801 38669 12835
rect 38669 12801 38703 12835
rect 38703 12801 38712 12835
rect 38660 12792 38712 12801
rect 36084 12724 36136 12776
rect 38568 12724 38620 12776
rect 29092 12588 29144 12640
rect 30380 12588 30432 12640
rect 30472 12588 30524 12640
rect 39488 12656 39540 12708
rect 39120 12631 39172 12640
rect 39120 12597 39129 12631
rect 39129 12597 39163 12631
rect 39163 12597 39172 12631
rect 39120 12588 39172 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 4712 12384 4764 12436
rect 4620 12316 4672 12368
rect 4712 12248 4764 12300
rect 5448 12384 5500 12436
rect 6368 12427 6420 12436
rect 6368 12393 6377 12427
rect 6377 12393 6411 12427
rect 6411 12393 6420 12427
rect 6368 12384 6420 12393
rect 6460 12384 6512 12436
rect 3976 12223 4028 12232
rect 3976 12189 3985 12223
rect 3985 12189 4019 12223
rect 4019 12189 4028 12223
rect 3976 12180 4028 12189
rect 5908 12316 5960 12368
rect 6276 12316 6328 12368
rect 5540 12248 5592 12300
rect 6092 12291 6144 12300
rect 6092 12257 6101 12291
rect 6101 12257 6135 12291
rect 6135 12257 6144 12291
rect 6092 12248 6144 12257
rect 7840 12384 7892 12436
rect 13084 12384 13136 12436
rect 17960 12427 18012 12436
rect 17960 12393 17969 12427
rect 17969 12393 18003 12427
rect 18003 12393 18012 12427
rect 17960 12384 18012 12393
rect 17040 12316 17092 12368
rect 18236 12316 18288 12368
rect 18972 12384 19024 12436
rect 19248 12384 19300 12436
rect 19340 12427 19392 12436
rect 19340 12393 19349 12427
rect 19349 12393 19383 12427
rect 19383 12393 19392 12427
rect 19340 12384 19392 12393
rect 19524 12427 19576 12436
rect 19524 12393 19533 12427
rect 19533 12393 19567 12427
rect 19567 12393 19576 12427
rect 19524 12384 19576 12393
rect 19708 12384 19760 12436
rect 19892 12384 19944 12436
rect 20352 12384 20404 12436
rect 21272 12384 21324 12436
rect 21732 12384 21784 12436
rect 18696 12316 18748 12368
rect 23388 12316 23440 12368
rect 23848 12316 23900 12368
rect 7012 12248 7064 12300
rect 7288 12248 7340 12300
rect 14556 12248 14608 12300
rect 5724 12155 5776 12164
rect 5724 12121 5733 12155
rect 5733 12121 5767 12155
rect 5767 12121 5776 12155
rect 5724 12112 5776 12121
rect 3792 12044 3844 12096
rect 5908 12155 5960 12164
rect 5908 12121 5943 12155
rect 5943 12121 5960 12155
rect 6184 12223 6236 12232
rect 6184 12189 6193 12223
rect 6193 12189 6227 12223
rect 6227 12189 6236 12223
rect 6184 12180 6236 12189
rect 6644 12223 6696 12232
rect 6644 12189 6653 12223
rect 6653 12189 6687 12223
rect 6687 12189 6696 12223
rect 6644 12180 6696 12189
rect 6736 12180 6788 12232
rect 7564 12223 7616 12232
rect 7564 12189 7573 12223
rect 7573 12189 7607 12223
rect 7607 12189 7616 12223
rect 7564 12180 7616 12189
rect 7748 12223 7800 12232
rect 7748 12189 7757 12223
rect 7757 12189 7791 12223
rect 7791 12189 7800 12223
rect 7748 12180 7800 12189
rect 12624 12180 12676 12232
rect 12900 12223 12952 12232
rect 12900 12189 12910 12223
rect 12910 12189 12944 12223
rect 12944 12189 12952 12223
rect 12900 12180 12952 12189
rect 13912 12180 13964 12232
rect 15200 12223 15252 12232
rect 15200 12189 15209 12223
rect 15209 12189 15243 12223
rect 15243 12189 15252 12223
rect 15200 12180 15252 12189
rect 17316 12180 17368 12232
rect 19432 12248 19484 12300
rect 20168 12248 20220 12300
rect 28080 12316 28132 12368
rect 29460 12384 29512 12436
rect 30932 12384 30984 12436
rect 33784 12384 33836 12436
rect 34796 12384 34848 12436
rect 37188 12384 37240 12436
rect 38660 12384 38712 12436
rect 33876 12316 33928 12368
rect 5908 12112 5960 12121
rect 8116 12112 8168 12164
rect 10508 12112 10560 12164
rect 15108 12155 15160 12164
rect 15108 12121 15117 12155
rect 15117 12121 15151 12155
rect 15151 12121 15160 12155
rect 15108 12112 15160 12121
rect 18512 12180 18564 12232
rect 18880 12180 18932 12232
rect 18972 12223 19024 12232
rect 18972 12189 18981 12223
rect 18981 12189 19015 12223
rect 19015 12189 19024 12223
rect 18972 12180 19024 12189
rect 19340 12112 19392 12164
rect 19800 12180 19852 12232
rect 20536 12223 20588 12232
rect 20536 12189 20545 12223
rect 20545 12189 20579 12223
rect 20579 12189 20588 12223
rect 20536 12180 20588 12189
rect 22376 12180 22428 12232
rect 22928 12180 22980 12232
rect 26056 12223 26108 12232
rect 26056 12189 26065 12223
rect 26065 12189 26099 12223
rect 26099 12189 26108 12223
rect 30012 12248 30064 12300
rect 26056 12180 26108 12189
rect 26332 12180 26384 12232
rect 27896 12223 27948 12232
rect 27896 12189 27905 12223
rect 27905 12189 27939 12223
rect 27939 12189 27948 12223
rect 27896 12180 27948 12189
rect 7472 12087 7524 12096
rect 7472 12053 7481 12087
rect 7481 12053 7515 12087
rect 7515 12053 7524 12087
rect 7472 12044 7524 12053
rect 8576 12044 8628 12096
rect 9496 12044 9548 12096
rect 12808 12044 12860 12096
rect 14832 12044 14884 12096
rect 15200 12044 15252 12096
rect 18604 12044 18656 12096
rect 19156 12044 19208 12096
rect 20720 12044 20772 12096
rect 20996 12112 21048 12164
rect 26424 12112 26476 12164
rect 28540 12180 28592 12232
rect 29920 12223 29972 12232
rect 29920 12189 29929 12223
rect 29929 12189 29963 12223
rect 29963 12189 29972 12223
rect 29920 12180 29972 12189
rect 30104 12223 30156 12232
rect 30104 12189 30113 12223
rect 30113 12189 30147 12223
rect 30147 12189 30156 12223
rect 30104 12180 30156 12189
rect 22192 12044 22244 12096
rect 25136 12044 25188 12096
rect 28724 12044 28776 12096
rect 29460 12044 29512 12096
rect 30748 12223 30800 12232
rect 30748 12189 30757 12223
rect 30757 12189 30791 12223
rect 30791 12189 30800 12223
rect 30748 12180 30800 12189
rect 33508 12248 33560 12300
rect 37832 12316 37884 12368
rect 33232 12180 33284 12232
rect 30840 12112 30892 12164
rect 34612 12248 34664 12300
rect 33968 12180 34020 12232
rect 36636 12248 36688 12300
rect 39580 12248 39632 12300
rect 35348 12180 35400 12232
rect 35532 12180 35584 12232
rect 38384 12223 38436 12232
rect 38384 12189 38393 12223
rect 38393 12189 38427 12223
rect 38427 12189 38436 12223
rect 38384 12180 38436 12189
rect 34520 12112 34572 12164
rect 34704 12112 34756 12164
rect 31300 12044 31352 12096
rect 31760 12044 31812 12096
rect 34244 12044 34296 12096
rect 34888 12044 34940 12096
rect 35072 12155 35124 12164
rect 35072 12121 35081 12155
rect 35081 12121 35115 12155
rect 35115 12121 35124 12155
rect 35072 12112 35124 12121
rect 35256 12044 35308 12096
rect 35440 12044 35492 12096
rect 38108 12155 38160 12164
rect 38108 12121 38117 12155
rect 38117 12121 38151 12155
rect 38151 12121 38160 12155
rect 38108 12112 38160 12121
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 4160 11840 4212 11892
rect 4712 11840 4764 11892
rect 5540 11840 5592 11892
rect 5724 11840 5776 11892
rect 6552 11840 6604 11892
rect 10508 11840 10560 11892
rect 3792 11815 3844 11824
rect 3792 11781 3801 11815
rect 3801 11781 3835 11815
rect 3835 11781 3844 11815
rect 3792 11772 3844 11781
rect 7656 11772 7708 11824
rect 3240 11636 3292 11688
rect 3516 11679 3568 11688
rect 3516 11645 3525 11679
rect 3525 11645 3559 11679
rect 3559 11645 3568 11679
rect 3516 11636 3568 11645
rect 6736 11747 6788 11756
rect 6736 11713 6745 11747
rect 6745 11713 6779 11747
rect 6779 11713 6788 11747
rect 6736 11704 6788 11713
rect 8300 11704 8352 11756
rect 8852 11815 8904 11824
rect 8852 11781 8861 11815
rect 8861 11781 8895 11815
rect 8895 11781 8904 11815
rect 8852 11772 8904 11781
rect 9588 11772 9640 11824
rect 8760 11747 8812 11756
rect 8760 11713 8769 11747
rect 8769 11713 8803 11747
rect 8803 11713 8812 11747
rect 8760 11704 8812 11713
rect 9312 11704 9364 11756
rect 10968 11772 11020 11824
rect 12992 11772 13044 11824
rect 14464 11840 14516 11892
rect 16856 11883 16908 11892
rect 16856 11849 16865 11883
rect 16865 11849 16899 11883
rect 16899 11849 16908 11883
rect 16856 11840 16908 11849
rect 18972 11840 19024 11892
rect 19156 11840 19208 11892
rect 15200 11815 15252 11824
rect 15200 11781 15209 11815
rect 15209 11781 15243 11815
rect 15243 11781 15252 11815
rect 15200 11772 15252 11781
rect 17408 11772 17460 11824
rect 17776 11772 17828 11824
rect 7748 11636 7800 11688
rect 9588 11636 9640 11688
rect 8852 11568 8904 11620
rect 13084 11747 13136 11756
rect 13084 11713 13093 11747
rect 13093 11713 13127 11747
rect 13127 11713 13136 11747
rect 13084 11704 13136 11713
rect 9864 11636 9916 11688
rect 10324 11636 10376 11688
rect 10968 11636 11020 11688
rect 11888 11636 11940 11688
rect 12256 11636 12308 11688
rect 12532 11636 12584 11688
rect 13452 11636 13504 11688
rect 13912 11636 13964 11688
rect 15476 11747 15528 11756
rect 15476 11713 15485 11747
rect 15485 11713 15519 11747
rect 15519 11713 15528 11747
rect 15476 11704 15528 11713
rect 16120 11704 16172 11756
rect 17040 11747 17092 11756
rect 17040 11713 17049 11747
rect 17049 11713 17083 11747
rect 17083 11713 17092 11747
rect 17040 11704 17092 11713
rect 17684 11704 17736 11756
rect 19524 11704 19576 11756
rect 20076 11747 20128 11756
rect 20076 11713 20085 11747
rect 20085 11713 20119 11747
rect 20119 11713 20128 11747
rect 20076 11704 20128 11713
rect 20260 11704 20312 11756
rect 20996 11772 21048 11824
rect 22008 11772 22060 11824
rect 24860 11772 24912 11824
rect 25596 11840 25648 11892
rect 25688 11840 25740 11892
rect 31208 11840 31260 11892
rect 33048 11840 33100 11892
rect 33600 11840 33652 11892
rect 8668 11500 8720 11552
rect 9588 11500 9640 11552
rect 10048 11500 10100 11552
rect 12164 11568 12216 11620
rect 12348 11568 12400 11620
rect 18236 11636 18288 11688
rect 20904 11704 20956 11756
rect 21548 11704 21600 11756
rect 22744 11704 22796 11756
rect 23388 11704 23440 11756
rect 24216 11704 24268 11756
rect 24492 11747 24544 11756
rect 24492 11713 24501 11747
rect 24501 11713 24535 11747
rect 24535 11713 24544 11747
rect 24492 11704 24544 11713
rect 24952 11747 25004 11756
rect 24952 11713 24961 11747
rect 24961 11713 24995 11747
rect 24995 11713 25004 11747
rect 24952 11704 25004 11713
rect 25136 11747 25188 11756
rect 25136 11713 25145 11747
rect 25145 11713 25179 11747
rect 25179 11713 25188 11747
rect 25136 11704 25188 11713
rect 25320 11704 25372 11756
rect 20720 11636 20772 11688
rect 21272 11636 21324 11688
rect 22100 11636 22152 11688
rect 23204 11679 23256 11688
rect 23204 11645 23213 11679
rect 23213 11645 23247 11679
rect 23247 11645 23256 11679
rect 23204 11636 23256 11645
rect 12256 11500 12308 11552
rect 13452 11543 13504 11552
rect 13452 11509 13461 11543
rect 13461 11509 13495 11543
rect 13495 11509 13504 11543
rect 13452 11500 13504 11509
rect 16764 11568 16816 11620
rect 17776 11568 17828 11620
rect 19800 11568 19852 11620
rect 20168 11568 20220 11620
rect 25412 11636 25464 11688
rect 25964 11772 26016 11824
rect 26332 11772 26384 11824
rect 26056 11636 26108 11688
rect 25228 11568 25280 11620
rect 25688 11568 25740 11620
rect 25964 11568 26016 11620
rect 26240 11704 26292 11756
rect 26424 11747 26476 11756
rect 26424 11713 26433 11747
rect 26433 11713 26467 11747
rect 26467 11713 26476 11747
rect 26424 11704 26476 11713
rect 30196 11772 30248 11824
rect 33508 11772 33560 11824
rect 34796 11840 34848 11892
rect 35072 11840 35124 11892
rect 38108 11840 38160 11892
rect 34888 11815 34940 11824
rect 34888 11781 34897 11815
rect 34897 11781 34931 11815
rect 34931 11781 34940 11815
rect 34888 11772 34940 11781
rect 27988 11704 28040 11756
rect 28448 11704 28500 11756
rect 29460 11704 29512 11756
rect 30104 11704 30156 11756
rect 32864 11704 32916 11756
rect 33600 11747 33652 11756
rect 33600 11713 33609 11747
rect 33609 11713 33643 11747
rect 33643 11713 33652 11747
rect 33600 11704 33652 11713
rect 34060 11704 34112 11756
rect 35348 11704 35400 11756
rect 36268 11704 36320 11756
rect 36544 11747 36596 11756
rect 36544 11713 36554 11747
rect 36554 11713 36588 11747
rect 36588 11713 36596 11747
rect 36544 11704 36596 11713
rect 36636 11704 36688 11756
rect 36820 11747 36872 11756
rect 36820 11713 36829 11747
rect 36829 11713 36863 11747
rect 36863 11713 36872 11747
rect 36820 11704 36872 11713
rect 29552 11636 29604 11688
rect 30564 11636 30616 11688
rect 31852 11636 31904 11688
rect 33508 11636 33560 11688
rect 38016 11747 38068 11756
rect 38016 11713 38025 11747
rect 38025 11713 38059 11747
rect 38059 11713 38068 11747
rect 38016 11704 38068 11713
rect 38292 11747 38344 11756
rect 38292 11713 38301 11747
rect 38301 11713 38335 11747
rect 38335 11713 38344 11747
rect 38292 11704 38344 11713
rect 38752 11747 38804 11756
rect 38752 11713 38761 11747
rect 38761 11713 38795 11747
rect 38795 11713 38804 11747
rect 38752 11704 38804 11713
rect 26516 11568 26568 11620
rect 26884 11568 26936 11620
rect 20076 11500 20128 11552
rect 20444 11500 20496 11552
rect 21364 11500 21416 11552
rect 24768 11543 24820 11552
rect 24768 11509 24777 11543
rect 24777 11509 24811 11543
rect 24811 11509 24820 11543
rect 24768 11500 24820 11509
rect 24952 11500 25004 11552
rect 25872 11543 25924 11552
rect 25872 11509 25881 11543
rect 25881 11509 25915 11543
rect 25915 11509 25924 11543
rect 25872 11500 25924 11509
rect 26240 11500 26292 11552
rect 27620 11500 27672 11552
rect 28356 11500 28408 11552
rect 28632 11543 28684 11552
rect 28632 11509 28641 11543
rect 28641 11509 28675 11543
rect 28675 11509 28684 11543
rect 28632 11500 28684 11509
rect 31944 11500 31996 11552
rect 33416 11500 33468 11552
rect 37372 11636 37424 11688
rect 38936 11679 38988 11688
rect 38936 11645 38945 11679
rect 38945 11645 38979 11679
rect 38979 11645 38988 11679
rect 38936 11636 38988 11645
rect 34612 11500 34664 11552
rect 38384 11500 38436 11552
rect 38568 11543 38620 11552
rect 38568 11509 38577 11543
rect 38577 11509 38611 11543
rect 38611 11509 38620 11543
rect 38568 11500 38620 11509
rect 39304 11500 39356 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 8668 11339 8720 11348
rect 8668 11305 8677 11339
rect 8677 11305 8711 11339
rect 8711 11305 8720 11339
rect 8668 11296 8720 11305
rect 9312 11296 9364 11348
rect 7104 11228 7156 11280
rect 9588 11160 9640 11212
rect 3516 11092 3568 11144
rect 7656 11092 7708 11144
rect 8392 11092 8444 11144
rect 7932 11067 7984 11076
rect 7932 11033 7941 11067
rect 7941 11033 7975 11067
rect 7975 11033 7984 11067
rect 7932 11024 7984 11033
rect 8208 11024 8260 11076
rect 9312 11092 9364 11144
rect 9496 11092 9548 11144
rect 9404 11024 9456 11076
rect 9956 11092 10008 11144
rect 10048 11135 10100 11144
rect 10048 11101 10057 11135
rect 10057 11101 10091 11135
rect 10091 11101 10100 11135
rect 10048 11092 10100 11101
rect 12164 11296 12216 11348
rect 12348 11296 12400 11348
rect 10324 11024 10376 11076
rect 10876 11135 10928 11144
rect 10876 11101 10885 11135
rect 10885 11101 10919 11135
rect 10919 11101 10928 11135
rect 10876 11092 10928 11101
rect 11152 11135 11204 11144
rect 11152 11101 11161 11135
rect 11161 11101 11195 11135
rect 11195 11101 11204 11135
rect 11152 11092 11204 11101
rect 11428 11092 11480 11144
rect 12440 11228 12492 11280
rect 12532 11135 12584 11144
rect 12532 11101 12541 11135
rect 12541 11101 12575 11135
rect 12575 11101 12584 11135
rect 12532 11092 12584 11101
rect 13820 11296 13872 11348
rect 15108 11296 15160 11348
rect 17316 11339 17368 11348
rect 17316 11305 17325 11339
rect 17325 11305 17359 11339
rect 17359 11305 17368 11339
rect 17316 11296 17368 11305
rect 17868 11296 17920 11348
rect 18236 11339 18288 11348
rect 18236 11305 18245 11339
rect 18245 11305 18279 11339
rect 18279 11305 18288 11339
rect 18236 11296 18288 11305
rect 19248 11296 19300 11348
rect 20996 11296 21048 11348
rect 21088 11296 21140 11348
rect 21272 11296 21324 11348
rect 22192 11296 22244 11348
rect 22468 11296 22520 11348
rect 24400 11339 24452 11348
rect 24400 11305 24409 11339
rect 24409 11305 24443 11339
rect 24443 11305 24452 11339
rect 24400 11296 24452 11305
rect 12808 11228 12860 11280
rect 15200 11160 15252 11212
rect 16120 11160 16172 11212
rect 17592 11160 17644 11212
rect 20536 11228 20588 11280
rect 24768 11296 24820 11348
rect 26056 11296 26108 11348
rect 26792 11296 26844 11348
rect 27988 11339 28040 11348
rect 27988 11305 27997 11339
rect 27997 11305 28031 11339
rect 28031 11305 28040 11339
rect 27988 11296 28040 11305
rect 28264 11296 28316 11348
rect 29552 11339 29604 11348
rect 29552 11305 29561 11339
rect 29561 11305 29595 11339
rect 29595 11305 29604 11339
rect 29552 11296 29604 11305
rect 30932 11296 30984 11348
rect 37280 11296 37332 11348
rect 12256 11024 12308 11076
rect 1860 10999 1912 11008
rect 1860 10965 1869 10999
rect 1869 10965 1903 10999
rect 1903 10965 1912 10999
rect 1860 10956 1912 10965
rect 8300 10999 8352 11008
rect 8300 10965 8309 10999
rect 8309 10965 8343 10999
rect 8343 10965 8352 10999
rect 8300 10956 8352 10965
rect 9496 10956 9548 11008
rect 9772 10956 9824 11008
rect 10692 10956 10744 11008
rect 12348 10956 12400 11008
rect 13452 11092 13504 11144
rect 14372 11092 14424 11144
rect 16580 11092 16632 11144
rect 16948 11092 17000 11144
rect 17776 11135 17828 11144
rect 17776 11101 17785 11135
rect 17785 11101 17819 11135
rect 17819 11101 17828 11135
rect 17776 11092 17828 11101
rect 20352 11203 20404 11212
rect 20352 11169 20361 11203
rect 20361 11169 20395 11203
rect 20395 11169 20404 11203
rect 20352 11160 20404 11169
rect 20812 11160 20864 11212
rect 18512 11135 18564 11144
rect 18512 11101 18521 11135
rect 18521 11101 18555 11135
rect 18555 11101 18564 11135
rect 18512 11092 18564 11101
rect 17408 10956 17460 11008
rect 19340 11024 19392 11076
rect 19708 11067 19760 11076
rect 19708 11033 19717 11067
rect 19717 11033 19751 11067
rect 19751 11033 19760 11067
rect 19708 11024 19760 11033
rect 20260 11024 20312 11076
rect 21456 11024 21508 11076
rect 22284 11203 22336 11212
rect 22284 11169 22293 11203
rect 22293 11169 22327 11203
rect 22327 11169 22336 11203
rect 22284 11160 22336 11169
rect 22468 11135 22520 11144
rect 22468 11101 22477 11135
rect 22477 11101 22511 11135
rect 22511 11101 22520 11135
rect 22468 11092 22520 11101
rect 25412 11228 25464 11280
rect 27988 11160 28040 11212
rect 23204 11135 23256 11144
rect 23204 11101 23213 11135
rect 23213 11101 23247 11135
rect 23247 11101 23256 11135
rect 23204 11092 23256 11101
rect 24768 11135 24820 11144
rect 24768 11101 24777 11135
rect 24777 11101 24811 11135
rect 24811 11101 24820 11135
rect 24768 11092 24820 11101
rect 25136 11092 25188 11144
rect 26332 11092 26384 11144
rect 26792 11135 26844 11144
rect 26792 11101 26801 11135
rect 26801 11101 26835 11135
rect 26835 11101 26844 11135
rect 26792 11092 26844 11101
rect 26976 11092 27028 11144
rect 26424 11024 26476 11076
rect 20720 10956 20772 11008
rect 21916 10999 21968 11008
rect 21916 10965 21925 10999
rect 21925 10965 21959 10999
rect 21959 10965 21968 10999
rect 21916 10956 21968 10965
rect 23020 10956 23072 11008
rect 27712 11092 27764 11144
rect 27896 11135 27948 11144
rect 27896 11101 27905 11135
rect 27905 11101 27939 11135
rect 27939 11101 27948 11135
rect 27896 11092 27948 11101
rect 28356 11092 28408 11144
rect 28816 11092 28868 11144
rect 29184 11135 29236 11144
rect 29184 11101 29193 11135
rect 29193 11101 29227 11135
rect 29227 11101 29236 11135
rect 29184 11092 29236 11101
rect 29460 11092 29512 11144
rect 30196 11160 30248 11212
rect 32220 11160 32272 11212
rect 33048 11160 33100 11212
rect 33968 11228 34020 11280
rect 33324 11203 33376 11212
rect 33324 11169 33333 11203
rect 33333 11169 33367 11203
rect 33367 11169 33376 11203
rect 33324 11160 33376 11169
rect 33600 11160 33652 11212
rect 28540 10956 28592 11008
rect 29092 10956 29144 11008
rect 29460 10956 29512 11008
rect 29828 10956 29880 11008
rect 30012 11024 30064 11076
rect 30288 11067 30340 11076
rect 30288 11033 30297 11067
rect 30297 11033 30331 11067
rect 30331 11033 30340 11067
rect 30288 11024 30340 11033
rect 30564 11135 30616 11144
rect 30564 11101 30573 11135
rect 30573 11101 30607 11135
rect 30607 11101 30616 11135
rect 30564 11092 30616 11101
rect 30840 11092 30892 11144
rect 30748 11024 30800 11076
rect 30472 10956 30524 11008
rect 31116 10956 31168 11008
rect 31668 11024 31720 11076
rect 32864 11135 32916 11144
rect 32864 11101 32873 11135
rect 32873 11101 32907 11135
rect 32907 11101 32916 11135
rect 32864 11092 32916 11101
rect 33416 11135 33468 11144
rect 33416 11101 33425 11135
rect 33425 11101 33459 11135
rect 33459 11101 33468 11135
rect 33416 11092 33468 11101
rect 33876 11135 33928 11144
rect 33876 11101 33893 11135
rect 33893 11101 33928 11135
rect 33324 11024 33376 11076
rect 33876 11092 33928 11101
rect 32128 10956 32180 11008
rect 32680 10956 32732 11008
rect 32772 10956 32824 11008
rect 33968 11067 34020 11076
rect 33968 11033 33977 11067
rect 33977 11033 34011 11067
rect 34011 11033 34020 11067
rect 33968 11024 34020 11033
rect 34336 11135 34388 11144
rect 34336 11101 34345 11135
rect 34345 11101 34379 11135
rect 34379 11101 34388 11135
rect 34336 11092 34388 11101
rect 34612 11092 34664 11144
rect 35348 11160 35400 11212
rect 34980 11135 35032 11144
rect 34980 11101 34989 11135
rect 34989 11101 35023 11135
rect 35023 11101 35032 11135
rect 34980 11092 35032 11101
rect 35992 11092 36044 11144
rect 36084 11024 36136 11076
rect 34612 10956 34664 11008
rect 34704 10999 34756 11008
rect 34704 10965 34713 10999
rect 34713 10965 34747 10999
rect 34747 10965 34756 10999
rect 34704 10956 34756 10965
rect 34888 10956 34940 11008
rect 38476 11228 38528 11280
rect 37096 11203 37148 11212
rect 37096 11169 37105 11203
rect 37105 11169 37139 11203
rect 37139 11169 37148 11203
rect 37096 11160 37148 11169
rect 36636 11135 36688 11144
rect 36636 11101 36645 11135
rect 36645 11101 36679 11135
rect 36679 11101 36688 11135
rect 36636 11092 36688 11101
rect 36728 11135 36780 11144
rect 36728 11101 36737 11135
rect 36737 11101 36771 11135
rect 36771 11101 36780 11135
rect 36728 11092 36780 11101
rect 39672 11160 39724 11212
rect 37280 11135 37332 11144
rect 37280 11101 37289 11135
rect 37289 11101 37323 11135
rect 37323 11101 37332 11135
rect 37280 11092 37332 11101
rect 38292 10956 38344 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 7380 10795 7432 10804
rect 7380 10761 7389 10795
rect 7389 10761 7423 10795
rect 7423 10761 7432 10795
rect 7380 10752 7432 10761
rect 5724 10684 5776 10736
rect 7656 10684 7708 10736
rect 6552 10659 6604 10668
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 6736 10659 6788 10668
rect 6736 10625 6745 10659
rect 6745 10625 6779 10659
rect 6779 10625 6788 10659
rect 6736 10616 6788 10625
rect 6920 10659 6972 10668
rect 6920 10625 6929 10659
rect 6929 10625 6963 10659
rect 6963 10625 6972 10659
rect 6920 10616 6972 10625
rect 7472 10659 7524 10668
rect 7472 10625 7481 10659
rect 7481 10625 7515 10659
rect 7515 10625 7524 10659
rect 7472 10616 7524 10625
rect 7932 10616 7984 10668
rect 8392 10727 8444 10736
rect 8392 10693 8401 10727
rect 8401 10693 8435 10727
rect 8435 10693 8444 10727
rect 8392 10684 8444 10693
rect 8208 10659 8260 10668
rect 8208 10625 8217 10659
rect 8217 10625 8251 10659
rect 8251 10625 8260 10659
rect 8208 10616 8260 10625
rect 8760 10684 8812 10736
rect 10048 10752 10100 10804
rect 10416 10752 10468 10804
rect 16948 10795 17000 10804
rect 16948 10761 16957 10795
rect 16957 10761 16991 10795
rect 16991 10761 17000 10795
rect 16948 10752 17000 10761
rect 9864 10659 9916 10668
rect 9864 10625 9872 10659
rect 9872 10625 9906 10659
rect 9906 10625 9916 10659
rect 9864 10616 9916 10625
rect 10876 10684 10928 10736
rect 12348 10684 12400 10736
rect 14740 10684 14792 10736
rect 6368 10455 6420 10464
rect 6368 10421 6377 10455
rect 6377 10421 6411 10455
rect 6411 10421 6420 10455
rect 6368 10412 6420 10421
rect 7012 10455 7064 10464
rect 7012 10421 7021 10455
rect 7021 10421 7055 10455
rect 7055 10421 7064 10455
rect 7012 10412 7064 10421
rect 7380 10412 7432 10464
rect 9772 10548 9824 10600
rect 10140 10616 10192 10668
rect 9312 10480 9364 10532
rect 11888 10616 11940 10668
rect 12440 10659 12492 10668
rect 12440 10625 12449 10659
rect 12449 10625 12483 10659
rect 12483 10625 12492 10659
rect 12440 10616 12492 10625
rect 12624 10659 12676 10668
rect 12624 10625 12633 10659
rect 12633 10625 12667 10659
rect 12667 10625 12676 10659
rect 12624 10616 12676 10625
rect 12992 10616 13044 10668
rect 14464 10616 14516 10668
rect 15384 10616 15436 10668
rect 21088 10684 21140 10736
rect 20812 10616 20864 10668
rect 20996 10659 21048 10668
rect 20996 10625 21005 10659
rect 21005 10625 21039 10659
rect 21039 10625 21048 10659
rect 20996 10616 21048 10625
rect 21824 10752 21876 10804
rect 22468 10752 22520 10804
rect 23112 10795 23164 10804
rect 23112 10761 23121 10795
rect 23121 10761 23155 10795
rect 23155 10761 23164 10795
rect 23112 10752 23164 10761
rect 24032 10795 24084 10804
rect 24032 10761 24041 10795
rect 24041 10761 24075 10795
rect 24075 10761 24084 10795
rect 24032 10752 24084 10761
rect 22100 10684 22152 10736
rect 25228 10752 25280 10804
rect 24308 10684 24360 10736
rect 24492 10684 24544 10736
rect 21272 10659 21324 10668
rect 21272 10625 21281 10659
rect 21281 10625 21315 10659
rect 21315 10625 21324 10659
rect 21272 10616 21324 10625
rect 21548 10616 21600 10668
rect 21824 10659 21876 10668
rect 21824 10625 21833 10659
rect 21833 10625 21867 10659
rect 21867 10625 21876 10659
rect 21824 10616 21876 10625
rect 22468 10616 22520 10668
rect 23020 10659 23072 10668
rect 23020 10625 23029 10659
rect 23029 10625 23063 10659
rect 23063 10625 23072 10659
rect 23020 10616 23072 10625
rect 23388 10616 23440 10668
rect 24768 10616 24820 10668
rect 15200 10548 15252 10600
rect 21732 10548 21784 10600
rect 21916 10548 21968 10600
rect 24860 10548 24912 10600
rect 25412 10727 25464 10736
rect 25412 10693 25421 10727
rect 25421 10693 25455 10727
rect 25455 10693 25464 10727
rect 25412 10684 25464 10693
rect 25320 10616 25372 10668
rect 26056 10795 26108 10804
rect 26056 10761 26065 10795
rect 26065 10761 26099 10795
rect 26099 10761 26108 10795
rect 26056 10752 26108 10761
rect 27804 10752 27856 10804
rect 27896 10752 27948 10804
rect 28356 10752 28408 10804
rect 31208 10795 31260 10804
rect 31208 10761 31217 10795
rect 31217 10761 31251 10795
rect 31251 10761 31260 10795
rect 31208 10752 31260 10761
rect 26424 10684 26476 10736
rect 26056 10616 26108 10668
rect 27620 10616 27672 10668
rect 28540 10684 28592 10736
rect 29644 10727 29696 10736
rect 29644 10693 29653 10727
rect 29653 10693 29687 10727
rect 29687 10693 29696 10727
rect 29644 10684 29696 10693
rect 32864 10795 32916 10804
rect 32864 10761 32873 10795
rect 32873 10761 32907 10795
rect 32907 10761 32916 10795
rect 32864 10752 32916 10761
rect 27988 10616 28040 10668
rect 28264 10616 28316 10668
rect 28816 10616 28868 10668
rect 29184 10616 29236 10668
rect 29828 10659 29880 10668
rect 29828 10625 29837 10659
rect 29837 10625 29871 10659
rect 29871 10625 29880 10659
rect 29828 10616 29880 10625
rect 30288 10659 30340 10668
rect 30288 10625 30297 10659
rect 30297 10625 30331 10659
rect 30331 10625 30340 10659
rect 30288 10616 30340 10625
rect 30840 10659 30892 10668
rect 30840 10625 30849 10659
rect 30849 10625 30883 10659
rect 30883 10625 30892 10659
rect 30840 10616 30892 10625
rect 32220 10684 32272 10736
rect 33968 10684 34020 10736
rect 34336 10684 34388 10736
rect 37556 10752 37608 10804
rect 39120 10684 39172 10736
rect 31116 10616 31168 10668
rect 11888 10480 11940 10532
rect 18696 10480 18748 10532
rect 24124 10480 24176 10532
rect 8116 10455 8168 10464
rect 8116 10421 8125 10455
rect 8125 10421 8159 10455
rect 8159 10421 8168 10455
rect 8116 10412 8168 10421
rect 8484 10412 8536 10464
rect 8760 10455 8812 10464
rect 8760 10421 8769 10455
rect 8769 10421 8803 10455
rect 8803 10421 8812 10455
rect 8760 10412 8812 10421
rect 10232 10412 10284 10464
rect 13452 10412 13504 10464
rect 14740 10455 14792 10464
rect 14740 10421 14749 10455
rect 14749 10421 14783 10455
rect 14783 10421 14792 10455
rect 14740 10412 14792 10421
rect 15016 10412 15068 10464
rect 17040 10412 17092 10464
rect 19524 10412 19576 10464
rect 20352 10412 20404 10464
rect 20996 10412 21048 10464
rect 21824 10412 21876 10464
rect 22008 10412 22060 10464
rect 22376 10412 22428 10464
rect 25044 10412 25096 10464
rect 28080 10480 28132 10532
rect 31392 10480 31444 10532
rect 31852 10616 31904 10668
rect 32312 10659 32364 10668
rect 32312 10625 32321 10659
rect 32321 10625 32355 10659
rect 32355 10625 32364 10659
rect 32312 10616 32364 10625
rect 32588 10616 32640 10668
rect 32864 10616 32916 10668
rect 32956 10616 33008 10668
rect 34704 10616 34756 10668
rect 37556 10659 37608 10668
rect 37556 10625 37565 10659
rect 37565 10625 37599 10659
rect 37599 10625 37608 10659
rect 37556 10616 37608 10625
rect 38292 10659 38344 10668
rect 38292 10625 38301 10659
rect 38301 10625 38335 10659
rect 38335 10625 38344 10659
rect 38292 10616 38344 10625
rect 39212 10616 39264 10668
rect 32128 10548 32180 10600
rect 31944 10480 31996 10532
rect 33232 10591 33284 10600
rect 33232 10557 33241 10591
rect 33241 10557 33275 10591
rect 33275 10557 33284 10591
rect 33232 10548 33284 10557
rect 37740 10548 37792 10600
rect 34060 10480 34112 10532
rect 36084 10480 36136 10532
rect 31116 10412 31168 10464
rect 34704 10412 34756 10464
rect 35348 10412 35400 10464
rect 38752 10480 38804 10532
rect 38660 10455 38712 10464
rect 38660 10421 38669 10455
rect 38669 10421 38703 10455
rect 38703 10421 38712 10455
rect 38660 10412 38712 10421
rect 39396 10412 39448 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 6368 10208 6420 10260
rect 6736 10208 6788 10260
rect 8668 10208 8720 10260
rect 8760 10208 8812 10260
rect 12624 10251 12676 10260
rect 12624 10217 12633 10251
rect 12633 10217 12667 10251
rect 12667 10217 12676 10251
rect 12624 10208 12676 10217
rect 5724 10183 5776 10192
rect 5724 10149 5733 10183
rect 5733 10149 5767 10183
rect 5767 10149 5776 10183
rect 5724 10140 5776 10149
rect 3516 10072 3568 10124
rect 4712 9936 4764 9988
rect 7104 10047 7156 10056
rect 7104 10013 7113 10047
rect 7113 10013 7147 10047
rect 7147 10013 7156 10047
rect 7104 10004 7156 10013
rect 6828 9979 6880 9988
rect 6828 9945 6837 9979
rect 6837 9945 6871 9979
rect 6871 9945 6880 9979
rect 6828 9936 6880 9945
rect 7380 10047 7432 10056
rect 7380 10013 7389 10047
rect 7389 10013 7423 10047
rect 7423 10013 7432 10047
rect 7380 10004 7432 10013
rect 8116 10072 8168 10124
rect 7564 10047 7616 10056
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 7656 10004 7708 10056
rect 7932 10004 7984 10056
rect 8300 10047 8352 10056
rect 8300 10013 8309 10047
rect 8309 10013 8343 10047
rect 8343 10013 8352 10047
rect 8300 10004 8352 10013
rect 9588 10140 9640 10192
rect 9036 10072 9088 10124
rect 10324 10140 10376 10192
rect 11796 10140 11848 10192
rect 14556 10208 14608 10260
rect 14924 10251 14976 10260
rect 14924 10217 14933 10251
rect 14933 10217 14967 10251
rect 14967 10217 14976 10251
rect 14924 10208 14976 10217
rect 16856 10251 16908 10260
rect 16856 10217 16865 10251
rect 16865 10217 16899 10251
rect 16899 10217 16908 10251
rect 16856 10208 16908 10217
rect 18696 10251 18748 10260
rect 18696 10217 18705 10251
rect 18705 10217 18739 10251
rect 18739 10217 18748 10251
rect 18696 10208 18748 10217
rect 12440 10072 12492 10124
rect 19524 10251 19576 10260
rect 19524 10217 19533 10251
rect 19533 10217 19567 10251
rect 19567 10217 19576 10251
rect 19524 10208 19576 10217
rect 20352 10208 20404 10260
rect 26608 10208 26660 10260
rect 27712 10208 27764 10260
rect 28080 10208 28132 10260
rect 29184 10208 29236 10260
rect 9588 9936 9640 9988
rect 10140 10004 10192 10056
rect 10232 10047 10284 10056
rect 10232 10013 10241 10047
rect 10241 10013 10275 10047
rect 10275 10013 10284 10047
rect 10232 10004 10284 10013
rect 10692 10004 10744 10056
rect 11520 10047 11572 10056
rect 11520 10013 11529 10047
rect 11529 10013 11563 10047
rect 11563 10013 11572 10047
rect 11520 10004 11572 10013
rect 11888 9936 11940 9988
rect 12532 9936 12584 9988
rect 12716 10047 12768 10056
rect 12716 10013 12725 10047
rect 12725 10013 12759 10047
rect 12759 10013 12768 10047
rect 12716 10004 12768 10013
rect 12808 10004 12860 10056
rect 15016 10004 15068 10056
rect 17224 10047 17276 10056
rect 17224 10013 17233 10047
rect 17233 10013 17267 10047
rect 17267 10013 17276 10047
rect 17224 10004 17276 10013
rect 17592 10047 17644 10056
rect 17592 10013 17601 10047
rect 17601 10013 17635 10047
rect 17635 10013 17644 10047
rect 17592 10004 17644 10013
rect 7288 9868 7340 9920
rect 7656 9911 7708 9920
rect 7656 9877 7665 9911
rect 7665 9877 7699 9911
rect 7699 9877 7708 9911
rect 7656 9868 7708 9877
rect 7748 9868 7800 9920
rect 9036 9868 9088 9920
rect 9312 9868 9364 9920
rect 11060 9868 11112 9920
rect 12808 9911 12860 9920
rect 12808 9877 12817 9911
rect 12817 9877 12851 9911
rect 12851 9877 12860 9911
rect 12808 9868 12860 9877
rect 14372 9936 14424 9988
rect 15384 9979 15436 9988
rect 15384 9945 15393 9979
rect 15393 9945 15427 9979
rect 15427 9945 15436 9979
rect 15384 9936 15436 9945
rect 14648 9868 14700 9920
rect 14832 9868 14884 9920
rect 17316 9979 17368 9988
rect 17316 9945 17325 9979
rect 17325 9945 17359 9979
rect 17359 9945 17368 9979
rect 17316 9936 17368 9945
rect 17408 9979 17460 9988
rect 17408 9945 17417 9979
rect 17417 9945 17451 9979
rect 17451 9945 17460 9979
rect 17408 9936 17460 9945
rect 17040 9911 17092 9920
rect 17040 9877 17049 9911
rect 17049 9877 17083 9911
rect 17083 9877 17092 9911
rect 17040 9868 17092 9877
rect 17776 9868 17828 9920
rect 18328 10004 18380 10056
rect 19064 10047 19116 10056
rect 19064 10013 19073 10047
rect 19073 10013 19107 10047
rect 19107 10013 19116 10047
rect 19064 10004 19116 10013
rect 19340 10115 19392 10124
rect 19340 10081 19349 10115
rect 19349 10081 19383 10115
rect 19383 10081 19392 10115
rect 19340 10072 19392 10081
rect 19616 10072 19668 10124
rect 19984 10140 20036 10192
rect 24308 10140 24360 10192
rect 19524 10047 19576 10056
rect 19524 10013 19533 10047
rect 19533 10013 19567 10047
rect 19567 10013 19576 10047
rect 19524 10004 19576 10013
rect 19248 9979 19300 9988
rect 19248 9945 19257 9979
rect 19257 9945 19291 9979
rect 19291 9945 19300 9979
rect 19248 9936 19300 9945
rect 19432 9936 19484 9988
rect 19984 10047 20036 10056
rect 19984 10013 19993 10047
rect 19993 10013 20027 10047
rect 20027 10013 20036 10047
rect 19984 10004 20036 10013
rect 25136 10072 25188 10124
rect 25780 10072 25832 10124
rect 23848 10004 23900 10056
rect 24308 10004 24360 10056
rect 24860 10047 24912 10056
rect 24860 10013 24869 10047
rect 24869 10013 24903 10047
rect 24903 10013 24912 10047
rect 24860 10004 24912 10013
rect 25320 10047 25372 10056
rect 25320 10013 25329 10047
rect 25329 10013 25363 10047
rect 25363 10013 25372 10047
rect 25320 10004 25372 10013
rect 25596 10047 25648 10056
rect 25596 10013 25605 10047
rect 25605 10013 25639 10047
rect 25639 10013 25648 10047
rect 25596 10004 25648 10013
rect 27804 10140 27856 10192
rect 27160 10072 27212 10124
rect 19800 9979 19852 9988
rect 19800 9945 19809 9979
rect 19809 9945 19843 9979
rect 19843 9945 19852 9979
rect 19800 9936 19852 9945
rect 25412 9936 25464 9988
rect 26240 9936 26292 9988
rect 24400 9868 24452 9920
rect 25136 9911 25188 9920
rect 25136 9877 25145 9911
rect 25145 9877 25179 9911
rect 25179 9877 25188 9911
rect 25136 9868 25188 9877
rect 26148 9911 26200 9920
rect 26148 9877 26157 9911
rect 26157 9877 26191 9911
rect 26191 9877 26200 9911
rect 26148 9868 26200 9877
rect 26424 10047 26476 10056
rect 26424 10013 26433 10047
rect 26433 10013 26467 10047
rect 26467 10013 26476 10047
rect 26424 10004 26476 10013
rect 27620 10004 27672 10056
rect 27344 9936 27396 9988
rect 28448 10047 28500 10056
rect 28448 10013 28457 10047
rect 28457 10013 28491 10047
rect 28491 10013 28500 10047
rect 28448 10004 28500 10013
rect 28632 10004 28684 10056
rect 30656 10208 30708 10260
rect 30932 10208 30984 10260
rect 29092 10004 29144 10056
rect 31116 10140 31168 10192
rect 31392 10140 31444 10192
rect 31760 10208 31812 10260
rect 32772 10251 32824 10260
rect 32772 10217 32781 10251
rect 32781 10217 32815 10251
rect 32815 10217 32824 10251
rect 32772 10208 32824 10217
rect 29552 10072 29604 10124
rect 33416 10208 33468 10260
rect 34704 10208 34756 10260
rect 37280 10208 37332 10260
rect 29828 10047 29880 10056
rect 29828 10013 29837 10047
rect 29837 10013 29871 10047
rect 29871 10013 29880 10047
rect 29828 10004 29880 10013
rect 30104 10004 30156 10056
rect 30748 10004 30800 10056
rect 35164 10072 35216 10124
rect 31392 10004 31444 10056
rect 32036 10004 32088 10056
rect 32680 10004 32732 10056
rect 33048 10004 33100 10056
rect 34520 10004 34572 10056
rect 35072 10004 35124 10056
rect 37188 10072 37240 10124
rect 38200 10072 38252 10124
rect 32128 9979 32180 9988
rect 26884 9868 26936 9920
rect 27896 9911 27948 9920
rect 27896 9877 27905 9911
rect 27905 9877 27939 9911
rect 27939 9877 27948 9911
rect 27896 9868 27948 9877
rect 28264 9911 28316 9920
rect 28264 9877 28273 9911
rect 28273 9877 28307 9911
rect 28307 9877 28316 9911
rect 28264 9868 28316 9877
rect 30472 9868 30524 9920
rect 32128 9945 32137 9979
rect 32137 9945 32171 9979
rect 32171 9945 32180 9979
rect 32128 9936 32180 9945
rect 32956 9936 33008 9988
rect 33784 9936 33836 9988
rect 37556 10004 37608 10056
rect 37832 10047 37884 10056
rect 37832 10013 37841 10047
rect 37841 10013 37875 10047
rect 37875 10013 37884 10047
rect 37832 10004 37884 10013
rect 37924 10004 37976 10056
rect 36360 9936 36412 9988
rect 36636 9936 36688 9988
rect 39396 9979 39448 9988
rect 39396 9945 39405 9979
rect 39405 9945 39439 9979
rect 39439 9945 39448 9979
rect 39396 9936 39448 9945
rect 30932 9911 30984 9920
rect 30932 9877 30941 9911
rect 30941 9877 30975 9911
rect 30975 9877 30984 9911
rect 30932 9868 30984 9877
rect 31392 9868 31444 9920
rect 35256 9868 35308 9920
rect 35440 9868 35492 9920
rect 37372 9868 37424 9920
rect 37464 9868 37516 9920
rect 37924 9911 37976 9920
rect 37924 9877 37933 9911
rect 37933 9877 37967 9911
rect 37967 9877 37976 9911
rect 37924 9868 37976 9877
rect 39028 9868 39080 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 8484 9664 8536 9716
rect 8668 9664 8720 9716
rect 6828 9571 6880 9580
rect 6828 9537 6837 9571
rect 6837 9537 6871 9571
rect 6871 9537 6880 9571
rect 6828 9528 6880 9537
rect 7012 9571 7064 9580
rect 7012 9537 7021 9571
rect 7021 9537 7055 9571
rect 7055 9537 7064 9571
rect 7012 9528 7064 9537
rect 7656 9528 7708 9580
rect 9312 9639 9364 9648
rect 9312 9605 9321 9639
rect 9321 9605 9355 9639
rect 9355 9605 9364 9639
rect 9312 9596 9364 9605
rect 11520 9664 11572 9716
rect 12348 9664 12400 9716
rect 14464 9707 14516 9716
rect 14464 9673 14473 9707
rect 14473 9673 14507 9707
rect 14507 9673 14516 9707
rect 14464 9664 14516 9673
rect 9128 9571 9180 9580
rect 9128 9537 9137 9571
rect 9137 9537 9171 9571
rect 9171 9537 9180 9571
rect 9128 9528 9180 9537
rect 9404 9571 9456 9580
rect 9404 9537 9413 9571
rect 9413 9537 9447 9571
rect 9447 9537 9456 9571
rect 9404 9528 9456 9537
rect 8392 9392 8444 9444
rect 8484 9392 8536 9444
rect 10232 9596 10284 9648
rect 10968 9596 11020 9648
rect 11060 9571 11112 9580
rect 11060 9537 11069 9571
rect 11069 9537 11103 9571
rect 11103 9537 11112 9571
rect 11060 9528 11112 9537
rect 11152 9571 11204 9580
rect 11152 9537 11161 9571
rect 11161 9537 11195 9571
rect 11195 9537 11204 9571
rect 11152 9528 11204 9537
rect 11428 9528 11480 9580
rect 11704 9571 11756 9580
rect 11704 9537 11713 9571
rect 11713 9537 11747 9571
rect 11747 9537 11756 9571
rect 11704 9528 11756 9537
rect 12256 9596 12308 9648
rect 15016 9664 15068 9716
rect 15384 9664 15436 9716
rect 22376 9664 22428 9716
rect 24124 9664 24176 9716
rect 10784 9503 10836 9512
rect 10784 9469 10793 9503
rect 10793 9469 10827 9503
rect 10827 9469 10836 9503
rect 10784 9460 10836 9469
rect 12808 9528 12860 9580
rect 11428 9392 11480 9444
rect 12256 9392 12308 9444
rect 12716 9460 12768 9512
rect 13176 9503 13228 9512
rect 13176 9469 13185 9503
rect 13185 9469 13219 9503
rect 13219 9469 13228 9503
rect 13176 9460 13228 9469
rect 13452 9571 13504 9580
rect 13452 9537 13461 9571
rect 13461 9537 13495 9571
rect 13495 9537 13504 9571
rect 13452 9528 13504 9537
rect 14372 9528 14424 9580
rect 14556 9460 14608 9512
rect 7104 9324 7156 9376
rect 7564 9324 7616 9376
rect 8944 9324 8996 9376
rect 9036 9324 9088 9376
rect 10876 9324 10928 9376
rect 11612 9324 11664 9376
rect 19064 9596 19116 9648
rect 15384 9571 15436 9580
rect 15384 9537 15393 9571
rect 15393 9537 15427 9571
rect 15427 9537 15436 9571
rect 15384 9528 15436 9537
rect 15844 9528 15896 9580
rect 15936 9571 15988 9580
rect 15936 9537 15945 9571
rect 15945 9537 15979 9571
rect 15979 9537 15988 9571
rect 15936 9528 15988 9537
rect 17040 9528 17092 9580
rect 17776 9528 17828 9580
rect 19248 9528 19300 9580
rect 19340 9528 19392 9580
rect 20536 9571 20588 9580
rect 20536 9537 20545 9571
rect 20545 9537 20579 9571
rect 20579 9537 20588 9571
rect 20536 9528 20588 9537
rect 20812 9528 20864 9580
rect 17500 9460 17552 9512
rect 15016 9392 15068 9444
rect 15936 9392 15988 9444
rect 18696 9460 18748 9512
rect 21180 9460 21232 9512
rect 19340 9392 19392 9444
rect 22560 9596 22612 9648
rect 23112 9596 23164 9648
rect 22008 9460 22060 9512
rect 22284 9528 22336 9580
rect 22192 9503 22244 9512
rect 22192 9469 22201 9503
rect 22201 9469 22235 9503
rect 22235 9469 22244 9503
rect 22192 9460 22244 9469
rect 23940 9528 23992 9580
rect 25320 9707 25372 9716
rect 25320 9673 25329 9707
rect 25329 9673 25363 9707
rect 25363 9673 25372 9707
rect 25320 9664 25372 9673
rect 28632 9707 28684 9716
rect 28632 9673 28641 9707
rect 28641 9673 28675 9707
rect 28675 9673 28684 9707
rect 28632 9664 28684 9673
rect 30748 9664 30800 9716
rect 34428 9664 34480 9716
rect 25596 9596 25648 9648
rect 26792 9596 26844 9648
rect 27068 9596 27120 9648
rect 27896 9596 27948 9648
rect 29092 9596 29144 9648
rect 29828 9639 29880 9648
rect 29828 9605 29837 9639
rect 29837 9605 29871 9639
rect 29871 9605 29880 9639
rect 29828 9596 29880 9605
rect 25136 9460 25188 9512
rect 26884 9528 26936 9580
rect 27436 9528 27488 9580
rect 28448 9528 28500 9580
rect 25688 9460 25740 9512
rect 26424 9460 26476 9512
rect 27068 9460 27120 9512
rect 27344 9503 27396 9512
rect 27344 9469 27353 9503
rect 27353 9469 27387 9503
rect 27387 9469 27396 9503
rect 27344 9460 27396 9469
rect 27896 9503 27948 9512
rect 27896 9469 27905 9503
rect 27905 9469 27939 9503
rect 27939 9469 27948 9503
rect 27896 9460 27948 9469
rect 29828 9460 29880 9512
rect 30932 9596 30984 9648
rect 31392 9639 31444 9648
rect 31392 9605 31401 9639
rect 31401 9605 31435 9639
rect 31435 9605 31444 9639
rect 31392 9596 31444 9605
rect 30380 9528 30432 9580
rect 31024 9571 31076 9580
rect 31024 9537 31033 9571
rect 31033 9537 31067 9571
rect 31067 9537 31076 9571
rect 31024 9528 31076 9537
rect 14464 9324 14516 9376
rect 15844 9324 15896 9376
rect 17592 9324 17644 9376
rect 20352 9324 20404 9376
rect 20904 9367 20956 9376
rect 20904 9333 20913 9367
rect 20913 9333 20947 9367
rect 20947 9333 20956 9367
rect 20904 9324 20956 9333
rect 22560 9367 22612 9376
rect 22560 9333 22569 9367
rect 22569 9333 22603 9367
rect 22603 9333 22612 9367
rect 22560 9324 22612 9333
rect 30104 9392 30156 9444
rect 30288 9435 30340 9444
rect 30288 9401 30297 9435
rect 30297 9401 30331 9435
rect 30331 9401 30340 9435
rect 30288 9392 30340 9401
rect 30748 9435 30800 9444
rect 30748 9401 30757 9435
rect 30757 9401 30791 9435
rect 30791 9401 30800 9435
rect 30748 9392 30800 9401
rect 25228 9324 25280 9376
rect 25412 9324 25464 9376
rect 25964 9324 26016 9376
rect 26240 9324 26292 9376
rect 27620 9324 27672 9376
rect 27804 9324 27856 9376
rect 28632 9324 28684 9376
rect 29000 9324 29052 9376
rect 30380 9367 30432 9376
rect 30380 9333 30389 9367
rect 30389 9333 30423 9367
rect 30423 9333 30432 9367
rect 30380 9324 30432 9333
rect 30472 9324 30524 9376
rect 35348 9664 35400 9716
rect 35624 9596 35676 9648
rect 36268 9664 36320 9716
rect 36636 9664 36688 9716
rect 36084 9639 36136 9648
rect 36084 9605 36093 9639
rect 36093 9605 36127 9639
rect 36127 9605 36136 9639
rect 36084 9596 36136 9605
rect 32128 9571 32180 9580
rect 32128 9537 32137 9571
rect 32137 9537 32171 9571
rect 32171 9537 32180 9571
rect 32128 9528 32180 9537
rect 32588 9528 32640 9580
rect 32680 9571 32732 9580
rect 32680 9537 32689 9571
rect 32689 9537 32723 9571
rect 32723 9537 32732 9571
rect 32680 9528 32732 9537
rect 32864 9571 32916 9580
rect 32864 9537 32873 9571
rect 32873 9537 32907 9571
rect 32907 9537 32916 9571
rect 32864 9528 32916 9537
rect 33324 9528 33376 9580
rect 33876 9528 33928 9580
rect 34152 9528 34204 9580
rect 33600 9460 33652 9512
rect 34520 9571 34572 9580
rect 34520 9537 34529 9571
rect 34529 9537 34563 9571
rect 34563 9537 34572 9571
rect 34520 9528 34572 9537
rect 34704 9571 34756 9580
rect 34704 9537 34718 9571
rect 34718 9537 34752 9571
rect 34752 9537 34756 9571
rect 34704 9528 34756 9537
rect 34888 9528 34940 9580
rect 35348 9571 35400 9580
rect 35348 9537 35357 9571
rect 35357 9537 35391 9571
rect 35391 9537 35400 9571
rect 35348 9528 35400 9537
rect 35532 9571 35584 9580
rect 35532 9537 35541 9571
rect 35541 9537 35575 9571
rect 35575 9537 35584 9571
rect 35532 9528 35584 9537
rect 35992 9571 36044 9580
rect 35992 9537 36009 9571
rect 36009 9537 36044 9571
rect 35992 9528 36044 9537
rect 36452 9596 36504 9648
rect 37740 9639 37792 9648
rect 37740 9605 37749 9639
rect 37749 9605 37783 9639
rect 37783 9605 37792 9639
rect 37740 9596 37792 9605
rect 38016 9639 38068 9648
rect 38016 9605 38025 9639
rect 38025 9605 38059 9639
rect 38059 9605 38068 9639
rect 38016 9596 38068 9605
rect 39948 9596 40000 9648
rect 36268 9571 36320 9580
rect 36268 9537 36277 9571
rect 36277 9537 36311 9571
rect 36311 9537 36320 9571
rect 36268 9528 36320 9537
rect 36544 9528 36596 9580
rect 37648 9571 37700 9580
rect 37648 9537 37657 9571
rect 37657 9537 37691 9571
rect 37691 9537 37700 9571
rect 37648 9528 37700 9537
rect 36360 9460 36412 9512
rect 37188 9460 37240 9512
rect 36176 9392 36228 9444
rect 36268 9392 36320 9444
rect 34612 9324 34664 9376
rect 35532 9324 35584 9376
rect 37464 9435 37516 9444
rect 37464 9401 37473 9435
rect 37473 9401 37507 9435
rect 37507 9401 37516 9435
rect 37464 9392 37516 9401
rect 37556 9392 37608 9444
rect 36820 9324 36872 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 9128 9120 9180 9172
rect 9864 9120 9916 9172
rect 10324 9120 10376 9172
rect 10692 9120 10744 9172
rect 5264 8984 5316 9036
rect 6828 8984 6880 9036
rect 7748 9052 7800 9104
rect 8024 9052 8076 9104
rect 7104 8916 7156 8968
rect 7288 8959 7340 8968
rect 7288 8925 7297 8959
rect 7297 8925 7331 8959
rect 7331 8925 7340 8959
rect 7288 8916 7340 8925
rect 8116 8984 8168 9036
rect 7012 8891 7064 8900
rect 7012 8857 7021 8891
rect 7021 8857 7055 8891
rect 7055 8857 7064 8891
rect 7012 8848 7064 8857
rect 7840 8916 7892 8968
rect 8944 8984 8996 9036
rect 9036 8916 9088 8968
rect 6644 8780 6696 8832
rect 7104 8780 7156 8832
rect 7472 8780 7524 8832
rect 10784 9052 10836 9104
rect 13176 9120 13228 9172
rect 20352 9163 20404 9172
rect 20352 9129 20361 9163
rect 20361 9129 20395 9163
rect 20395 9129 20404 9163
rect 20352 9120 20404 9129
rect 20996 9163 21048 9172
rect 20996 9129 21005 9163
rect 21005 9129 21039 9163
rect 21039 9129 21048 9163
rect 20996 9120 21048 9129
rect 22192 9120 22244 9172
rect 10416 8916 10468 8968
rect 10508 8959 10560 8968
rect 10508 8925 10517 8959
rect 10517 8925 10551 8959
rect 10551 8925 10560 8959
rect 10508 8916 10560 8925
rect 10600 8959 10652 8968
rect 10600 8925 10609 8959
rect 10609 8925 10643 8959
rect 10643 8925 10652 8959
rect 10600 8916 10652 8925
rect 11336 8984 11388 9036
rect 11152 8959 11204 8968
rect 11152 8925 11161 8959
rect 11161 8925 11195 8959
rect 11195 8925 11204 8959
rect 11152 8916 11204 8925
rect 11428 8959 11480 8968
rect 11428 8925 11437 8959
rect 11437 8925 11471 8959
rect 11471 8925 11480 8959
rect 11428 8916 11480 8925
rect 11060 8848 11112 8900
rect 12532 9052 12584 9104
rect 20812 9052 20864 9104
rect 23480 9120 23532 9172
rect 24584 9163 24636 9172
rect 24584 9129 24593 9163
rect 24593 9129 24627 9163
rect 24627 9129 24636 9163
rect 24584 9120 24636 9129
rect 25044 9163 25096 9172
rect 25044 9129 25053 9163
rect 25053 9129 25087 9163
rect 25087 9129 25096 9163
rect 25044 9120 25096 9129
rect 22560 9052 22612 9104
rect 24124 9052 24176 9104
rect 25136 9052 25188 9104
rect 25320 9120 25372 9172
rect 26148 9120 26200 9172
rect 26240 9120 26292 9172
rect 26884 9163 26936 9172
rect 26884 9129 26893 9163
rect 26893 9129 26927 9163
rect 26927 9129 26936 9163
rect 26884 9120 26936 9129
rect 27620 9120 27672 9172
rect 27712 9163 27764 9172
rect 27712 9129 27721 9163
rect 27721 9129 27755 9163
rect 27755 9129 27764 9163
rect 27712 9120 27764 9129
rect 28356 9120 28408 9172
rect 31116 9120 31168 9172
rect 31484 9163 31536 9172
rect 31484 9129 31493 9163
rect 31493 9129 31527 9163
rect 31527 9129 31536 9163
rect 31484 9120 31536 9129
rect 28540 9052 28592 9104
rect 28908 9095 28960 9104
rect 28908 9061 28917 9095
rect 28917 9061 28951 9095
rect 28951 9061 28960 9095
rect 28908 9052 28960 9061
rect 12256 8916 12308 8968
rect 12348 8959 12400 8968
rect 12348 8925 12357 8959
rect 12357 8925 12391 8959
rect 12391 8925 12400 8959
rect 12348 8916 12400 8925
rect 12716 8984 12768 9036
rect 15476 9027 15528 9036
rect 15476 8993 15485 9027
rect 15485 8993 15519 9027
rect 15519 8993 15528 9027
rect 15476 8984 15528 8993
rect 17408 8984 17460 9036
rect 14648 8916 14700 8968
rect 16488 8916 16540 8968
rect 18236 8984 18288 9036
rect 8392 8780 8444 8832
rect 10324 8823 10376 8832
rect 10324 8789 10333 8823
rect 10333 8789 10367 8823
rect 10367 8789 10376 8823
rect 10324 8780 10376 8789
rect 10416 8780 10468 8832
rect 11152 8780 11204 8832
rect 12532 8848 12584 8900
rect 18328 8916 18380 8968
rect 17776 8848 17828 8900
rect 19616 8848 19668 8900
rect 20168 8848 20220 8900
rect 20260 8848 20312 8900
rect 20720 8891 20772 8900
rect 20720 8857 20729 8891
rect 20729 8857 20763 8891
rect 20763 8857 20772 8891
rect 20720 8848 20772 8857
rect 26240 8984 26292 9036
rect 26424 8984 26476 9036
rect 27528 8984 27580 9036
rect 30472 9052 30524 9104
rect 30564 9052 30616 9104
rect 33692 9120 33744 9172
rect 35348 9120 35400 9172
rect 37648 9163 37700 9172
rect 37648 9129 37657 9163
rect 37657 9129 37691 9163
rect 37691 9129 37700 9163
rect 37648 9120 37700 9129
rect 38016 9120 38068 9172
rect 11888 8780 11940 8832
rect 12256 8780 12308 8832
rect 15384 8780 15436 8832
rect 19984 8780 20036 8832
rect 20628 8780 20680 8832
rect 23112 8916 23164 8968
rect 24216 8959 24268 8968
rect 24216 8925 24225 8959
rect 24225 8925 24259 8959
rect 24259 8925 24268 8959
rect 24216 8916 24268 8925
rect 24768 8916 24820 8968
rect 25044 8916 25096 8968
rect 22744 8848 22796 8900
rect 23020 8848 23072 8900
rect 24400 8891 24452 8900
rect 24400 8857 24409 8891
rect 24409 8857 24443 8891
rect 24443 8857 24452 8891
rect 24400 8848 24452 8857
rect 22928 8780 22980 8832
rect 24032 8780 24084 8832
rect 25412 8916 25464 8968
rect 26056 8916 26108 8968
rect 26332 8959 26384 8968
rect 26332 8925 26341 8959
rect 26341 8925 26375 8959
rect 26375 8925 26384 8959
rect 26332 8916 26384 8925
rect 27068 8916 27120 8968
rect 27344 8959 27396 8968
rect 27344 8925 27353 8959
rect 27353 8925 27387 8959
rect 27387 8925 27396 8959
rect 27344 8916 27396 8925
rect 24768 8823 24820 8832
rect 24768 8789 24777 8823
rect 24777 8789 24811 8823
rect 24811 8789 24820 8823
rect 24768 8780 24820 8789
rect 25320 8891 25372 8900
rect 25320 8857 25329 8891
rect 25329 8857 25363 8891
rect 25363 8857 25372 8891
rect 25320 8848 25372 8857
rect 25228 8823 25280 8832
rect 25228 8789 25237 8823
rect 25237 8789 25271 8823
rect 25271 8789 25280 8823
rect 25228 8780 25280 8789
rect 25688 8823 25740 8832
rect 25688 8789 25697 8823
rect 25697 8789 25731 8823
rect 25731 8789 25740 8823
rect 25688 8780 25740 8789
rect 26700 8848 26752 8900
rect 29184 8984 29236 9036
rect 28264 8959 28316 8968
rect 28264 8925 28273 8959
rect 28273 8925 28307 8959
rect 28307 8925 28316 8959
rect 28264 8916 28316 8925
rect 28724 8959 28776 8968
rect 28724 8925 28733 8959
rect 28733 8925 28767 8959
rect 28767 8925 28776 8959
rect 28724 8916 28776 8925
rect 28632 8848 28684 8900
rect 29736 8959 29788 8968
rect 29736 8925 29745 8959
rect 29745 8925 29779 8959
rect 29779 8925 29788 8959
rect 29736 8916 29788 8925
rect 30104 8959 30156 8968
rect 30104 8925 30113 8959
rect 30113 8925 30147 8959
rect 30147 8925 30156 8959
rect 30104 8916 30156 8925
rect 30656 8959 30708 8968
rect 30656 8925 30665 8959
rect 30665 8925 30699 8959
rect 30699 8925 30708 8959
rect 30656 8916 30708 8925
rect 29092 8848 29144 8900
rect 30380 8891 30432 8900
rect 30380 8857 30389 8891
rect 30389 8857 30423 8891
rect 30423 8857 30432 8891
rect 30380 8848 30432 8857
rect 31116 8959 31168 8968
rect 31116 8925 31125 8959
rect 31125 8925 31159 8959
rect 31159 8925 31168 8959
rect 31116 8916 31168 8925
rect 31208 8916 31260 8968
rect 32404 8984 32456 9036
rect 32588 8916 32640 8968
rect 32864 8916 32916 8968
rect 33416 8984 33468 9036
rect 35164 8916 35216 8968
rect 35440 8916 35492 8968
rect 36084 8916 36136 8968
rect 37556 8916 37608 8968
rect 31484 8848 31536 8900
rect 33324 8891 33376 8900
rect 33324 8857 33333 8891
rect 33333 8857 33367 8891
rect 33367 8857 33376 8891
rect 33324 8848 33376 8857
rect 33600 8848 33652 8900
rect 34428 8848 34480 8900
rect 36176 8848 36228 8900
rect 37740 8916 37792 8968
rect 37924 8959 37976 8968
rect 37924 8925 37933 8959
rect 37933 8925 37967 8959
rect 37967 8925 37976 8959
rect 37924 8916 37976 8925
rect 26332 8780 26384 8832
rect 28540 8780 28592 8832
rect 28908 8780 28960 8832
rect 30932 8780 30984 8832
rect 32680 8780 32732 8832
rect 34520 8780 34572 8832
rect 34980 8780 35032 8832
rect 35256 8780 35308 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 5632 8576 5684 8628
rect 6920 8576 6972 8628
rect 7564 8576 7616 8628
rect 8484 8576 8536 8628
rect 4712 8508 4764 8560
rect 8300 8508 8352 8560
rect 6644 8483 6696 8492
rect 6644 8449 6653 8483
rect 6653 8449 6687 8483
rect 6687 8449 6696 8483
rect 6644 8440 6696 8449
rect 6828 8483 6880 8492
rect 6828 8449 6837 8483
rect 6837 8449 6871 8483
rect 6871 8449 6880 8483
rect 6828 8440 6880 8449
rect 7104 8440 7156 8492
rect 7196 8440 7248 8492
rect 7472 8483 7524 8492
rect 7472 8449 7481 8483
rect 7481 8449 7515 8483
rect 7515 8449 7524 8483
rect 7472 8440 7524 8449
rect 5724 8415 5776 8424
rect 5724 8381 5733 8415
rect 5733 8381 5767 8415
rect 5767 8381 5776 8415
rect 5724 8372 5776 8381
rect 7012 8372 7064 8424
rect 7288 8372 7340 8424
rect 7748 8483 7800 8492
rect 7748 8449 7757 8483
rect 7757 8449 7791 8483
rect 7791 8449 7800 8483
rect 7748 8440 7800 8449
rect 6460 8279 6512 8288
rect 6460 8245 6469 8279
rect 6469 8245 6503 8279
rect 6503 8245 6512 8279
rect 6460 8236 6512 8245
rect 8208 8483 8260 8492
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 8484 8440 8536 8492
rect 8944 8619 8996 8628
rect 8944 8585 8953 8619
rect 8953 8585 8987 8619
rect 8987 8585 8996 8619
rect 8944 8576 8996 8585
rect 11428 8576 11480 8628
rect 9864 8508 9916 8560
rect 9036 8483 9088 8492
rect 9036 8449 9045 8483
rect 9045 8449 9079 8483
rect 9079 8449 9088 8483
rect 9036 8440 9088 8449
rect 9128 8440 9180 8492
rect 10416 8440 10468 8492
rect 7932 8415 7984 8424
rect 7932 8381 7941 8415
rect 7941 8381 7975 8415
rect 7975 8381 7984 8415
rect 7932 8372 7984 8381
rect 8300 8415 8352 8424
rect 8300 8381 8334 8415
rect 8334 8381 8352 8415
rect 8300 8372 8352 8381
rect 8668 8372 8720 8424
rect 10876 8483 10928 8492
rect 10876 8449 10885 8483
rect 10885 8449 10919 8483
rect 10919 8449 10928 8483
rect 10876 8440 10928 8449
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 12532 8440 12584 8492
rect 10968 8372 11020 8424
rect 15568 8576 15620 8628
rect 14372 8508 14424 8560
rect 14740 8508 14792 8560
rect 17868 8576 17920 8628
rect 18788 8576 18840 8628
rect 20076 8576 20128 8628
rect 15200 8483 15252 8492
rect 15200 8449 15209 8483
rect 15209 8449 15243 8483
rect 15243 8449 15252 8483
rect 15200 8440 15252 8449
rect 15292 8483 15344 8492
rect 15292 8449 15301 8483
rect 15301 8449 15335 8483
rect 15335 8449 15344 8483
rect 15292 8440 15344 8449
rect 8116 8236 8168 8288
rect 8484 8304 8536 8356
rect 14740 8372 14792 8424
rect 15384 8372 15436 8424
rect 15660 8483 15712 8492
rect 15660 8449 15669 8483
rect 15669 8449 15703 8483
rect 15703 8449 15712 8483
rect 15660 8440 15712 8449
rect 17592 8483 17644 8492
rect 17592 8449 17601 8483
rect 17601 8449 17635 8483
rect 17635 8449 17644 8483
rect 17592 8440 17644 8449
rect 19432 8508 19484 8560
rect 18696 8483 18748 8492
rect 18696 8449 18705 8483
rect 18705 8449 18739 8483
rect 18739 8449 18748 8483
rect 18696 8440 18748 8449
rect 18788 8440 18840 8492
rect 19156 8440 19208 8492
rect 19616 8483 19668 8492
rect 19616 8449 19625 8483
rect 19625 8449 19659 8483
rect 19659 8449 19668 8483
rect 19616 8440 19668 8449
rect 17316 8372 17368 8424
rect 17684 8415 17736 8424
rect 17684 8381 17693 8415
rect 17693 8381 17727 8415
rect 17727 8381 17736 8415
rect 17684 8372 17736 8381
rect 17960 8372 18012 8424
rect 19248 8372 19300 8424
rect 20260 8508 20312 8560
rect 19984 8440 20036 8492
rect 20076 8483 20128 8492
rect 20076 8449 20085 8483
rect 20085 8449 20119 8483
rect 20119 8449 20128 8483
rect 20076 8440 20128 8449
rect 20996 8576 21048 8628
rect 20720 8508 20772 8560
rect 20628 8483 20680 8492
rect 20628 8449 20637 8483
rect 20637 8449 20671 8483
rect 20671 8449 20680 8483
rect 20628 8440 20680 8449
rect 20812 8483 20864 8492
rect 20812 8449 20821 8483
rect 20821 8449 20855 8483
rect 20855 8449 20864 8483
rect 20812 8440 20864 8449
rect 21180 8440 21232 8492
rect 22284 8508 22336 8560
rect 22744 8440 22796 8492
rect 21732 8372 21784 8424
rect 22652 8372 22704 8424
rect 23112 8619 23164 8628
rect 23112 8585 23121 8619
rect 23121 8585 23155 8619
rect 23155 8585 23164 8619
rect 23112 8576 23164 8585
rect 23296 8576 23348 8628
rect 23848 8576 23900 8628
rect 23756 8551 23808 8560
rect 23756 8517 23765 8551
rect 23765 8517 23799 8551
rect 23799 8517 23808 8551
rect 23756 8508 23808 8517
rect 24124 8551 24176 8560
rect 24124 8517 24133 8551
rect 24133 8517 24167 8551
rect 24167 8517 24176 8551
rect 24124 8508 24176 8517
rect 24216 8551 24268 8560
rect 24216 8517 24225 8551
rect 24225 8517 24259 8551
rect 24259 8517 24268 8551
rect 24216 8508 24268 8517
rect 24952 8576 25004 8628
rect 27068 8619 27120 8628
rect 27068 8585 27077 8619
rect 27077 8585 27111 8619
rect 27111 8585 27120 8619
rect 27068 8576 27120 8585
rect 26148 8508 26200 8560
rect 27436 8508 27488 8560
rect 24032 8483 24084 8492
rect 24032 8449 24041 8483
rect 24041 8449 24075 8483
rect 24075 8449 24084 8483
rect 24032 8440 24084 8449
rect 24584 8440 24636 8492
rect 24768 8372 24820 8424
rect 25228 8483 25280 8492
rect 25228 8449 25237 8483
rect 25237 8449 25271 8483
rect 25271 8449 25280 8483
rect 25228 8440 25280 8449
rect 25688 8483 25740 8492
rect 25688 8449 25697 8483
rect 25697 8449 25731 8483
rect 25731 8449 25740 8483
rect 25688 8440 25740 8449
rect 25780 8440 25832 8492
rect 26700 8483 26752 8492
rect 26700 8449 26709 8483
rect 26709 8449 26743 8483
rect 26743 8449 26752 8483
rect 26700 8440 26752 8449
rect 27528 8440 27580 8492
rect 27712 8508 27764 8560
rect 28632 8619 28684 8628
rect 28632 8585 28641 8619
rect 28641 8585 28675 8619
rect 28675 8585 28684 8619
rect 28632 8576 28684 8585
rect 28724 8619 28776 8628
rect 28724 8585 28733 8619
rect 28733 8585 28767 8619
rect 28767 8585 28776 8619
rect 28724 8576 28776 8585
rect 28816 8576 28868 8628
rect 31208 8576 31260 8628
rect 33784 8619 33836 8628
rect 33784 8585 33793 8619
rect 33793 8585 33827 8619
rect 33827 8585 33836 8619
rect 33784 8576 33836 8585
rect 33968 8576 34020 8628
rect 29000 8508 29052 8560
rect 27068 8372 27120 8424
rect 27344 8372 27396 8424
rect 28908 8483 28960 8492
rect 28908 8449 28917 8483
rect 28917 8449 28951 8483
rect 28951 8449 28960 8483
rect 28908 8440 28960 8449
rect 29092 8440 29144 8492
rect 29828 8508 29880 8560
rect 29736 8483 29788 8492
rect 29736 8449 29745 8483
rect 29745 8449 29779 8483
rect 29779 8449 29788 8483
rect 29736 8440 29788 8449
rect 30012 8415 30064 8424
rect 30012 8381 30021 8415
rect 30021 8381 30055 8415
rect 30055 8381 30064 8415
rect 30012 8372 30064 8381
rect 30656 8483 30708 8492
rect 30656 8449 30665 8483
rect 30665 8449 30699 8483
rect 30699 8449 30708 8483
rect 30656 8440 30708 8449
rect 31576 8440 31628 8492
rect 31760 8440 31812 8492
rect 34060 8508 34112 8560
rect 34244 8619 34296 8628
rect 34244 8585 34253 8619
rect 34253 8585 34287 8619
rect 34287 8585 34296 8619
rect 34244 8576 34296 8585
rect 34520 8619 34572 8628
rect 34520 8585 34529 8619
rect 34529 8585 34563 8619
rect 34563 8585 34572 8619
rect 34520 8576 34572 8585
rect 36084 8619 36136 8628
rect 36084 8585 36093 8619
rect 36093 8585 36127 8619
rect 36127 8585 36136 8619
rect 36084 8576 36136 8585
rect 36176 8619 36228 8628
rect 36176 8585 36185 8619
rect 36185 8585 36219 8619
rect 36219 8585 36228 8619
rect 36176 8576 36228 8585
rect 37740 8576 37792 8628
rect 38568 8576 38620 8628
rect 35440 8508 35492 8560
rect 37464 8508 37516 8560
rect 39028 8508 39080 8560
rect 32588 8483 32640 8492
rect 32588 8449 32597 8483
rect 32597 8449 32631 8483
rect 32631 8449 32640 8483
rect 32588 8440 32640 8449
rect 33968 8440 34020 8492
rect 30748 8372 30800 8424
rect 30932 8372 30984 8424
rect 33048 8372 33100 8424
rect 33876 8372 33928 8424
rect 36544 8440 36596 8492
rect 37740 8483 37792 8492
rect 37740 8449 37749 8483
rect 37749 8449 37783 8483
rect 37783 8449 37792 8483
rect 37740 8440 37792 8449
rect 8392 8236 8444 8288
rect 9128 8236 9180 8288
rect 15108 8236 15160 8288
rect 18328 8304 18380 8356
rect 18880 8304 18932 8356
rect 22192 8347 22244 8356
rect 22192 8313 22201 8347
rect 22201 8313 22235 8347
rect 22235 8313 22244 8347
rect 22192 8304 22244 8313
rect 23940 8304 23992 8356
rect 28264 8304 28316 8356
rect 28448 8304 28500 8356
rect 15844 8236 15896 8288
rect 18420 8279 18472 8288
rect 18420 8245 18429 8279
rect 18429 8245 18463 8279
rect 18463 8245 18472 8279
rect 18420 8236 18472 8245
rect 20444 8236 20496 8288
rect 20904 8236 20956 8288
rect 21640 8236 21692 8288
rect 21824 8236 21876 8288
rect 23480 8236 23532 8288
rect 23848 8279 23900 8288
rect 23848 8245 23857 8279
rect 23857 8245 23891 8279
rect 23891 8245 23900 8279
rect 23848 8236 23900 8245
rect 26424 8236 26476 8288
rect 26976 8236 27028 8288
rect 27804 8236 27856 8288
rect 28632 8236 28684 8288
rect 29000 8347 29052 8356
rect 29000 8313 29009 8347
rect 29009 8313 29043 8347
rect 29043 8313 29052 8347
rect 29000 8304 29052 8313
rect 29828 8236 29880 8288
rect 30196 8236 30248 8288
rect 30380 8236 30432 8288
rect 31024 8236 31076 8288
rect 32312 8236 32364 8288
rect 33692 8347 33744 8356
rect 33692 8313 33701 8347
rect 33701 8313 33735 8347
rect 33735 8313 33744 8347
rect 33692 8304 33744 8313
rect 34520 8372 34572 8424
rect 34704 8304 34756 8356
rect 34980 8372 35032 8424
rect 36176 8304 36228 8356
rect 38476 8415 38528 8424
rect 38476 8381 38485 8415
rect 38485 8381 38519 8415
rect 38519 8381 38528 8415
rect 38476 8372 38528 8381
rect 37556 8304 37608 8356
rect 35164 8236 35216 8288
rect 37832 8236 37884 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 5724 8032 5776 8084
rect 6736 8032 6788 8084
rect 7932 8032 7984 8084
rect 8208 8032 8260 8084
rect 7196 7964 7248 8016
rect 5632 7939 5684 7948
rect 5632 7905 5641 7939
rect 5641 7905 5675 7939
rect 5675 7905 5684 7939
rect 5632 7896 5684 7905
rect 6552 7896 6604 7948
rect 6460 7828 6512 7880
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 7932 7939 7984 7948
rect 7932 7905 7941 7939
rect 7941 7905 7975 7939
rect 7975 7905 7984 7939
rect 7932 7896 7984 7905
rect 7564 7871 7616 7880
rect 7564 7837 7573 7871
rect 7573 7837 7607 7871
rect 7607 7837 7616 7871
rect 7564 7828 7616 7837
rect 7840 7871 7892 7880
rect 7840 7837 7849 7871
rect 7849 7837 7883 7871
rect 7883 7837 7892 7871
rect 7840 7828 7892 7837
rect 9036 7964 9088 8016
rect 11888 8032 11940 8084
rect 11980 8032 12032 8084
rect 12716 8032 12768 8084
rect 15200 8032 15252 8084
rect 15292 8075 15344 8084
rect 15292 8041 15301 8075
rect 15301 8041 15335 8075
rect 15335 8041 15344 8075
rect 15292 8032 15344 8041
rect 8300 7896 8352 7948
rect 8392 7939 8444 7948
rect 8392 7905 8401 7939
rect 8401 7905 8435 7939
rect 8435 7905 8444 7939
rect 8392 7896 8444 7905
rect 10968 7964 11020 8016
rect 11428 7964 11480 8016
rect 15108 8007 15160 8016
rect 15108 7973 15117 8007
rect 15117 7973 15151 8007
rect 15151 7973 15160 8007
rect 15108 7964 15160 7973
rect 15568 7964 15620 8016
rect 9864 7939 9916 7948
rect 9864 7905 9873 7939
rect 9873 7905 9907 7939
rect 9907 7905 9916 7939
rect 9864 7896 9916 7905
rect 10324 7896 10376 7948
rect 10692 7896 10744 7948
rect 14004 7828 14056 7880
rect 14096 7871 14148 7880
rect 14096 7837 14105 7871
rect 14105 7837 14139 7871
rect 14139 7837 14148 7871
rect 14096 7828 14148 7837
rect 11612 7760 11664 7812
rect 11796 7760 11848 7812
rect 14740 7828 14792 7880
rect 15292 7828 15344 7880
rect 16672 8032 16724 8084
rect 17316 8032 17368 8084
rect 18788 8075 18840 8084
rect 18788 8041 18797 8075
rect 18797 8041 18831 8075
rect 18831 8041 18840 8075
rect 18788 8032 18840 8041
rect 19432 8075 19484 8084
rect 19432 8041 19441 8075
rect 19441 8041 19475 8075
rect 19475 8041 19484 8075
rect 19432 8032 19484 8041
rect 15752 7896 15804 7948
rect 16304 7896 16356 7948
rect 20352 7964 20404 8016
rect 20628 7964 20680 8016
rect 22376 7964 22428 8016
rect 22836 7964 22888 8016
rect 15844 7871 15896 7880
rect 15844 7837 15853 7871
rect 15853 7837 15887 7871
rect 15887 7837 15896 7871
rect 15844 7828 15896 7837
rect 15936 7871 15988 7880
rect 15936 7837 15945 7871
rect 15945 7837 15979 7871
rect 15979 7837 15988 7871
rect 15936 7828 15988 7837
rect 18144 7828 18196 7880
rect 19340 7896 19392 7948
rect 19156 7828 19208 7880
rect 20720 7896 20772 7948
rect 20904 7939 20956 7948
rect 20904 7905 20913 7939
rect 20913 7905 20947 7939
rect 20947 7905 20956 7939
rect 20904 7896 20956 7905
rect 21824 7896 21876 7948
rect 16764 7760 16816 7812
rect 17776 7760 17828 7812
rect 18972 7760 19024 7812
rect 20076 7828 20128 7880
rect 20352 7871 20404 7880
rect 20352 7837 20361 7871
rect 20361 7837 20395 7871
rect 20395 7837 20404 7871
rect 20352 7828 20404 7837
rect 20536 7828 20588 7880
rect 22100 7871 22152 7880
rect 22100 7837 22109 7871
rect 22109 7837 22143 7871
rect 22143 7837 22152 7871
rect 22100 7828 22152 7837
rect 20628 7760 20680 7812
rect 22284 7871 22336 7880
rect 22284 7837 22293 7871
rect 22293 7837 22327 7871
rect 22327 7837 22336 7871
rect 22284 7828 22336 7837
rect 22468 7828 22520 7880
rect 22744 7871 22796 7880
rect 22744 7837 22753 7871
rect 22753 7837 22787 7871
rect 22787 7837 22796 7871
rect 22744 7828 22796 7837
rect 23020 7939 23072 7948
rect 23020 7905 23029 7939
rect 23029 7905 23063 7939
rect 23063 7905 23072 7939
rect 23020 7896 23072 7905
rect 23388 8075 23440 8084
rect 23388 8041 23397 8075
rect 23397 8041 23431 8075
rect 23431 8041 23440 8075
rect 23388 8032 23440 8041
rect 24676 8075 24728 8084
rect 24676 8041 24685 8075
rect 24685 8041 24719 8075
rect 24719 8041 24728 8075
rect 24676 8032 24728 8041
rect 25504 8075 25556 8084
rect 25504 8041 25513 8075
rect 25513 8041 25547 8075
rect 25547 8041 25556 8075
rect 25504 8032 25556 8041
rect 26056 8032 26108 8084
rect 25780 7896 25832 7948
rect 9496 7735 9548 7744
rect 9496 7701 9505 7735
rect 9505 7701 9539 7735
rect 9539 7701 9548 7735
rect 9496 7692 9548 7701
rect 13820 7735 13872 7744
rect 13820 7701 13829 7735
rect 13829 7701 13863 7735
rect 13863 7701 13872 7735
rect 13820 7692 13872 7701
rect 14556 7692 14608 7744
rect 15292 7692 15344 7744
rect 20076 7692 20128 7744
rect 22652 7760 22704 7812
rect 24124 7871 24176 7880
rect 24124 7837 24133 7871
rect 24133 7837 24167 7871
rect 24167 7837 24176 7871
rect 24124 7828 24176 7837
rect 26424 8032 26476 8084
rect 26516 8032 26568 8084
rect 27436 8032 27488 8084
rect 28264 8075 28316 8084
rect 28264 8041 28273 8075
rect 28273 8041 28307 8075
rect 28307 8041 28316 8075
rect 28264 8032 28316 8041
rect 28632 8075 28684 8084
rect 28632 8041 28641 8075
rect 28641 8041 28675 8075
rect 28675 8041 28684 8075
rect 28632 8032 28684 8041
rect 30288 8032 30340 8084
rect 30380 8075 30432 8084
rect 30380 8041 30389 8075
rect 30389 8041 30423 8075
rect 30423 8041 30432 8075
rect 30380 8032 30432 8041
rect 30748 8032 30800 8084
rect 31576 8032 31628 8084
rect 26792 8007 26844 8016
rect 26792 7973 26801 8007
rect 26801 7973 26835 8007
rect 26835 7973 26844 8007
rect 26792 7964 26844 7973
rect 26240 7939 26292 7948
rect 26240 7905 26249 7939
rect 26249 7905 26283 7939
rect 26283 7905 26292 7939
rect 26240 7896 26292 7905
rect 26608 7896 26660 7948
rect 27528 7964 27580 8016
rect 28172 7964 28224 8016
rect 36176 8032 36228 8084
rect 36820 8032 36872 8084
rect 27068 7939 27120 7948
rect 27068 7905 27077 7939
rect 27077 7905 27111 7939
rect 27111 7905 27120 7939
rect 27068 7896 27120 7905
rect 27160 7896 27212 7948
rect 29000 7896 29052 7948
rect 31392 7939 31444 7948
rect 22928 7692 22980 7744
rect 24492 7692 24544 7744
rect 24768 7692 24820 7744
rect 25044 7735 25096 7744
rect 25044 7701 25053 7735
rect 25053 7701 25087 7735
rect 25087 7701 25096 7735
rect 25044 7692 25096 7701
rect 27804 7828 27856 7880
rect 28816 7871 28868 7880
rect 28816 7837 28825 7871
rect 28825 7837 28859 7871
rect 28859 7837 28868 7871
rect 28816 7828 28868 7837
rect 29184 7871 29236 7880
rect 29184 7837 29193 7871
rect 29193 7837 29227 7871
rect 29227 7837 29236 7871
rect 29184 7828 29236 7837
rect 29644 7828 29696 7880
rect 28080 7803 28132 7812
rect 28080 7769 28089 7803
rect 28089 7769 28123 7803
rect 28123 7769 28132 7803
rect 28080 7760 28132 7769
rect 29828 7871 29880 7880
rect 29828 7837 29837 7871
rect 29837 7837 29871 7871
rect 29871 7837 29880 7871
rect 29828 7828 29880 7837
rect 30288 7828 30340 7880
rect 31392 7905 31401 7939
rect 31401 7905 31435 7939
rect 31435 7905 31444 7939
rect 31392 7896 31444 7905
rect 31484 7939 31536 7948
rect 31484 7905 31493 7939
rect 31493 7905 31527 7939
rect 31527 7905 31536 7939
rect 31484 7896 31536 7905
rect 31024 7828 31076 7880
rect 32312 7896 32364 7948
rect 33048 7896 33100 7948
rect 33416 7896 33468 7948
rect 33508 7939 33560 7948
rect 33508 7905 33517 7939
rect 33517 7905 33551 7939
rect 33551 7905 33560 7939
rect 33508 7896 33560 7905
rect 34796 7896 34848 7948
rect 33784 7828 33836 7880
rect 34704 7828 34756 7880
rect 35992 7964 36044 8016
rect 35440 7896 35492 7948
rect 38200 7896 38252 7948
rect 28264 7735 28316 7744
rect 28264 7701 28289 7735
rect 28289 7701 28316 7735
rect 28264 7692 28316 7701
rect 30840 7692 30892 7744
rect 31300 7692 31352 7744
rect 33324 7760 33376 7812
rect 32312 7692 32364 7744
rect 33968 7692 34020 7744
rect 34520 7760 34572 7812
rect 36084 7828 36136 7880
rect 40040 7828 40092 7880
rect 34612 7692 34664 7744
rect 35072 7692 35124 7744
rect 36360 7692 36412 7744
rect 37004 7803 37056 7812
rect 37004 7769 37013 7803
rect 37013 7769 37047 7803
rect 37047 7769 37056 7803
rect 37004 7760 37056 7769
rect 37464 7760 37516 7812
rect 37280 7692 37332 7744
rect 39028 7692 39080 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 7288 7488 7340 7540
rect 8668 7488 8720 7540
rect 8208 7395 8260 7404
rect 8208 7361 8217 7395
rect 8217 7361 8251 7395
rect 8251 7361 8260 7395
rect 8208 7352 8260 7361
rect 8300 7395 8352 7404
rect 8300 7361 8309 7395
rect 8309 7361 8343 7395
rect 8343 7361 8352 7395
rect 8300 7352 8352 7361
rect 12072 7531 12124 7540
rect 12072 7497 12081 7531
rect 12081 7497 12115 7531
rect 12115 7497 12124 7531
rect 12072 7488 12124 7497
rect 12348 7488 12400 7540
rect 12440 7488 12492 7540
rect 14280 7488 14332 7540
rect 14556 7488 14608 7540
rect 9496 7463 9548 7472
rect 9496 7429 9505 7463
rect 9505 7429 9539 7463
rect 9539 7429 9548 7463
rect 9496 7420 9548 7429
rect 10968 7420 11020 7472
rect 10600 7352 10652 7404
rect 4712 7284 4764 7336
rect 10692 7284 10744 7336
rect 12624 7352 12676 7404
rect 14372 7420 14424 7472
rect 15292 7395 15344 7404
rect 15292 7361 15301 7395
rect 15301 7361 15335 7395
rect 15335 7361 15344 7395
rect 15292 7352 15344 7361
rect 15936 7488 15988 7540
rect 17592 7488 17644 7540
rect 17960 7531 18012 7540
rect 17960 7497 17969 7531
rect 17969 7497 18003 7531
rect 18003 7497 18012 7531
rect 17960 7488 18012 7497
rect 20444 7488 20496 7540
rect 21272 7488 21324 7540
rect 16488 7463 16540 7472
rect 16488 7429 16497 7463
rect 16497 7429 16531 7463
rect 16531 7429 16540 7463
rect 16488 7420 16540 7429
rect 17776 7420 17828 7472
rect 16304 7352 16356 7404
rect 16764 7352 16816 7404
rect 17224 7352 17276 7404
rect 18236 7352 18288 7404
rect 18972 7420 19024 7472
rect 20812 7420 20864 7472
rect 22008 7531 22060 7540
rect 22008 7497 22017 7531
rect 22017 7497 22051 7531
rect 22051 7497 22060 7531
rect 22008 7488 22060 7497
rect 22192 7531 22244 7540
rect 22192 7497 22219 7531
rect 22219 7497 22244 7531
rect 22192 7488 22244 7497
rect 18788 7352 18840 7404
rect 20720 7352 20772 7404
rect 12532 7284 12584 7336
rect 12992 7327 13044 7336
rect 12992 7293 13001 7327
rect 13001 7293 13035 7327
rect 13035 7293 13044 7327
rect 12992 7284 13044 7293
rect 14004 7284 14056 7336
rect 14648 7284 14700 7336
rect 14188 7148 14240 7200
rect 14556 7191 14608 7200
rect 14556 7157 14565 7191
rect 14565 7157 14599 7191
rect 14599 7157 14608 7191
rect 14556 7148 14608 7157
rect 14740 7148 14792 7200
rect 15936 7284 15988 7336
rect 16580 7284 16632 7336
rect 16672 7216 16724 7268
rect 17684 7216 17736 7268
rect 20904 7327 20956 7336
rect 20904 7293 20913 7327
rect 20913 7293 20947 7327
rect 20947 7293 20956 7327
rect 20904 7284 20956 7293
rect 21088 7395 21140 7404
rect 21088 7361 21097 7395
rect 21097 7361 21131 7395
rect 21131 7361 21140 7395
rect 21088 7352 21140 7361
rect 22376 7463 22428 7472
rect 22376 7429 22385 7463
rect 22385 7429 22419 7463
rect 22419 7429 22428 7463
rect 22376 7420 22428 7429
rect 24768 7488 24820 7540
rect 25044 7531 25096 7540
rect 25044 7497 25053 7531
rect 25053 7497 25087 7531
rect 25087 7497 25096 7531
rect 25044 7488 25096 7497
rect 26332 7488 26384 7540
rect 29368 7488 29420 7540
rect 30196 7488 30248 7540
rect 30288 7488 30340 7540
rect 33416 7488 33468 7540
rect 34704 7488 34756 7540
rect 37740 7488 37792 7540
rect 39948 7488 40000 7540
rect 29552 7463 29604 7472
rect 29552 7429 29561 7463
rect 29561 7429 29595 7463
rect 29595 7429 29604 7463
rect 29552 7420 29604 7429
rect 31392 7420 31444 7472
rect 21272 7284 21324 7336
rect 23296 7352 23348 7404
rect 24308 7352 24360 7404
rect 24492 7352 24544 7404
rect 26516 7395 26568 7404
rect 26516 7361 26525 7395
rect 26525 7361 26559 7395
rect 26559 7361 26568 7395
rect 26516 7352 26568 7361
rect 26608 7395 26660 7404
rect 26608 7361 26617 7395
rect 26617 7361 26651 7395
rect 26651 7361 26660 7395
rect 26608 7352 26660 7361
rect 27068 7352 27120 7404
rect 24400 7216 24452 7268
rect 25320 7327 25372 7336
rect 25320 7293 25329 7327
rect 25329 7293 25363 7327
rect 25363 7293 25372 7327
rect 25320 7284 25372 7293
rect 27436 7352 27488 7404
rect 27620 7352 27672 7404
rect 29184 7352 29236 7404
rect 30656 7352 30708 7404
rect 31024 7352 31076 7404
rect 32404 7352 32456 7404
rect 33784 7395 33836 7404
rect 33784 7361 33793 7395
rect 33793 7361 33827 7395
rect 33827 7361 33836 7395
rect 33784 7352 33836 7361
rect 33968 7395 34020 7404
rect 33968 7361 33977 7395
rect 33977 7361 34011 7395
rect 34011 7361 34020 7395
rect 33968 7352 34020 7361
rect 34336 7395 34388 7404
rect 34336 7361 34345 7395
rect 34345 7361 34379 7395
rect 34379 7361 34388 7395
rect 34336 7352 34388 7361
rect 34612 7352 34664 7404
rect 27068 7216 27120 7268
rect 27252 7284 27304 7336
rect 31300 7284 31352 7336
rect 31576 7327 31628 7336
rect 31576 7293 31585 7327
rect 31585 7293 31619 7327
rect 31619 7293 31628 7327
rect 31576 7284 31628 7293
rect 31668 7284 31720 7336
rect 32312 7327 32364 7336
rect 32312 7293 32330 7327
rect 32330 7293 32364 7327
rect 32312 7284 32364 7293
rect 34060 7284 34112 7336
rect 35072 7352 35124 7404
rect 35440 7395 35492 7404
rect 35440 7361 35449 7395
rect 35449 7361 35483 7395
rect 35483 7361 35492 7395
rect 35440 7352 35492 7361
rect 35992 7352 36044 7404
rect 37280 7395 37332 7404
rect 37280 7361 37289 7395
rect 37289 7361 37323 7395
rect 37323 7361 37332 7395
rect 37280 7352 37332 7361
rect 38476 7420 38528 7472
rect 38660 7420 38712 7472
rect 39028 7420 39080 7472
rect 27804 7216 27856 7268
rect 28264 7216 28316 7268
rect 15568 7148 15620 7200
rect 17316 7191 17368 7200
rect 17316 7157 17325 7191
rect 17325 7157 17359 7191
rect 17359 7157 17368 7191
rect 17316 7148 17368 7157
rect 18144 7191 18196 7200
rect 18144 7157 18153 7191
rect 18153 7157 18187 7191
rect 18187 7157 18196 7191
rect 18144 7148 18196 7157
rect 18420 7191 18472 7200
rect 18420 7157 18429 7191
rect 18429 7157 18463 7191
rect 18463 7157 18472 7191
rect 18420 7148 18472 7157
rect 19340 7148 19392 7200
rect 20720 7148 20772 7200
rect 21456 7191 21508 7200
rect 21456 7157 21465 7191
rect 21465 7157 21499 7191
rect 21499 7157 21508 7191
rect 21456 7148 21508 7157
rect 22560 7148 22612 7200
rect 25504 7148 25556 7200
rect 27988 7148 28040 7200
rect 28816 7148 28868 7200
rect 31208 7148 31260 7200
rect 31300 7148 31352 7200
rect 35072 7216 35124 7268
rect 35348 7284 35400 7336
rect 35532 7284 35584 7336
rect 37464 7148 37516 7200
rect 39028 7148 39080 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 12716 6944 12768 6996
rect 12992 6944 13044 6996
rect 12900 6808 12952 6860
rect 13820 6808 13872 6860
rect 14188 6919 14240 6928
rect 14188 6885 14197 6919
rect 14197 6885 14231 6919
rect 14231 6885 14240 6919
rect 14188 6876 14240 6885
rect 14372 6876 14424 6928
rect 15384 6876 15436 6928
rect 15108 6808 15160 6860
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 11520 6740 11572 6749
rect 11796 6783 11848 6792
rect 11796 6749 11805 6783
rect 11805 6749 11839 6783
rect 11839 6749 11848 6783
rect 11796 6740 11848 6749
rect 11980 6740 12032 6792
rect 12256 6740 12308 6792
rect 12532 6740 12584 6792
rect 13636 6783 13688 6792
rect 13636 6749 13645 6783
rect 13645 6749 13679 6783
rect 13679 6749 13688 6783
rect 13636 6740 13688 6749
rect 14556 6740 14608 6792
rect 15292 6740 15344 6792
rect 15568 6808 15620 6860
rect 16580 6808 16632 6860
rect 17132 6944 17184 6996
rect 20536 6944 20588 6996
rect 20628 6944 20680 6996
rect 24216 6944 24268 6996
rect 33876 6944 33928 6996
rect 19616 6876 19668 6928
rect 21456 6876 21508 6928
rect 22284 6876 22336 6928
rect 28264 6876 28316 6928
rect 35532 6944 35584 6996
rect 36360 6987 36412 6996
rect 36360 6953 36369 6987
rect 36369 6953 36403 6987
rect 36403 6953 36412 6987
rect 36360 6944 36412 6953
rect 37280 6944 37332 6996
rect 37372 6944 37424 6996
rect 18880 6808 18932 6860
rect 24952 6808 25004 6860
rect 25964 6808 26016 6860
rect 29000 6808 29052 6860
rect 20536 6740 20588 6792
rect 29276 6740 29328 6792
rect 29920 6783 29972 6792
rect 29920 6749 29929 6783
rect 29929 6749 29963 6783
rect 29963 6749 29972 6783
rect 29920 6740 29972 6749
rect 11888 6715 11940 6724
rect 11888 6681 11897 6715
rect 11897 6681 11931 6715
rect 11931 6681 11940 6715
rect 11888 6672 11940 6681
rect 15936 6672 15988 6724
rect 18604 6672 18656 6724
rect 21548 6672 21600 6724
rect 29460 6672 29512 6724
rect 33600 6808 33652 6860
rect 30196 6783 30248 6792
rect 30196 6749 30205 6783
rect 30205 6749 30239 6783
rect 30239 6749 30248 6783
rect 30196 6740 30248 6749
rect 33692 6740 33744 6792
rect 37464 6808 37516 6860
rect 38200 6808 38252 6860
rect 15016 6604 15068 6656
rect 16672 6604 16724 6656
rect 16764 6647 16816 6656
rect 16764 6613 16773 6647
rect 16773 6613 16807 6647
rect 16807 6613 16816 6647
rect 16764 6604 16816 6613
rect 17132 6647 17184 6656
rect 17132 6613 17141 6647
rect 17141 6613 17175 6647
rect 17175 6613 17184 6647
rect 17132 6604 17184 6613
rect 25320 6604 25372 6656
rect 28080 6604 28132 6656
rect 30104 6647 30156 6656
rect 30104 6613 30113 6647
rect 30113 6613 30147 6647
rect 30147 6613 30156 6647
rect 30104 6604 30156 6613
rect 30196 6604 30248 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 11888 6443 11940 6452
rect 11888 6409 11897 6443
rect 11897 6409 11931 6443
rect 11931 6409 11940 6443
rect 11888 6400 11940 6409
rect 13636 6400 13688 6452
rect 15108 6400 15160 6452
rect 16396 6443 16448 6452
rect 16396 6409 16405 6443
rect 16405 6409 16439 6443
rect 16439 6409 16448 6443
rect 16396 6400 16448 6409
rect 17132 6400 17184 6452
rect 19064 6400 19116 6452
rect 21272 6400 21324 6452
rect 24492 6400 24544 6452
rect 26516 6400 26568 6452
rect 26884 6400 26936 6452
rect 29184 6400 29236 6452
rect 29552 6400 29604 6452
rect 30104 6400 30156 6452
rect 15200 6332 15252 6384
rect 15384 6332 15436 6384
rect 16856 6332 16908 6384
rect 17684 6332 17736 6384
rect 19340 6375 19392 6384
rect 19340 6341 19349 6375
rect 19349 6341 19383 6375
rect 19383 6341 19392 6375
rect 19340 6332 19392 6341
rect 20260 6332 20312 6384
rect 22376 6332 22428 6384
rect 26240 6332 26292 6384
rect 24952 6307 25004 6316
rect 24952 6273 24961 6307
rect 24961 6273 24995 6307
rect 24995 6273 25004 6307
rect 24952 6264 25004 6273
rect 12256 6196 12308 6248
rect 16764 6196 16816 6248
rect 17224 6196 17276 6248
rect 20444 6196 20496 6248
rect 23020 6196 23072 6248
rect 23756 6196 23808 6248
rect 25412 6264 25464 6316
rect 26792 6307 26844 6316
rect 26792 6273 26801 6307
rect 26801 6273 26835 6307
rect 26835 6273 26844 6307
rect 26792 6264 26844 6273
rect 26884 6264 26936 6316
rect 26240 6196 26292 6248
rect 27344 6307 27396 6316
rect 27344 6273 27353 6307
rect 27353 6273 27387 6307
rect 27387 6273 27396 6307
rect 27344 6264 27396 6273
rect 12992 6128 13044 6180
rect 15936 6128 15988 6180
rect 22284 6128 22336 6180
rect 25596 6128 25648 6180
rect 29368 6332 29420 6384
rect 30196 6332 30248 6384
rect 28724 6264 28776 6316
rect 31300 6264 31352 6316
rect 31668 6264 31720 6316
rect 10692 6060 10744 6112
rect 16212 6060 16264 6112
rect 17960 6060 18012 6112
rect 19524 6060 19576 6112
rect 21272 6060 21324 6112
rect 22192 6060 22244 6112
rect 22376 6103 22428 6112
rect 22376 6069 22385 6103
rect 22385 6069 22419 6103
rect 22419 6069 22428 6103
rect 22376 6060 22428 6069
rect 23572 6060 23624 6112
rect 24768 6060 24820 6112
rect 25136 6103 25188 6112
rect 25136 6069 25145 6103
rect 25145 6069 25179 6103
rect 25179 6069 25188 6103
rect 25136 6060 25188 6069
rect 27252 6060 27304 6112
rect 27344 6060 27396 6112
rect 29460 6060 29512 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 18788 5856 18840 5908
rect 19340 5788 19392 5840
rect 19984 5899 20036 5908
rect 19984 5865 19993 5899
rect 19993 5865 20027 5899
rect 20027 5865 20036 5899
rect 19984 5856 20036 5865
rect 20444 5899 20496 5908
rect 20444 5865 20453 5899
rect 20453 5865 20487 5899
rect 20487 5865 20496 5899
rect 20444 5856 20496 5865
rect 21548 5856 21600 5908
rect 10784 5720 10836 5772
rect 18604 5720 18656 5772
rect 18696 5720 18748 5772
rect 18512 5695 18564 5704
rect 18512 5661 18521 5695
rect 18521 5661 18555 5695
rect 18555 5661 18564 5695
rect 18512 5652 18564 5661
rect 18788 5695 18840 5704
rect 18788 5661 18797 5695
rect 18797 5661 18831 5695
rect 18831 5661 18840 5695
rect 18788 5652 18840 5661
rect 19156 5652 19208 5704
rect 19432 5652 19484 5704
rect 19524 5695 19576 5704
rect 19524 5661 19533 5695
rect 19533 5661 19567 5695
rect 19567 5661 19576 5695
rect 19524 5652 19576 5661
rect 10692 5627 10744 5636
rect 10692 5593 10701 5627
rect 10701 5593 10735 5627
rect 10735 5593 10744 5627
rect 10692 5584 10744 5593
rect 10600 5516 10652 5568
rect 18144 5584 18196 5636
rect 11336 5516 11388 5568
rect 12256 5516 12308 5568
rect 17040 5559 17092 5568
rect 17040 5525 17049 5559
rect 17049 5525 17083 5559
rect 17083 5525 17092 5559
rect 17040 5516 17092 5525
rect 19248 5516 19300 5568
rect 19892 5652 19944 5704
rect 20076 5695 20128 5704
rect 20076 5661 20085 5695
rect 20085 5661 20119 5695
rect 20119 5661 20128 5695
rect 20076 5652 20128 5661
rect 20720 5788 20772 5840
rect 21364 5788 21416 5840
rect 20536 5695 20588 5704
rect 20536 5661 20545 5695
rect 20545 5661 20579 5695
rect 20579 5661 20588 5695
rect 20536 5652 20588 5661
rect 21272 5652 21324 5704
rect 21548 5695 21600 5704
rect 21548 5661 21557 5695
rect 21557 5661 21591 5695
rect 21591 5661 21600 5695
rect 21548 5652 21600 5661
rect 21732 5652 21784 5704
rect 23204 5720 23256 5772
rect 24216 5763 24268 5772
rect 24216 5729 24225 5763
rect 24225 5729 24259 5763
rect 24259 5729 24268 5763
rect 24216 5720 24268 5729
rect 22100 5652 22152 5704
rect 24492 5695 24544 5704
rect 24492 5661 24501 5695
rect 24501 5661 24535 5695
rect 24535 5661 24544 5695
rect 24492 5652 24544 5661
rect 24860 5788 24912 5840
rect 24952 5788 25004 5840
rect 25504 5856 25556 5908
rect 26424 5856 26476 5908
rect 25412 5788 25464 5840
rect 26700 5788 26752 5840
rect 27252 5763 27304 5772
rect 27252 5729 27261 5763
rect 27261 5729 27295 5763
rect 27295 5729 27304 5763
rect 27252 5720 27304 5729
rect 25136 5652 25188 5704
rect 22192 5584 22244 5636
rect 22468 5627 22520 5636
rect 22468 5593 22477 5627
rect 22477 5593 22511 5627
rect 22511 5593 22520 5627
rect 22468 5584 22520 5593
rect 24584 5584 24636 5636
rect 21732 5516 21784 5568
rect 22376 5516 22428 5568
rect 24768 5627 24820 5636
rect 24768 5593 24777 5627
rect 24777 5593 24811 5627
rect 24811 5593 24820 5627
rect 24768 5584 24820 5593
rect 24952 5516 25004 5568
rect 25044 5559 25096 5568
rect 25044 5525 25053 5559
rect 25053 5525 25087 5559
rect 25087 5525 25096 5559
rect 25044 5516 25096 5525
rect 25136 5559 25188 5568
rect 25136 5525 25145 5559
rect 25145 5525 25179 5559
rect 25179 5525 25188 5559
rect 25136 5516 25188 5525
rect 25412 5627 25464 5636
rect 25412 5593 25421 5627
rect 25421 5593 25455 5627
rect 25455 5593 25464 5627
rect 25412 5584 25464 5593
rect 25504 5627 25556 5636
rect 25504 5593 25513 5627
rect 25513 5593 25547 5627
rect 25547 5593 25556 5627
rect 25504 5584 25556 5593
rect 25688 5695 25740 5704
rect 25688 5661 25697 5695
rect 25697 5661 25731 5695
rect 25731 5661 25740 5695
rect 25688 5652 25740 5661
rect 25780 5695 25832 5704
rect 25780 5661 25789 5695
rect 25789 5661 25823 5695
rect 25823 5661 25832 5695
rect 25780 5652 25832 5661
rect 26240 5695 26292 5704
rect 26240 5661 26249 5695
rect 26249 5661 26283 5695
rect 26283 5661 26292 5695
rect 26240 5652 26292 5661
rect 26884 5652 26936 5704
rect 28724 5899 28776 5908
rect 28724 5865 28733 5899
rect 28733 5865 28767 5899
rect 28767 5865 28776 5899
rect 28724 5856 28776 5865
rect 29552 5899 29604 5908
rect 29552 5865 29561 5899
rect 29561 5865 29595 5899
rect 29595 5865 29604 5899
rect 29552 5856 29604 5865
rect 31300 5763 31352 5772
rect 31300 5729 31309 5763
rect 31309 5729 31343 5763
rect 31343 5729 31352 5763
rect 31300 5720 31352 5729
rect 29184 5695 29236 5704
rect 29184 5661 29193 5695
rect 29193 5661 29227 5695
rect 29227 5661 29236 5695
rect 29184 5652 29236 5661
rect 26424 5627 26476 5636
rect 26424 5593 26433 5627
rect 26433 5593 26467 5627
rect 26467 5593 26476 5627
rect 26424 5584 26476 5593
rect 26516 5627 26568 5636
rect 26516 5593 26525 5627
rect 26525 5593 26559 5627
rect 26559 5593 26568 5627
rect 26516 5584 26568 5593
rect 25688 5516 25740 5568
rect 25964 5559 26016 5568
rect 25964 5525 25973 5559
rect 25973 5525 26007 5559
rect 26007 5525 26016 5559
rect 25964 5516 26016 5525
rect 27344 5584 27396 5636
rect 28080 5516 28132 5568
rect 29460 5584 29512 5636
rect 30288 5584 30340 5636
rect 29092 5516 29144 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 13820 5312 13872 5364
rect 13360 5244 13412 5296
rect 18512 5312 18564 5364
rect 21364 5355 21416 5364
rect 21364 5321 21373 5355
rect 21373 5321 21407 5355
rect 21407 5321 21416 5355
rect 21364 5312 21416 5321
rect 22284 5312 22336 5364
rect 22468 5312 22520 5364
rect 25780 5312 25832 5364
rect 26792 5312 26844 5364
rect 15384 5244 15436 5296
rect 17040 5244 17092 5296
rect 17684 5244 17736 5296
rect 10968 5176 11020 5228
rect 20076 5244 20128 5296
rect 18604 5176 18656 5228
rect 19340 5219 19392 5228
rect 19340 5185 19349 5219
rect 19349 5185 19383 5219
rect 19383 5185 19392 5219
rect 19340 5176 19392 5185
rect 20628 5176 20680 5228
rect 22376 5244 22428 5296
rect 12072 5151 12124 5160
rect 12072 5117 12081 5151
rect 12081 5117 12115 5151
rect 12115 5117 12124 5151
rect 12072 5108 12124 5117
rect 14280 5108 14332 5160
rect 14924 5040 14976 5092
rect 15200 4972 15252 5024
rect 15384 5015 15436 5024
rect 15384 4981 15393 5015
rect 15393 4981 15427 5015
rect 15427 4981 15436 5015
rect 17040 5108 17092 5160
rect 17500 5108 17552 5160
rect 18972 5108 19024 5160
rect 19340 5040 19392 5092
rect 20076 5040 20128 5092
rect 21456 5219 21508 5228
rect 21456 5185 21465 5219
rect 21465 5185 21499 5219
rect 21499 5185 21508 5219
rect 21456 5176 21508 5185
rect 22100 5176 22152 5228
rect 23020 5176 23072 5228
rect 24216 5244 24268 5296
rect 22376 5151 22428 5160
rect 22376 5117 22385 5151
rect 22385 5117 22419 5151
rect 22419 5117 22428 5151
rect 22376 5108 22428 5117
rect 22836 5040 22888 5092
rect 23940 5176 23992 5228
rect 24860 5244 24912 5296
rect 25044 5244 25096 5296
rect 29092 5312 29144 5364
rect 30288 5355 30340 5364
rect 30288 5321 30297 5355
rect 30297 5321 30331 5355
rect 30331 5321 30340 5355
rect 30288 5312 30340 5321
rect 28172 5244 28224 5296
rect 31300 5244 31352 5296
rect 29000 5219 29052 5228
rect 29000 5185 29009 5219
rect 29009 5185 29043 5219
rect 29043 5185 29052 5219
rect 29000 5176 29052 5185
rect 29184 5219 29236 5228
rect 29184 5185 29193 5219
rect 29193 5185 29227 5219
rect 29227 5185 29236 5219
rect 29184 5176 29236 5185
rect 30196 5219 30248 5228
rect 30196 5185 30205 5219
rect 30205 5185 30239 5219
rect 30239 5185 30248 5219
rect 30196 5176 30248 5185
rect 25688 5108 25740 5160
rect 26148 5108 26200 5160
rect 28080 5108 28132 5160
rect 15384 4972 15436 4981
rect 18144 4972 18196 5024
rect 19524 4972 19576 5024
rect 20628 4972 20680 5024
rect 20904 5015 20956 5024
rect 20904 4981 20913 5015
rect 20913 4981 20947 5015
rect 20947 4981 20956 5015
rect 20904 4972 20956 4981
rect 21272 4972 21324 5024
rect 28632 4972 28684 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 12072 4768 12124 4820
rect 14280 4811 14332 4820
rect 14280 4777 14289 4811
rect 14289 4777 14323 4811
rect 14323 4777 14332 4811
rect 14280 4768 14332 4777
rect 13912 4700 13964 4752
rect 18972 4768 19024 4820
rect 19708 4768 19760 4820
rect 20536 4768 20588 4820
rect 21456 4768 21508 4820
rect 12992 4675 13044 4684
rect 12992 4641 13001 4675
rect 13001 4641 13035 4675
rect 13035 4641 13044 4675
rect 12992 4632 13044 4641
rect 14924 4700 14976 4752
rect 20628 4700 20680 4752
rect 15016 4632 15068 4684
rect 15200 4632 15252 4684
rect 16580 4632 16632 4684
rect 12256 4607 12308 4616
rect 12256 4573 12265 4607
rect 12265 4573 12299 4607
rect 12299 4573 12308 4607
rect 12256 4564 12308 4573
rect 12348 4564 12400 4616
rect 13820 4607 13872 4616
rect 13820 4573 13829 4607
rect 13829 4573 13863 4607
rect 13863 4573 13872 4607
rect 13820 4564 13872 4573
rect 14280 4564 14332 4616
rect 17224 4564 17276 4616
rect 19524 4675 19576 4684
rect 19524 4641 19533 4675
rect 19533 4641 19567 4675
rect 19567 4641 19576 4675
rect 19524 4632 19576 4641
rect 20076 4632 20128 4684
rect 23112 4632 23164 4684
rect 24768 4675 24820 4684
rect 24768 4641 24777 4675
rect 24777 4641 24811 4675
rect 24811 4641 24820 4675
rect 24768 4632 24820 4641
rect 39948 4632 40000 4684
rect 26148 4564 26200 4616
rect 26700 4564 26752 4616
rect 14188 4496 14240 4548
rect 15200 4496 15252 4548
rect 15476 4496 15528 4548
rect 16028 4496 16080 4548
rect 11612 4471 11664 4480
rect 11612 4437 11621 4471
rect 11621 4437 11655 4471
rect 11655 4437 11664 4471
rect 11612 4428 11664 4437
rect 16856 4428 16908 4480
rect 17684 4496 17736 4548
rect 20168 4496 20220 4548
rect 21640 4496 21692 4548
rect 22652 4539 22704 4548
rect 22652 4505 22661 4539
rect 22661 4505 22695 4539
rect 22695 4505 22704 4539
rect 22652 4496 22704 4505
rect 25136 4496 25188 4548
rect 18328 4428 18380 4480
rect 24768 4428 24820 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 11612 4224 11664 4276
rect 12716 4267 12768 4276
rect 12716 4233 12725 4267
rect 12725 4233 12759 4267
rect 12759 4233 12768 4267
rect 12716 4224 12768 4233
rect 16028 4224 16080 4276
rect 17960 4224 18012 4276
rect 11888 4199 11940 4208
rect 11888 4165 11897 4199
rect 11897 4165 11931 4199
rect 11931 4165 11940 4199
rect 11888 4156 11940 4165
rect 16948 4156 17000 4208
rect 17684 4156 17736 4208
rect 16672 4131 16724 4140
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 19340 4156 19392 4208
rect 20168 4156 20220 4208
rect 20904 4224 20956 4276
rect 21272 4199 21324 4208
rect 21272 4165 21281 4199
rect 21281 4165 21315 4199
rect 21315 4165 21324 4199
rect 21272 4156 21324 4165
rect 22652 4267 22704 4276
rect 22652 4233 22661 4267
rect 22661 4233 22695 4267
rect 22695 4233 22704 4267
rect 22652 4224 22704 4233
rect 23020 4224 23072 4276
rect 29184 4224 29236 4276
rect 21456 4156 21508 4208
rect 18696 4131 18748 4140
rect 18696 4097 18705 4131
rect 18705 4097 18739 4131
rect 18739 4097 18748 4131
rect 18696 4088 18748 4097
rect 18880 4088 18932 4140
rect 19708 4131 19760 4140
rect 19708 4097 19717 4131
rect 19717 4097 19751 4131
rect 19751 4097 19760 4131
rect 19708 4088 19760 4097
rect 19892 4088 19944 4140
rect 20076 4131 20128 4140
rect 20076 4097 20085 4131
rect 20085 4097 20119 4131
rect 20119 4097 20128 4131
rect 20076 4088 20128 4097
rect 12992 4063 13044 4072
rect 12992 4029 13001 4063
rect 13001 4029 13035 4063
rect 13035 4029 13044 4063
rect 12992 4020 13044 4029
rect 13820 4020 13872 4072
rect 14004 4020 14056 4072
rect 15660 4020 15712 4072
rect 16856 4020 16908 4072
rect 18328 4063 18380 4072
rect 18328 4029 18337 4063
rect 18337 4029 18371 4063
rect 18371 4029 18380 4063
rect 18328 4020 18380 4029
rect 18604 4063 18656 4072
rect 18604 4029 18613 4063
rect 18613 4029 18647 4063
rect 18647 4029 18656 4063
rect 18604 4020 18656 4029
rect 15016 3952 15068 4004
rect 19432 3952 19484 4004
rect 11060 3884 11112 3936
rect 11888 3884 11940 3936
rect 12992 3884 13044 3936
rect 14832 3884 14884 3936
rect 17040 3884 17092 3936
rect 17132 3927 17184 3936
rect 17132 3893 17141 3927
rect 17141 3893 17175 3927
rect 17175 3893 17184 3927
rect 17132 3884 17184 3893
rect 18788 3884 18840 3936
rect 23940 4156 23992 4208
rect 30196 4156 30248 4208
rect 20720 4088 20772 4140
rect 21548 4131 21600 4140
rect 21548 4097 21557 4131
rect 21557 4097 21591 4131
rect 21591 4097 21600 4131
rect 21548 4088 21600 4097
rect 21732 4088 21784 4140
rect 21824 4088 21876 4140
rect 21180 4020 21232 4072
rect 23020 4088 23072 4140
rect 23296 4131 23348 4140
rect 23296 4097 23305 4131
rect 23305 4097 23339 4131
rect 23339 4097 23348 4131
rect 23296 4088 23348 4097
rect 23480 4131 23532 4140
rect 23480 4097 23489 4131
rect 23489 4097 23523 4131
rect 23523 4097 23532 4131
rect 23480 4088 23532 4097
rect 28172 4131 28224 4140
rect 28172 4097 28181 4131
rect 28181 4097 28215 4131
rect 28215 4097 28224 4131
rect 28172 4088 28224 4097
rect 28632 4088 28684 4140
rect 23388 4020 23440 4072
rect 29276 3952 29328 4004
rect 22376 3884 22428 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 11612 3680 11664 3732
rect 12256 3680 12308 3732
rect 20076 3680 20128 3732
rect 21548 3680 21600 3732
rect 10968 3544 11020 3596
rect 12992 3587 13044 3596
rect 12992 3553 13001 3587
rect 13001 3553 13035 3587
rect 13035 3553 13044 3587
rect 12992 3544 13044 3553
rect 13084 3544 13136 3596
rect 14832 3587 14884 3596
rect 14832 3553 14841 3587
rect 14841 3553 14875 3587
rect 14875 3553 14884 3587
rect 14832 3544 14884 3553
rect 15016 3587 15068 3596
rect 15016 3553 15025 3587
rect 15025 3553 15059 3587
rect 15059 3553 15068 3587
rect 17868 3612 17920 3664
rect 15016 3544 15068 3553
rect 12900 3519 12952 3528
rect 12900 3485 12909 3519
rect 12909 3485 12943 3519
rect 12943 3485 12952 3519
rect 12900 3476 12952 3485
rect 13912 3476 13964 3528
rect 14648 3476 14700 3528
rect 15568 3519 15620 3528
rect 15568 3485 15577 3519
rect 15577 3485 15611 3519
rect 15611 3485 15620 3519
rect 15568 3476 15620 3485
rect 16948 3476 17000 3528
rect 18788 3476 18840 3528
rect 19248 3519 19300 3528
rect 19248 3485 19257 3519
rect 19257 3485 19291 3519
rect 19291 3485 19300 3519
rect 19248 3476 19300 3485
rect 21364 3519 21416 3528
rect 21364 3485 21373 3519
rect 21373 3485 21407 3519
rect 21407 3485 21416 3519
rect 21364 3476 21416 3485
rect 21640 3476 21692 3528
rect 11060 3408 11112 3460
rect 10600 3340 10652 3392
rect 15752 3408 15804 3460
rect 22928 3680 22980 3732
rect 23296 3680 23348 3732
rect 39948 3655 40000 3664
rect 39948 3621 39957 3655
rect 39957 3621 39991 3655
rect 39991 3621 40000 3655
rect 39948 3612 40000 3621
rect 22744 3544 22796 3596
rect 23112 3544 23164 3596
rect 24860 3544 24912 3596
rect 12532 3383 12584 3392
rect 12532 3349 12541 3383
rect 12541 3349 12575 3383
rect 12575 3349 12584 3383
rect 12532 3340 12584 3349
rect 14096 3340 14148 3392
rect 17408 3383 17460 3392
rect 17408 3349 17417 3383
rect 17417 3349 17451 3383
rect 17451 3349 17460 3383
rect 17408 3340 17460 3349
rect 21548 3340 21600 3392
rect 24768 3476 24820 3528
rect 26792 3519 26844 3528
rect 26792 3485 26801 3519
rect 26801 3485 26835 3519
rect 26835 3485 26844 3519
rect 26792 3476 26844 3485
rect 40132 3451 40184 3460
rect 40132 3417 40141 3451
rect 40141 3417 40175 3451
rect 40175 3417 40184 3451
rect 40132 3408 40184 3417
rect 24216 3383 24268 3392
rect 24216 3349 24225 3383
rect 24225 3349 24259 3383
rect 24259 3349 24268 3383
rect 24216 3340 24268 3349
rect 24308 3340 24360 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 11612 3043 11664 3052
rect 11612 3009 11621 3043
rect 11621 3009 11655 3043
rect 11655 3009 11664 3043
rect 11612 3000 11664 3009
rect 11796 2932 11848 2984
rect 12532 3068 12584 3120
rect 13360 3000 13412 3052
rect 15568 3136 15620 3188
rect 16672 3136 16724 3188
rect 17040 3179 17092 3188
rect 17040 3145 17049 3179
rect 17049 3145 17083 3179
rect 17083 3145 17092 3179
rect 17040 3136 17092 3145
rect 17132 3179 17184 3188
rect 17132 3145 17141 3179
rect 17141 3145 17175 3179
rect 17175 3145 17184 3179
rect 17132 3136 17184 3145
rect 14096 3111 14148 3120
rect 14096 3077 14105 3111
rect 14105 3077 14139 3111
rect 14139 3077 14148 3111
rect 14096 3068 14148 3077
rect 15752 3111 15804 3120
rect 15752 3077 15761 3111
rect 15761 3077 15795 3111
rect 15795 3077 15804 3111
rect 15752 3068 15804 3077
rect 15200 3000 15252 3052
rect 15476 3000 15528 3052
rect 16672 3000 16724 3052
rect 17224 3000 17276 3052
rect 18788 3068 18840 3120
rect 21640 3179 21692 3188
rect 21640 3145 21649 3179
rect 21649 3145 21683 3179
rect 21683 3145 21692 3179
rect 21640 3136 21692 3145
rect 22836 3136 22888 3188
rect 26792 3136 26844 3188
rect 21548 3068 21600 3120
rect 12808 2932 12860 2984
rect 17868 2932 17920 2984
rect 19340 2932 19392 2984
rect 20168 2975 20220 2984
rect 20168 2941 20177 2975
rect 20177 2941 20211 2975
rect 20211 2941 20220 2975
rect 20168 2932 20220 2941
rect 20812 2932 20864 2984
rect 21916 2932 21968 2984
rect 22468 2932 22520 2984
rect 23112 3000 23164 3052
rect 23480 3068 23532 3120
rect 23940 3111 23992 3120
rect 23940 3077 23949 3111
rect 23949 3077 23983 3111
rect 23983 3077 23992 3111
rect 23940 3068 23992 3077
rect 24216 3068 24268 3120
rect 24308 3043 24360 3052
rect 24308 3009 24317 3043
rect 24317 3009 24351 3043
rect 24351 3009 24360 3043
rect 24308 3000 24360 3009
rect 23388 2932 23440 2984
rect 13820 2864 13872 2916
rect 15660 2864 15712 2916
rect 16580 2864 16632 2916
rect 12348 2796 12400 2848
rect 19800 2839 19852 2848
rect 19800 2805 19809 2839
rect 19809 2805 19843 2839
rect 19843 2805 19852 2839
rect 19800 2796 19852 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 19248 2592 19300 2644
rect 19340 2635 19392 2644
rect 19340 2601 19349 2635
rect 19349 2601 19383 2635
rect 19383 2601 19392 2635
rect 19340 2592 19392 2601
rect 20168 2592 20220 2644
rect 12900 2524 12952 2576
rect 13544 2524 13596 2576
rect 11796 2456 11848 2508
rect 11336 2431 11388 2440
rect 11336 2397 11345 2431
rect 11345 2397 11379 2431
rect 11379 2397 11388 2431
rect 11336 2388 11388 2397
rect 14004 2388 14056 2440
rect 14280 2431 14332 2440
rect 14280 2397 14289 2431
rect 14289 2397 14323 2431
rect 14323 2397 14332 2431
rect 14280 2388 14332 2397
rect 15384 2456 15436 2508
rect 16672 2456 16724 2508
rect 17408 2499 17460 2508
rect 17408 2465 17417 2499
rect 17417 2465 17451 2499
rect 17451 2465 17460 2499
rect 17408 2456 17460 2465
rect 19800 2456 19852 2508
rect 11888 2320 11940 2372
rect 12808 2320 12860 2372
rect 13820 2320 13872 2372
rect 15568 2388 15620 2440
rect 16856 2388 16908 2440
rect 19340 2388 19392 2440
rect 20628 2388 20680 2440
rect 22744 2456 22796 2508
rect 23020 2388 23072 2440
rect 17960 2320 18012 2372
rect 20720 2320 20772 2372
rect 22468 2320 22520 2372
rect 11612 2252 11664 2304
rect 14188 2252 14240 2304
rect 14832 2252 14884 2304
rect 16120 2252 16172 2304
rect 16764 2252 16816 2304
rect 21364 2252 21416 2304
rect 23848 2252 23900 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
<< metal2 >>
rect 7102 43101 7158 43901
rect 23846 43101 23902 43901
rect 24490 43101 24546 43901
rect 25134 43101 25190 43901
rect 25778 43101 25834 43901
rect 26422 43101 26478 43901
rect 27066 43101 27122 43901
rect 27710 43101 27766 43901
rect 28354 43101 28410 43901
rect 30930 43101 30986 43901
rect 7116 41414 7144 43101
rect 7024 41386 7144 41414
rect 4874 41372 5182 41381
rect 4874 41370 4880 41372
rect 4936 41370 4960 41372
rect 5016 41370 5040 41372
rect 5096 41370 5120 41372
rect 5176 41370 5182 41372
rect 4936 41318 4938 41370
rect 5118 41318 5120 41370
rect 4874 41316 4880 41318
rect 4936 41316 4960 41318
rect 5016 41316 5040 41318
rect 5096 41316 5120 41318
rect 5176 41316 5182 41318
rect 4874 41307 5182 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4874 40284 5182 40293
rect 4874 40282 4880 40284
rect 4936 40282 4960 40284
rect 5016 40282 5040 40284
rect 5096 40282 5120 40284
rect 5176 40282 5182 40284
rect 4936 40230 4938 40282
rect 5118 40230 5120 40282
rect 4874 40228 4880 40230
rect 4936 40228 4960 40230
rect 5016 40228 5040 40230
rect 5096 40228 5120 40230
rect 5176 40228 5182 40230
rect 4874 40219 5182 40228
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4874 39196 5182 39205
rect 4874 39194 4880 39196
rect 4936 39194 4960 39196
rect 5016 39194 5040 39196
rect 5096 39194 5120 39196
rect 5176 39194 5182 39196
rect 4936 39142 4938 39194
rect 5118 39142 5120 39194
rect 4874 39140 4880 39142
rect 4936 39140 4960 39142
rect 5016 39140 5040 39142
rect 5096 39140 5120 39142
rect 5176 39140 5182 39142
rect 4874 39131 5182 39140
rect 6828 38888 6880 38894
rect 3422 38856 3478 38865
rect 6828 38830 6880 38836
rect 3422 38791 3478 38800
rect 2962 36136 3018 36145
rect 2962 36071 3018 36080
rect 2976 36038 3004 36071
rect 2964 36032 3016 36038
rect 2964 35974 3016 35980
rect 2976 35766 3004 35974
rect 1308 35760 1360 35766
rect 1308 35702 1360 35708
rect 2964 35760 3016 35766
rect 2964 35702 3016 35708
rect 1320 35018 1348 35702
rect 2228 35692 2280 35698
rect 2228 35634 2280 35640
rect 1308 35012 1360 35018
rect 1308 34954 1360 34960
rect 1320 34785 1348 34954
rect 1306 34776 1362 34785
rect 1306 34711 1362 34720
rect 1674 34096 1730 34105
rect 1674 34031 1730 34040
rect 1688 33930 1716 34031
rect 1676 33924 1728 33930
rect 1676 33866 1728 33872
rect 2240 33658 2268 35634
rect 3148 35488 3200 35494
rect 3148 35430 3200 35436
rect 3160 35154 3188 35430
rect 3148 35148 3200 35154
rect 3148 35090 3200 35096
rect 2688 35012 2740 35018
rect 2688 34954 2740 34960
rect 2700 34746 2728 34954
rect 2688 34740 2740 34746
rect 2688 34682 2740 34688
rect 2320 34536 2372 34542
rect 2320 34478 2372 34484
rect 2332 33930 2360 34478
rect 2320 33924 2372 33930
rect 2320 33866 2372 33872
rect 2228 33652 2280 33658
rect 2228 33594 2280 33600
rect 1492 33584 1544 33590
rect 1492 33526 1544 33532
rect 1504 32842 1532 33526
rect 2240 33522 2268 33594
rect 2228 33516 2280 33522
rect 2228 33458 2280 33464
rect 1676 33448 1728 33454
rect 1674 33416 1676 33425
rect 1728 33416 1730 33425
rect 1674 33351 1730 33360
rect 1492 32836 1544 32842
rect 1492 32778 1544 32784
rect 1504 32745 1532 32778
rect 1490 32736 1546 32745
rect 1490 32671 1546 32680
rect 1688 32502 1716 33351
rect 2700 32824 2728 34682
rect 2872 33380 2924 33386
rect 2872 33322 2924 33328
rect 2884 32978 2912 33322
rect 2872 32972 2924 32978
rect 2872 32914 2924 32920
rect 2780 32836 2832 32842
rect 2608 32796 2780 32824
rect 2608 32502 2636 32796
rect 2780 32778 2832 32784
rect 1676 32496 1728 32502
rect 1676 32438 1728 32444
rect 2596 32496 2648 32502
rect 2596 32438 2648 32444
rect 2608 32026 2636 32438
rect 2596 32020 2648 32026
rect 2596 31962 2648 31968
rect 2608 31754 2636 31962
rect 2608 31726 2728 31754
rect 2700 31414 2728 31726
rect 2872 31476 2924 31482
rect 2872 31418 2924 31424
rect 2688 31408 2740 31414
rect 2688 31350 2740 31356
rect 1582 30696 1638 30705
rect 2700 30666 2728 31350
rect 1582 30631 1584 30640
rect 1636 30631 1638 30640
rect 2688 30660 2740 30666
rect 1584 30602 1636 30608
rect 2688 30602 2740 30608
rect 1596 30394 1624 30602
rect 1584 30388 1636 30394
rect 1584 30330 1636 30336
rect 2884 30258 2912 31418
rect 3238 31376 3294 31385
rect 3238 31311 3294 31320
rect 3252 31278 3280 31311
rect 3240 31272 3292 31278
rect 3240 31214 3292 31220
rect 3252 30802 3280 31214
rect 3240 30796 3292 30802
rect 3240 30738 3292 30744
rect 3332 30660 3384 30666
rect 3332 30602 3384 30608
rect 3344 30326 3372 30602
rect 3332 30320 3384 30326
rect 3332 30262 3384 30268
rect 848 30252 900 30258
rect 848 30194 900 30200
rect 2872 30252 2924 30258
rect 2872 30194 2924 30200
rect 860 30161 888 30194
rect 846 30152 902 30161
rect 846 30087 902 30096
rect 3148 27056 3200 27062
rect 3148 26998 3200 27004
rect 3056 26580 3108 26586
rect 3056 26522 3108 26528
rect 2780 26444 2832 26450
rect 2780 26386 2832 26392
rect 1860 26240 1912 26246
rect 1860 26182 1912 26188
rect 1872 25974 1900 26182
rect 1860 25968 1912 25974
rect 1860 25910 1912 25916
rect 1584 25832 1636 25838
rect 1584 25774 1636 25780
rect 1596 25362 1624 25774
rect 1584 25356 1636 25362
rect 1584 25298 1636 25304
rect 1860 25220 1912 25226
rect 1860 25162 1912 25168
rect 1872 24954 1900 25162
rect 1860 24948 1912 24954
rect 1860 24890 1912 24896
rect 1676 24132 1728 24138
rect 1676 24074 1728 24080
rect 1688 23866 1716 24074
rect 1676 23860 1728 23866
rect 1676 23802 1728 23808
rect 2596 22976 2648 22982
rect 2596 22918 2648 22924
rect 2608 22778 2636 22918
rect 2596 22772 2648 22778
rect 2596 22714 2648 22720
rect 2228 22432 2280 22438
rect 2228 22374 2280 22380
rect 2240 22234 2268 22374
rect 2228 22228 2280 22234
rect 2228 22170 2280 22176
rect 2792 22114 2820 26386
rect 2872 25356 2924 25362
rect 2872 25298 2924 25304
rect 2884 24274 2912 25298
rect 2964 24608 3016 24614
rect 2964 24550 3016 24556
rect 2872 24268 2924 24274
rect 2872 24210 2924 24216
rect 2884 23118 2912 24210
rect 2976 23866 3004 24550
rect 2964 23860 3016 23866
rect 2964 23802 3016 23808
rect 3068 23730 3096 26522
rect 3160 26450 3188 26998
rect 3148 26444 3200 26450
rect 3148 26386 3200 26392
rect 3148 25968 3200 25974
rect 3148 25910 3200 25916
rect 3160 25226 3188 25910
rect 3148 25220 3200 25226
rect 3148 25162 3200 25168
rect 3160 24206 3188 25162
rect 3148 24200 3200 24206
rect 3148 24142 3200 24148
rect 3056 23724 3108 23730
rect 3056 23666 3108 23672
rect 2872 23112 2924 23118
rect 2872 23054 2924 23060
rect 2884 22642 2912 23054
rect 3068 22778 3096 23666
rect 3240 23180 3292 23186
rect 3240 23122 3292 23128
rect 3056 22772 3108 22778
rect 3108 22732 3188 22760
rect 3056 22714 3108 22720
rect 2872 22636 2924 22642
rect 2872 22578 2924 22584
rect 2872 22500 2924 22506
rect 2872 22442 2924 22448
rect 2700 22086 2820 22114
rect 1492 22024 1544 22030
rect 1492 21966 1544 21972
rect 1504 21486 1532 21966
rect 1492 21480 1544 21486
rect 1492 21422 1544 21428
rect 2700 21434 2728 22086
rect 1504 21026 1532 21422
rect 2700 21406 2820 21434
rect 1504 20998 1624 21026
rect 1596 20942 1624 20998
rect 1584 20936 1636 20942
rect 1584 20878 1636 20884
rect 1596 20602 1624 20878
rect 2136 20868 2188 20874
rect 2136 20810 2188 20816
rect 1584 20596 1636 20602
rect 1584 20538 1636 20544
rect 1596 19310 1624 20538
rect 2148 20330 2176 20810
rect 2792 20398 2820 21406
rect 2884 21010 2912 22442
rect 3056 22024 3108 22030
rect 3056 21966 3108 21972
rect 3068 21622 3096 21966
rect 3056 21616 3108 21622
rect 3056 21558 3108 21564
rect 2872 21004 2924 21010
rect 2872 20946 2924 20952
rect 3160 20618 3188 22732
rect 3252 22234 3280 23122
rect 3332 22568 3384 22574
rect 3332 22510 3384 22516
rect 3240 22228 3292 22234
rect 3240 22170 3292 22176
rect 3344 21690 3372 22510
rect 3332 21684 3384 21690
rect 3332 21626 3384 21632
rect 3332 21004 3384 21010
rect 3332 20946 3384 20952
rect 3160 20590 3280 20618
rect 3056 20460 3108 20466
rect 3056 20402 3108 20408
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 2136 20324 2188 20330
rect 2136 20266 2188 20272
rect 3068 20058 3096 20402
rect 3148 20392 3200 20398
rect 3148 20334 3200 20340
rect 3056 20052 3108 20058
rect 3056 19994 3108 20000
rect 3056 19372 3108 19378
rect 3056 19314 3108 19320
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1596 18834 1624 19246
rect 3068 18834 3096 19314
rect 1584 18828 1636 18834
rect 1584 18770 1636 18776
rect 3056 18828 3108 18834
rect 3056 18770 3108 18776
rect 1860 18692 1912 18698
rect 1860 18634 1912 18640
rect 1872 18426 1900 18634
rect 1860 18420 1912 18426
rect 1860 18362 1912 18368
rect 2504 18352 2556 18358
rect 2504 18294 2556 18300
rect 2516 17202 2544 18294
rect 3160 17610 3188 20334
rect 3252 19334 3280 20590
rect 3344 20398 3372 20946
rect 3436 20913 3464 38791
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 5448 38344 5500 38350
rect 5448 38286 5500 38292
rect 5724 38344 5776 38350
rect 5724 38286 5776 38292
rect 4436 38208 4488 38214
rect 4436 38150 4488 38156
rect 4448 37942 4476 38150
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 4436 37936 4488 37942
rect 4436 37878 4488 37884
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 5460 37262 5488 38286
rect 5540 37664 5592 37670
rect 5540 37606 5592 37612
rect 5448 37256 5500 37262
rect 5448 37198 5500 37204
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 5460 36786 5488 37198
rect 5448 36780 5500 36786
rect 5448 36722 5500 36728
rect 3976 36644 4028 36650
rect 3976 36586 4028 36592
rect 3988 36174 4016 36586
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 5460 36378 5488 36722
rect 5448 36372 5500 36378
rect 5448 36314 5500 36320
rect 3976 36168 4028 36174
rect 3976 36110 4028 36116
rect 4620 36168 4672 36174
rect 4620 36110 4672 36116
rect 4252 36032 4304 36038
rect 4252 35974 4304 35980
rect 4264 35766 4292 35974
rect 3792 35760 3844 35766
rect 3792 35702 3844 35708
rect 4252 35760 4304 35766
rect 4252 35702 4304 35708
rect 3608 33312 3660 33318
rect 3608 33254 3660 33260
rect 3620 32502 3648 33254
rect 3804 33114 3832 35702
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4068 34536 4120 34542
rect 4068 34478 4120 34484
rect 4080 34202 4108 34478
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4068 34196 4120 34202
rect 4068 34138 4120 34144
rect 4632 33998 4660 36110
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 5448 35760 5500 35766
rect 5448 35702 5500 35708
rect 5460 35290 5488 35702
rect 5552 35698 5580 37606
rect 5632 37256 5684 37262
rect 5632 37198 5684 37204
rect 5644 36582 5672 37198
rect 5632 36576 5684 36582
rect 5632 36518 5684 36524
rect 5644 35834 5672 36518
rect 5736 36174 5764 38286
rect 5908 37868 5960 37874
rect 5908 37810 5960 37816
rect 5816 37120 5868 37126
rect 5816 37062 5868 37068
rect 5828 36786 5856 37062
rect 5816 36780 5868 36786
rect 5816 36722 5868 36728
rect 5724 36168 5776 36174
rect 5724 36110 5776 36116
rect 5816 36100 5868 36106
rect 5816 36042 5868 36048
rect 5632 35828 5684 35834
rect 5632 35770 5684 35776
rect 5540 35692 5592 35698
rect 5540 35634 5592 35640
rect 5448 35284 5500 35290
rect 5448 35226 5500 35232
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 4160 33992 4212 33998
rect 4160 33934 4212 33940
rect 4620 33992 4672 33998
rect 4620 33934 4672 33940
rect 4172 33658 4200 33934
rect 4160 33652 4212 33658
rect 4160 33594 4212 33600
rect 4172 33454 4200 33594
rect 4160 33448 4212 33454
rect 4160 33390 4212 33396
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 3792 33108 3844 33114
rect 3792 33050 3844 33056
rect 3608 32496 3660 32502
rect 3608 32438 3660 32444
rect 3804 31822 3832 33050
rect 3884 32904 3936 32910
rect 3884 32846 3936 32852
rect 3896 32366 3924 32846
rect 3884 32360 3936 32366
rect 3884 32302 3936 32308
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 3792 31816 3844 31822
rect 3792 31758 3844 31764
rect 4632 31754 4660 33934
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 5172 33312 5224 33318
rect 5172 33254 5224 33260
rect 5184 32978 5212 33254
rect 5172 32972 5224 32978
rect 5172 32914 5224 32920
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 5460 31754 5488 35226
rect 5552 35154 5580 35634
rect 5828 35630 5856 36042
rect 5816 35624 5868 35630
rect 5816 35566 5868 35572
rect 5816 35488 5868 35494
rect 5816 35430 5868 35436
rect 5540 35148 5592 35154
rect 5540 35090 5592 35096
rect 5552 34610 5580 35090
rect 5540 34604 5592 34610
rect 5540 34546 5592 34552
rect 5632 33992 5684 33998
rect 5632 33934 5684 33940
rect 5540 33652 5592 33658
rect 5540 33594 5592 33600
rect 5552 32842 5580 33594
rect 5644 33522 5672 33934
rect 5632 33516 5684 33522
rect 5632 33458 5684 33464
rect 5644 33114 5672 33458
rect 5828 33454 5856 35430
rect 5920 34950 5948 37810
rect 6644 37800 6696 37806
rect 6644 37742 6696 37748
rect 6656 37466 6684 37742
rect 6840 37670 6868 38830
rect 7024 38282 7052 41386
rect 17040 40656 17092 40662
rect 17040 40598 17092 40604
rect 15016 40588 15068 40594
rect 15016 40530 15068 40536
rect 13452 40112 13504 40118
rect 13452 40054 13504 40060
rect 12256 39976 12308 39982
rect 12256 39918 12308 39924
rect 12164 39840 12216 39846
rect 12164 39782 12216 39788
rect 11980 39636 12032 39642
rect 11980 39578 12032 39584
rect 8484 39500 8536 39506
rect 8484 39442 8536 39448
rect 8392 39432 8444 39438
rect 8392 39374 8444 39380
rect 8300 39296 8352 39302
rect 8300 39238 8352 39244
rect 8312 38350 8340 39238
rect 8404 38554 8432 39374
rect 8392 38548 8444 38554
rect 8392 38490 8444 38496
rect 8024 38344 8076 38350
rect 8022 38312 8024 38321
rect 8116 38344 8168 38350
rect 8076 38312 8078 38321
rect 7012 38276 7064 38282
rect 8116 38286 8168 38292
rect 8300 38344 8352 38350
rect 8300 38286 8352 38292
rect 8392 38344 8444 38350
rect 8392 38286 8444 38292
rect 8022 38247 8078 38256
rect 7012 38218 7064 38224
rect 7024 38010 7052 38218
rect 7012 38004 7064 38010
rect 7012 37946 7064 37952
rect 6828 37664 6880 37670
rect 6828 37606 6880 37612
rect 7932 37664 7984 37670
rect 7932 37606 7984 37612
rect 6644 37460 6696 37466
rect 6644 37402 6696 37408
rect 7012 37392 7064 37398
rect 7012 37334 7064 37340
rect 6000 37256 6052 37262
rect 6000 37198 6052 37204
rect 6012 36922 6040 37198
rect 6000 36916 6052 36922
rect 6000 36858 6052 36864
rect 6368 36780 6420 36786
rect 6368 36722 6420 36728
rect 6092 36712 6144 36718
rect 6092 36654 6144 36660
rect 6000 35828 6052 35834
rect 6000 35770 6052 35776
rect 6012 35154 6040 35770
rect 6000 35148 6052 35154
rect 6000 35090 6052 35096
rect 5908 34944 5960 34950
rect 5908 34886 5960 34892
rect 5920 34678 5948 34886
rect 5908 34672 5960 34678
rect 5908 34614 5960 34620
rect 6104 34610 6132 36654
rect 6380 36174 6408 36722
rect 6368 36168 6420 36174
rect 6368 36110 6420 36116
rect 6276 36100 6328 36106
rect 6276 36042 6328 36048
rect 6184 35692 6236 35698
rect 6184 35634 6236 35640
rect 6196 34678 6224 35634
rect 6288 35329 6316 36042
rect 6274 35320 6330 35329
rect 6274 35255 6330 35264
rect 6184 34672 6236 34678
rect 6184 34614 6236 34620
rect 6092 34604 6144 34610
rect 6092 34546 6144 34552
rect 6104 34474 6132 34546
rect 6092 34468 6144 34474
rect 6092 34410 6144 34416
rect 6380 33522 6408 36110
rect 7024 35698 7052 37334
rect 7944 37312 7972 37606
rect 8128 37466 8156 38286
rect 8404 38196 8432 38286
rect 8220 38168 8432 38196
rect 8116 37460 8168 37466
rect 8116 37402 8168 37408
rect 8220 37398 8248 38168
rect 8208 37392 8260 37398
rect 8208 37334 8260 37340
rect 8496 37330 8524 39442
rect 9404 39432 9456 39438
rect 9404 39374 9456 39380
rect 11244 39432 11296 39438
rect 11244 39374 11296 39380
rect 11520 39432 11572 39438
rect 11520 39374 11572 39380
rect 8576 38888 8628 38894
rect 8576 38830 8628 38836
rect 9312 38888 9364 38894
rect 9416 38876 9444 39374
rect 11060 39296 11112 39302
rect 11060 39238 11112 39244
rect 10876 39092 10928 39098
rect 10876 39034 10928 39040
rect 10232 38956 10284 38962
rect 10232 38898 10284 38904
rect 9364 38848 9444 38876
rect 9312 38830 9364 38836
rect 8588 38554 8616 38830
rect 9416 38554 9444 38848
rect 9588 38820 9640 38826
rect 9588 38762 9640 38768
rect 8576 38548 8628 38554
rect 8576 38490 8628 38496
rect 9404 38548 9456 38554
rect 9404 38490 9456 38496
rect 8852 38480 8904 38486
rect 8588 38428 8852 38434
rect 8588 38422 8904 38428
rect 8588 38418 8892 38422
rect 8576 38412 8892 38418
rect 8628 38406 8892 38412
rect 9312 38412 9364 38418
rect 8576 38354 8628 38360
rect 9312 38354 9364 38360
rect 8668 38344 8720 38350
rect 9036 38344 9088 38350
rect 8668 38286 8720 38292
rect 8850 38312 8906 38321
rect 8680 38010 8708 38286
rect 8850 38247 8906 38256
rect 9034 38312 9036 38321
rect 9088 38312 9090 38321
rect 9034 38247 9090 38256
rect 8668 38004 8720 38010
rect 8668 37946 8720 37952
rect 8864 37466 8892 38247
rect 9324 37890 9352 38354
rect 9600 38350 9628 38762
rect 9956 38752 10008 38758
rect 9956 38694 10008 38700
rect 10140 38752 10192 38758
rect 10140 38694 10192 38700
rect 9588 38344 9640 38350
rect 9588 38286 9640 38292
rect 8956 37874 9352 37890
rect 8944 37868 9364 37874
rect 8996 37862 9312 37868
rect 8944 37810 8996 37816
rect 8852 37460 8904 37466
rect 8852 37402 8904 37408
rect 8024 37324 8076 37330
rect 7944 37284 8024 37312
rect 7840 37256 7892 37262
rect 7840 37198 7892 37204
rect 7852 36378 7880 37198
rect 7472 36372 7524 36378
rect 7472 36314 7524 36320
rect 7840 36372 7892 36378
rect 7840 36314 7892 36320
rect 7288 36168 7340 36174
rect 7286 36136 7288 36145
rect 7340 36136 7342 36145
rect 7286 36071 7342 36080
rect 7012 35692 7064 35698
rect 7012 35634 7064 35640
rect 6736 35624 6788 35630
rect 6736 35566 6788 35572
rect 6552 35556 6604 35562
rect 6552 35498 6604 35504
rect 6458 35184 6514 35193
rect 6564 35154 6592 35498
rect 6748 35290 6776 35566
rect 7196 35488 7248 35494
rect 7196 35430 7248 35436
rect 6736 35284 6788 35290
rect 6736 35226 6788 35232
rect 6458 35119 6460 35128
rect 6512 35119 6514 35128
rect 6552 35148 6604 35154
rect 6460 35090 6512 35096
rect 6552 35090 6604 35096
rect 6644 35080 6696 35086
rect 6748 35068 6776 35226
rect 7208 35086 7236 35430
rect 6696 35040 6776 35068
rect 6644 35022 6696 35028
rect 6552 34944 6604 34950
rect 6552 34886 6604 34892
rect 6564 34610 6592 34886
rect 6552 34604 6604 34610
rect 6552 34546 6604 34552
rect 6644 34604 6696 34610
rect 6644 34546 6696 34552
rect 6552 34196 6604 34202
rect 6552 34138 6604 34144
rect 6000 33516 6052 33522
rect 6000 33458 6052 33464
rect 6368 33516 6420 33522
rect 6368 33458 6420 33464
rect 5816 33448 5868 33454
rect 5816 33390 5868 33396
rect 5632 33108 5684 33114
rect 5632 33050 5684 33056
rect 5540 32836 5592 32842
rect 5540 32778 5592 32784
rect 5552 32570 5580 32778
rect 5540 32564 5592 32570
rect 5644 32552 5672 33050
rect 5816 32768 5868 32774
rect 5816 32710 5868 32716
rect 5644 32524 5764 32552
rect 5540 32506 5592 32512
rect 5632 32428 5684 32434
rect 5632 32370 5684 32376
rect 5540 32360 5592 32366
rect 5540 32302 5592 32308
rect 5552 31958 5580 32302
rect 5540 31952 5592 31958
rect 5540 31894 5592 31900
rect 4632 31726 4844 31754
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4816 30841 4844 31726
rect 5264 31748 5316 31754
rect 5264 31690 5316 31696
rect 5368 31726 5488 31754
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 5276 31482 5304 31690
rect 5264 31476 5316 31482
rect 5264 31418 5316 31424
rect 4988 31272 5040 31278
rect 4988 31214 5040 31220
rect 4896 31136 4948 31142
rect 4896 31078 4948 31084
rect 4802 30832 4858 30841
rect 4802 30767 4804 30776
rect 4856 30767 4858 30776
rect 4804 30738 4856 30744
rect 3792 30728 3844 30734
rect 3792 30670 3844 30676
rect 3804 29646 3832 30670
rect 4816 30326 4844 30738
rect 4908 30734 4936 31078
rect 5000 30938 5028 31214
rect 4988 30932 5040 30938
rect 4988 30874 5040 30880
rect 4896 30728 4948 30734
rect 4896 30670 4948 30676
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 4804 30320 4856 30326
rect 4804 30262 4856 30268
rect 4896 30320 4948 30326
rect 4896 30262 4948 30268
rect 4908 30190 4936 30262
rect 4620 30184 4672 30190
rect 4620 30126 4672 30132
rect 4804 30184 4856 30190
rect 4804 30126 4856 30132
rect 4896 30184 4948 30190
rect 4896 30126 4948 30132
rect 5264 30184 5316 30190
rect 5264 30126 5316 30132
rect 4068 30048 4120 30054
rect 4068 29990 4120 29996
rect 4080 29714 4108 29990
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4632 29850 4660 30126
rect 4620 29844 4672 29850
rect 4620 29786 4672 29792
rect 4068 29708 4120 29714
rect 4068 29650 4120 29656
rect 3792 29640 3844 29646
rect 3792 29582 3844 29588
rect 3804 29306 3832 29582
rect 3792 29300 3844 29306
rect 3792 29242 3844 29248
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4632 28490 4660 29786
rect 4816 29714 4844 30126
rect 4804 29708 4856 29714
rect 4804 29650 4856 29656
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4804 29096 4856 29102
rect 4804 29038 4856 29044
rect 3884 28484 3936 28490
rect 3884 28426 3936 28432
rect 4620 28484 4672 28490
rect 4620 28426 4672 28432
rect 3792 27872 3844 27878
rect 3792 27814 3844 27820
rect 3804 27538 3832 27814
rect 3792 27532 3844 27538
rect 3792 27474 3844 27480
rect 3700 25900 3752 25906
rect 3804 25888 3832 27474
rect 3752 25860 3832 25888
rect 3700 25842 3752 25848
rect 3712 25362 3740 25842
rect 3896 25378 3924 28426
rect 4068 28416 4120 28422
rect 4068 28358 4120 28364
rect 4080 28150 4108 28358
rect 4068 28144 4120 28150
rect 4068 28086 4120 28092
rect 4080 27554 4108 28086
rect 4712 28076 4764 28082
rect 4712 28018 4764 28024
rect 4620 27940 4672 27946
rect 4620 27882 4672 27888
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3988 27526 4108 27554
rect 3988 25974 4016 27526
rect 4068 27396 4120 27402
rect 4068 27338 4120 27344
rect 4080 27130 4108 27338
rect 4344 27328 4396 27334
rect 4344 27270 4396 27276
rect 4356 27130 4384 27270
rect 4068 27124 4120 27130
rect 4068 27066 4120 27072
rect 4344 27124 4396 27130
rect 4344 27066 4396 27072
rect 4632 26926 4660 27882
rect 4620 26920 4672 26926
rect 4620 26862 4672 26868
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4344 26376 4396 26382
rect 4344 26318 4396 26324
rect 4356 26042 4384 26318
rect 4344 26036 4396 26042
rect 4344 25978 4396 25984
rect 3976 25968 4028 25974
rect 3976 25910 4028 25916
rect 4436 25968 4488 25974
rect 4436 25910 4488 25916
rect 3976 25832 4028 25838
rect 3976 25774 4028 25780
rect 4448 25786 4476 25910
rect 3988 25498 4016 25774
rect 4448 25758 4660 25786
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 3976 25492 4028 25498
rect 3976 25434 4028 25440
rect 3700 25356 3752 25362
rect 3896 25350 4016 25378
rect 3700 25298 3752 25304
rect 3792 25152 3844 25158
rect 3792 25094 3844 25100
rect 3804 24954 3832 25094
rect 3792 24948 3844 24954
rect 3792 24890 3844 24896
rect 3516 24880 3568 24886
rect 3516 24822 3568 24828
rect 3528 21593 3556 24822
rect 3884 24744 3936 24750
rect 3884 24686 3936 24692
rect 3700 24676 3752 24682
rect 3700 24618 3752 24624
rect 3712 24274 3740 24618
rect 3896 24410 3924 24686
rect 3884 24404 3936 24410
rect 3884 24346 3936 24352
rect 3700 24268 3752 24274
rect 3700 24210 3752 24216
rect 3712 23798 3740 24210
rect 3700 23792 3752 23798
rect 3700 23734 3752 23740
rect 3896 23730 3924 24346
rect 3884 23724 3936 23730
rect 3884 23666 3936 23672
rect 3988 23118 4016 25350
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4632 24138 4660 25758
rect 4724 24886 4752 28018
rect 4816 25401 4844 29038
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 5276 26586 5304 30126
rect 5368 26586 5396 31726
rect 5644 31464 5672 32370
rect 5736 32026 5764 32524
rect 5828 32366 5856 32710
rect 5816 32360 5868 32366
rect 5816 32302 5868 32308
rect 5908 32292 5960 32298
rect 5908 32234 5960 32240
rect 5724 32020 5776 32026
rect 5724 31962 5776 31968
rect 5816 31884 5868 31890
rect 5816 31826 5868 31832
rect 5724 31476 5776 31482
rect 5644 31436 5724 31464
rect 5724 31418 5776 31424
rect 5828 31414 5856 31826
rect 5920 31822 5948 32234
rect 6012 32230 6040 33458
rect 6092 33380 6144 33386
rect 6092 33322 6144 33328
rect 6000 32224 6052 32230
rect 6000 32166 6052 32172
rect 6104 31890 6132 33322
rect 6276 32836 6328 32842
rect 6276 32778 6328 32784
rect 6184 32428 6236 32434
rect 6184 32370 6236 32376
rect 6092 31884 6144 31890
rect 6092 31826 6144 31832
rect 5908 31816 5960 31822
rect 5908 31758 5960 31764
rect 5816 31408 5868 31414
rect 5816 31350 5868 31356
rect 5448 31340 5500 31346
rect 5448 31282 5500 31288
rect 5264 26580 5316 26586
rect 5264 26522 5316 26528
rect 5356 26580 5408 26586
rect 5356 26522 5408 26528
rect 5264 26444 5316 26450
rect 5264 26386 5316 26392
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4802 25392 4858 25401
rect 5276 25362 5304 26386
rect 5356 26036 5408 26042
rect 5356 25978 5408 25984
rect 5368 25362 5396 25978
rect 4802 25327 4804 25336
rect 4856 25327 4858 25336
rect 5264 25356 5316 25362
rect 4804 25298 4856 25304
rect 5264 25298 5316 25304
rect 5356 25356 5408 25362
rect 5356 25298 5408 25304
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 5276 24954 5304 25298
rect 5264 24948 5316 24954
rect 5264 24890 5316 24896
rect 4712 24880 4764 24886
rect 4712 24822 4764 24828
rect 5276 24818 5304 24890
rect 5368 24818 5396 25298
rect 5264 24812 5316 24818
rect 5264 24754 5316 24760
rect 5356 24812 5408 24818
rect 5356 24754 5408 24760
rect 4068 24132 4120 24138
rect 4068 24074 4120 24080
rect 4620 24132 4672 24138
rect 4620 24074 4672 24080
rect 4080 23594 4108 24074
rect 4632 23882 4660 24074
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4632 23854 4752 23882
rect 4620 23792 4672 23798
rect 4620 23734 4672 23740
rect 4068 23588 4120 23594
rect 4068 23530 4120 23536
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 3976 23112 4028 23118
rect 3976 23054 4028 23060
rect 3792 22568 3844 22574
rect 3792 22510 3844 22516
rect 3804 22030 3832 22510
rect 3884 22432 3936 22438
rect 3884 22374 3936 22380
rect 3792 22024 3844 22030
rect 3792 21966 3844 21972
rect 3514 21584 3570 21593
rect 3896 21554 3924 22374
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 22030 4660 23734
rect 4724 23322 4752 23854
rect 5078 23760 5134 23769
rect 5078 23695 5134 23704
rect 5092 23662 5120 23695
rect 5276 23662 5304 24754
rect 5460 23798 5488 31282
rect 5920 31278 5948 31758
rect 5540 31272 5592 31278
rect 5540 31214 5592 31220
rect 5908 31272 5960 31278
rect 5908 31214 5960 31220
rect 5552 29306 5580 31214
rect 6092 30728 6144 30734
rect 6092 30670 6144 30676
rect 5908 30116 5960 30122
rect 5908 30058 5960 30064
rect 5724 29504 5776 29510
rect 5724 29446 5776 29452
rect 5540 29300 5592 29306
rect 5540 29242 5592 29248
rect 5552 28626 5580 29242
rect 5736 28966 5764 29446
rect 5724 28960 5776 28966
rect 5724 28902 5776 28908
rect 5540 28620 5592 28626
rect 5540 28562 5592 28568
rect 5816 28484 5868 28490
rect 5816 28426 5868 28432
rect 5828 28218 5856 28426
rect 5816 28212 5868 28218
rect 5816 28154 5868 28160
rect 5540 27600 5592 27606
rect 5540 27542 5592 27548
rect 5552 27130 5580 27542
rect 5920 27130 5948 30058
rect 6000 29640 6052 29646
rect 6000 29582 6052 29588
rect 6012 29034 6040 29582
rect 6000 29028 6052 29034
rect 6000 28970 6052 28976
rect 6000 28144 6052 28150
rect 5998 28112 6000 28121
rect 6052 28112 6054 28121
rect 5998 28047 6054 28056
rect 5540 27124 5592 27130
rect 5540 27066 5592 27072
rect 5908 27124 5960 27130
rect 5908 27066 5960 27072
rect 5552 26840 5580 27066
rect 6104 27062 6132 30670
rect 6196 30598 6224 32370
rect 6288 32230 6316 32778
rect 6380 32298 6408 33458
rect 6564 32978 6592 34138
rect 6656 33590 6684 34546
rect 6748 34066 6776 35040
rect 7104 35080 7156 35086
rect 7104 35022 7156 35028
rect 7196 35080 7248 35086
rect 7196 35022 7248 35028
rect 7116 34746 7144 35022
rect 7104 34740 7156 34746
rect 7104 34682 7156 34688
rect 6828 34536 6880 34542
rect 6880 34496 6960 34524
rect 6828 34478 6880 34484
rect 6736 34060 6788 34066
rect 6736 34002 6788 34008
rect 6644 33584 6696 33590
rect 6644 33526 6696 33532
rect 6552 32972 6604 32978
rect 6552 32914 6604 32920
rect 6552 32768 6604 32774
rect 6552 32710 6604 32716
rect 6564 32502 6592 32710
rect 6552 32496 6604 32502
rect 6552 32438 6604 32444
rect 6644 32496 6696 32502
rect 6748 32484 6776 34002
rect 6828 33448 6880 33454
rect 6828 33390 6880 33396
rect 6840 32570 6868 33390
rect 6932 32978 6960 34496
rect 7104 34468 7156 34474
rect 7104 34410 7156 34416
rect 7116 33454 7144 34410
rect 7300 34202 7328 36071
rect 7380 35556 7432 35562
rect 7380 35498 7432 35504
rect 7392 35193 7420 35498
rect 7378 35184 7434 35193
rect 7378 35119 7434 35128
rect 7392 35086 7420 35119
rect 7484 35086 7512 36314
rect 7564 36100 7616 36106
rect 7564 36042 7616 36048
rect 7748 36100 7800 36106
rect 7748 36042 7800 36048
rect 7576 35834 7604 36042
rect 7564 35828 7616 35834
rect 7564 35770 7616 35776
rect 7760 35698 7788 36042
rect 7564 35692 7616 35698
rect 7564 35634 7616 35640
rect 7748 35692 7800 35698
rect 7748 35634 7800 35640
rect 7576 35329 7604 35634
rect 7562 35320 7618 35329
rect 7760 35290 7788 35634
rect 7562 35255 7618 35264
rect 7748 35284 7800 35290
rect 7748 35226 7800 35232
rect 7380 35080 7432 35086
rect 7380 35022 7432 35028
rect 7472 35080 7524 35086
rect 7472 35022 7524 35028
rect 7288 34196 7340 34202
rect 7288 34138 7340 34144
rect 7196 33516 7248 33522
rect 7196 33458 7248 33464
rect 7288 33516 7340 33522
rect 7288 33458 7340 33464
rect 7104 33448 7156 33454
rect 7104 33390 7156 33396
rect 7012 33380 7064 33386
rect 7012 33322 7064 33328
rect 6920 32972 6972 32978
rect 6920 32914 6972 32920
rect 6828 32564 6880 32570
rect 6828 32506 6880 32512
rect 6932 32502 6960 32914
rect 6696 32456 6776 32484
rect 6920 32496 6972 32502
rect 6644 32438 6696 32444
rect 6920 32438 6972 32444
rect 6368 32292 6420 32298
rect 6368 32234 6420 32240
rect 6276 32224 6328 32230
rect 6276 32166 6328 32172
rect 6552 32224 6604 32230
rect 6552 32166 6604 32172
rect 6276 32020 6328 32026
rect 6276 31962 6328 31968
rect 6184 30592 6236 30598
rect 6184 30534 6236 30540
rect 6196 30122 6224 30534
rect 6184 30116 6236 30122
rect 6184 30058 6236 30064
rect 6184 29504 6236 29510
rect 6184 29446 6236 29452
rect 6196 29170 6224 29446
rect 6184 29164 6236 29170
rect 6184 29106 6236 29112
rect 6184 29028 6236 29034
rect 6184 28970 6236 28976
rect 6196 28762 6224 28970
rect 6184 28756 6236 28762
rect 6184 28698 6236 28704
rect 6092 27056 6144 27062
rect 6092 26998 6144 27004
rect 5816 26988 5868 26994
rect 5816 26930 5868 26936
rect 5908 26988 5960 26994
rect 5908 26930 5960 26936
rect 5552 26812 5764 26840
rect 5632 26308 5684 26314
rect 5632 26250 5684 26256
rect 5644 26042 5672 26250
rect 5632 26036 5684 26042
rect 5632 25978 5684 25984
rect 5540 25696 5592 25702
rect 5540 25638 5592 25644
rect 5552 25294 5580 25638
rect 5644 25294 5672 25978
rect 5540 25288 5592 25294
rect 5540 25230 5592 25236
rect 5632 25288 5684 25294
rect 5632 25230 5684 25236
rect 5540 25152 5592 25158
rect 5540 25094 5592 25100
rect 5552 24818 5580 25094
rect 5736 24818 5764 26812
rect 5828 26246 5856 26930
rect 5816 26240 5868 26246
rect 5816 26182 5868 26188
rect 5816 25220 5868 25226
rect 5920 25208 5948 26930
rect 6000 26784 6052 26790
rect 6000 26726 6052 26732
rect 6012 26382 6040 26726
rect 6000 26376 6052 26382
rect 6000 26318 6052 26324
rect 6092 26376 6144 26382
rect 6092 26318 6144 26324
rect 5868 25180 5948 25208
rect 5816 25162 5868 25168
rect 5540 24812 5592 24818
rect 5540 24754 5592 24760
rect 5724 24812 5776 24818
rect 5724 24754 5776 24760
rect 5448 23792 5500 23798
rect 5448 23734 5500 23740
rect 5552 23662 5580 24754
rect 5724 24268 5776 24274
rect 5724 24210 5776 24216
rect 5632 24064 5684 24070
rect 5632 24006 5684 24012
rect 5644 23866 5672 24006
rect 5632 23860 5684 23866
rect 5632 23802 5684 23808
rect 5080 23656 5132 23662
rect 4816 23616 5080 23644
rect 4712 23316 4764 23322
rect 4712 23258 4764 23264
rect 4724 22710 4752 23258
rect 4712 22704 4764 22710
rect 4712 22646 4764 22652
rect 4712 22500 4764 22506
rect 4712 22442 4764 22448
rect 4620 22024 4672 22030
rect 4618 21992 4620 22001
rect 4672 21992 4674 22001
rect 4618 21927 4674 21936
rect 4724 21690 4752 22442
rect 4712 21684 4764 21690
rect 4712 21626 4764 21632
rect 4816 21570 4844 23616
rect 5080 23598 5132 23604
rect 5264 23656 5316 23662
rect 5264 23598 5316 23604
rect 5540 23656 5592 23662
rect 5540 23598 5592 23604
rect 5632 23520 5684 23526
rect 5446 23488 5502 23497
rect 5632 23462 5684 23468
rect 5446 23423 5502 23432
rect 5264 23112 5316 23118
rect 5264 23054 5316 23060
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 5276 22506 5304 23054
rect 5264 22500 5316 22506
rect 5264 22442 5316 22448
rect 5460 22094 5488 23423
rect 5644 23254 5672 23462
rect 5632 23248 5684 23254
rect 5632 23190 5684 23196
rect 5632 23044 5684 23050
rect 5632 22986 5684 22992
rect 5644 22438 5672 22986
rect 5736 22642 5764 24210
rect 5724 22636 5776 22642
rect 5724 22578 5776 22584
rect 5632 22432 5684 22438
rect 5632 22374 5684 22380
rect 5276 22066 5488 22094
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4448 21554 4844 21570
rect 3514 21519 3570 21528
rect 3608 21548 3660 21554
rect 3422 20904 3478 20913
rect 3422 20839 3478 20848
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 3424 19848 3476 19854
rect 3424 19790 3476 19796
rect 3436 19514 3464 19790
rect 3424 19508 3476 19514
rect 3424 19450 3476 19456
rect 3528 19446 3556 21519
rect 3608 21490 3660 21496
rect 3700 21548 3752 21554
rect 3700 21490 3752 21496
rect 3884 21548 3936 21554
rect 3884 21490 3936 21496
rect 4436 21548 4844 21554
rect 4488 21542 4844 21548
rect 5170 21584 5226 21593
rect 4436 21490 4488 21496
rect 3620 21457 3648 21490
rect 3606 21448 3662 21457
rect 3606 21383 3662 21392
rect 3608 20800 3660 20806
rect 3712 20788 3740 21490
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 3792 20868 3844 20874
rect 3792 20810 3844 20816
rect 3660 20760 3740 20788
rect 3608 20742 3660 20748
rect 3620 19922 3648 20742
rect 3804 20534 3832 20810
rect 4436 20800 4488 20806
rect 4436 20742 4488 20748
rect 3792 20528 3844 20534
rect 3792 20470 3844 20476
rect 3608 19916 3660 19922
rect 3608 19858 3660 19864
rect 3516 19440 3568 19446
rect 3516 19382 3568 19388
rect 3252 19306 3372 19334
rect 3240 18692 3292 18698
rect 3240 18634 3292 18640
rect 3148 17604 3200 17610
rect 3148 17546 3200 17552
rect 2780 17536 2832 17542
rect 2780 17478 2832 17484
rect 2792 17270 2820 17478
rect 2780 17264 2832 17270
rect 2780 17206 2832 17212
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 3252 16182 3280 18634
rect 3344 18426 3372 19306
rect 3804 18902 3832 20470
rect 4448 20398 4476 20742
rect 4436 20392 4488 20398
rect 4436 20334 4488 20340
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3884 19712 3936 19718
rect 3884 19654 3936 19660
rect 3896 19514 3924 19654
rect 3884 19508 3936 19514
rect 3884 19450 3936 19456
rect 4632 19310 4660 21542
rect 5170 21519 5226 21528
rect 5184 21486 5212 21519
rect 5172 21480 5224 21486
rect 5172 21422 5224 21428
rect 5080 21412 5132 21418
rect 5080 21354 5132 21360
rect 5092 21049 5120 21354
rect 4894 21040 4950 21049
rect 4894 20975 4950 20984
rect 5078 21040 5134 21049
rect 5078 20975 5080 20984
rect 4908 20942 4936 20975
rect 5132 20975 5134 20984
rect 5080 20946 5132 20952
rect 4896 20936 4948 20942
rect 4896 20878 4948 20884
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 5276 20466 5304 22066
rect 5632 22024 5684 22030
rect 5632 21966 5684 21972
rect 5448 21956 5500 21962
rect 5448 21898 5500 21904
rect 5356 21888 5408 21894
rect 5356 21830 5408 21836
rect 5368 21690 5396 21830
rect 5356 21684 5408 21690
rect 5356 21626 5408 21632
rect 5460 21486 5488 21898
rect 5448 21480 5500 21486
rect 5448 21422 5500 21428
rect 5644 21350 5672 21966
rect 5724 21956 5776 21962
rect 5724 21898 5776 21904
rect 5736 21554 5764 21898
rect 5828 21690 5856 25162
rect 6104 25129 6132 26318
rect 6196 25378 6224 28698
rect 6288 26858 6316 31962
rect 6564 30734 6592 32166
rect 6656 31958 6684 32438
rect 6920 32360 6972 32366
rect 7024 32348 7052 33322
rect 7208 32434 7236 33458
rect 7300 32842 7328 33458
rect 7392 33386 7420 35022
rect 7840 33516 7892 33522
rect 7840 33458 7892 33464
rect 7472 33448 7524 33454
rect 7472 33390 7524 33396
rect 7380 33380 7432 33386
rect 7380 33322 7432 33328
rect 7288 32836 7340 32842
rect 7288 32778 7340 32784
rect 7196 32428 7248 32434
rect 7196 32370 7248 32376
rect 6972 32320 7052 32348
rect 6920 32302 6972 32308
rect 6644 31952 6696 31958
rect 6644 31894 6696 31900
rect 6552 30728 6604 30734
rect 6552 30670 6604 30676
rect 6552 29708 6604 29714
rect 6552 29650 6604 29656
rect 6460 28416 6512 28422
rect 6380 28376 6460 28404
rect 6380 28082 6408 28376
rect 6460 28358 6512 28364
rect 6460 28212 6512 28218
rect 6460 28154 6512 28160
rect 6368 28076 6420 28082
rect 6368 28018 6420 28024
rect 6472 27606 6500 28154
rect 6564 28150 6592 29650
rect 6552 28144 6604 28150
rect 6552 28086 6604 28092
rect 6460 27600 6512 27606
rect 6460 27542 6512 27548
rect 6368 26988 6420 26994
rect 6368 26930 6420 26936
rect 6276 26852 6328 26858
rect 6276 26794 6328 26800
rect 6380 26450 6408 26930
rect 6460 26784 6512 26790
rect 6460 26726 6512 26732
rect 6472 26586 6500 26726
rect 6460 26580 6512 26586
rect 6460 26522 6512 26528
rect 6656 26450 6684 31894
rect 7300 31482 7328 32778
rect 7380 32564 7432 32570
rect 7380 32506 7432 32512
rect 7392 32026 7420 32506
rect 7484 32434 7512 33390
rect 7656 33312 7708 33318
rect 7656 33254 7708 33260
rect 7668 32978 7696 33254
rect 7656 32972 7708 32978
rect 7656 32914 7708 32920
rect 7852 32570 7880 33458
rect 7840 32564 7892 32570
rect 7840 32506 7892 32512
rect 7472 32428 7524 32434
rect 7472 32370 7524 32376
rect 7380 32020 7432 32026
rect 7380 31962 7432 31968
rect 7840 31748 7892 31754
rect 7840 31690 7892 31696
rect 7288 31476 7340 31482
rect 7288 31418 7340 31424
rect 7380 31340 7432 31346
rect 7380 31282 7432 31288
rect 7392 31142 7420 31282
rect 7852 31278 7880 31690
rect 7748 31272 7800 31278
rect 7748 31214 7800 31220
rect 7840 31272 7892 31278
rect 7840 31214 7892 31220
rect 7380 31136 7432 31142
rect 7380 31078 7432 31084
rect 7392 30258 7420 31078
rect 7760 30818 7788 31214
rect 7668 30790 7788 30818
rect 7668 30734 7696 30790
rect 7656 30728 7708 30734
rect 7656 30670 7708 30676
rect 7380 30252 7432 30258
rect 7380 30194 7432 30200
rect 6828 29844 6880 29850
rect 6828 29786 6880 29792
rect 6840 29306 6868 29786
rect 7196 29572 7248 29578
rect 7196 29514 7248 29520
rect 6828 29300 6880 29306
rect 6828 29242 6880 29248
rect 7208 29238 7236 29514
rect 7196 29232 7248 29238
rect 7196 29174 7248 29180
rect 7208 29102 7236 29174
rect 6828 29096 6880 29102
rect 6828 29038 6880 29044
rect 7104 29096 7156 29102
rect 7104 29038 7156 29044
rect 7196 29096 7248 29102
rect 7196 29038 7248 29044
rect 6840 28626 6868 29038
rect 7116 28762 7144 29038
rect 7104 28756 7156 28762
rect 7104 28698 7156 28704
rect 6828 28620 6880 28626
rect 6828 28562 6880 28568
rect 6840 27538 6868 28562
rect 7288 28416 7340 28422
rect 7288 28358 7340 28364
rect 7104 28144 7156 28150
rect 7102 28112 7104 28121
rect 7156 28112 7158 28121
rect 7102 28047 7158 28056
rect 7300 27878 7328 28358
rect 6920 27872 6972 27878
rect 6920 27814 6972 27820
rect 7288 27872 7340 27878
rect 7288 27814 7340 27820
rect 6828 27532 6880 27538
rect 6828 27474 6880 27480
rect 6736 27124 6788 27130
rect 6736 27066 6788 27072
rect 6748 26761 6776 27066
rect 6828 26988 6880 26994
rect 6828 26930 6880 26936
rect 6734 26752 6790 26761
rect 6734 26687 6790 26696
rect 6368 26444 6420 26450
rect 6644 26444 6696 26450
rect 6420 26404 6500 26432
rect 6368 26386 6420 26392
rect 6276 26308 6328 26314
rect 6276 26250 6328 26256
rect 6288 25974 6316 26250
rect 6276 25968 6328 25974
rect 6276 25910 6328 25916
rect 6368 25900 6420 25906
rect 6368 25842 6420 25848
rect 6380 25498 6408 25842
rect 6368 25492 6420 25498
rect 6368 25434 6420 25440
rect 6196 25350 6316 25378
rect 6288 25294 6316 25350
rect 6472 25294 6500 26404
rect 6644 26386 6696 26392
rect 6656 26058 6684 26386
rect 6748 26314 6776 26687
rect 6840 26586 6868 26930
rect 6828 26580 6880 26586
rect 6828 26522 6880 26528
rect 6828 26376 6880 26382
rect 6828 26318 6880 26324
rect 6736 26308 6788 26314
rect 6736 26250 6788 26256
rect 6656 26030 6776 26058
rect 6552 25900 6604 25906
rect 6604 25860 6684 25888
rect 6552 25842 6604 25848
rect 6552 25764 6604 25770
rect 6552 25706 6604 25712
rect 6184 25288 6236 25294
rect 6184 25230 6236 25236
rect 6276 25288 6328 25294
rect 6460 25288 6512 25294
rect 6276 25230 6328 25236
rect 6380 25248 6460 25276
rect 6090 25120 6146 25129
rect 6090 25055 6146 25064
rect 6092 24812 6144 24818
rect 6196 24800 6224 25230
rect 6144 24772 6224 24800
rect 6092 24754 6144 24760
rect 5908 24608 5960 24614
rect 5908 24550 5960 24556
rect 5816 21684 5868 21690
rect 5816 21626 5868 21632
rect 5920 21554 5948 24550
rect 6000 24132 6052 24138
rect 6000 24074 6052 24080
rect 6012 23866 6040 24074
rect 6104 23905 6132 24754
rect 6380 24449 6408 25248
rect 6460 25230 6512 25236
rect 6460 25152 6512 25158
rect 6460 25094 6512 25100
rect 6366 24440 6422 24449
rect 6366 24375 6422 24384
rect 6380 24342 6408 24375
rect 6368 24336 6420 24342
rect 6368 24278 6420 24284
rect 6276 24200 6328 24206
rect 6196 24148 6276 24154
rect 6196 24142 6328 24148
rect 6196 24126 6316 24142
rect 6090 23896 6146 23905
rect 6000 23860 6052 23866
rect 6090 23831 6146 23840
rect 6000 23802 6052 23808
rect 6196 23730 6224 24126
rect 6184 23724 6236 23730
rect 6184 23666 6236 23672
rect 6276 23724 6328 23730
rect 6276 23666 6328 23672
rect 6196 23633 6224 23666
rect 6182 23624 6238 23633
rect 6182 23559 6238 23568
rect 6184 23520 6236 23526
rect 6184 23462 6236 23468
rect 6092 23112 6144 23118
rect 6092 23054 6144 23060
rect 6104 21842 6132 23054
rect 6196 22642 6224 23462
rect 6288 23186 6316 23666
rect 6368 23520 6420 23526
rect 6368 23462 6420 23468
rect 6276 23180 6328 23186
rect 6276 23122 6328 23128
rect 6380 23118 6408 23462
rect 6368 23112 6420 23118
rect 6368 23054 6420 23060
rect 6276 23044 6328 23050
rect 6276 22986 6328 22992
rect 6184 22636 6236 22642
rect 6184 22578 6236 22584
rect 6012 21814 6132 21842
rect 5724 21548 5776 21554
rect 5724 21490 5776 21496
rect 5908 21548 5960 21554
rect 5908 21490 5960 21496
rect 5816 21412 5868 21418
rect 5816 21354 5868 21360
rect 5632 21344 5684 21350
rect 5632 21286 5684 21292
rect 5448 20936 5500 20942
rect 5448 20878 5500 20884
rect 5356 20868 5408 20874
rect 5356 20810 5408 20816
rect 5368 20602 5396 20810
rect 5356 20596 5408 20602
rect 5356 20538 5408 20544
rect 5460 20482 5488 20878
rect 5538 20632 5594 20641
rect 5538 20567 5594 20576
rect 5552 20534 5580 20567
rect 5644 20534 5672 21286
rect 5722 21176 5778 21185
rect 5722 21111 5778 21120
rect 5264 20460 5316 20466
rect 5264 20402 5316 20408
rect 5368 20454 5488 20482
rect 5540 20528 5592 20534
rect 5540 20470 5592 20476
rect 5632 20528 5684 20534
rect 5632 20470 5684 20476
rect 5736 20466 5764 21111
rect 5724 20460 5776 20466
rect 4804 20256 4856 20262
rect 4804 20198 4856 20204
rect 4816 19514 4844 20198
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4804 19508 4856 19514
rect 4804 19450 4856 19456
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 4068 19304 4120 19310
rect 4068 19246 4120 19252
rect 4620 19304 4672 19310
rect 4620 19246 4672 19252
rect 3792 18896 3844 18902
rect 3792 18838 3844 18844
rect 3804 18630 3832 18838
rect 4080 18834 4108 19246
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4068 18828 4120 18834
rect 4068 18770 4120 18776
rect 4436 18828 4488 18834
rect 4436 18770 4488 18776
rect 3792 18624 3844 18630
rect 3792 18566 3844 18572
rect 4068 18624 4120 18630
rect 4068 18566 4120 18572
rect 3332 18420 3384 18426
rect 3332 18362 3384 18368
rect 3700 18420 3752 18426
rect 3700 18362 3752 18368
rect 3712 18193 3740 18362
rect 3804 18204 3832 18566
rect 4080 18358 4108 18566
rect 4068 18352 4120 18358
rect 4068 18294 4120 18300
rect 4160 18352 4212 18358
rect 4160 18294 4212 18300
rect 4172 18204 4200 18294
rect 3698 18184 3754 18193
rect 3698 18119 3754 18128
rect 3804 18176 4200 18204
rect 3804 17270 3832 18176
rect 4448 18086 4476 18770
rect 4632 18222 4660 19110
rect 4724 18766 4752 19110
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4816 18426 4844 19450
rect 4896 19304 4948 19310
rect 4896 19246 4948 19252
rect 4908 18970 4936 19246
rect 4988 19236 5040 19242
rect 4988 19178 5040 19184
rect 4896 18964 4948 18970
rect 4896 18906 4948 18912
rect 5000 18766 5028 19178
rect 5080 18964 5132 18970
rect 5080 18906 5132 18912
rect 5092 18834 5120 18906
rect 5184 18834 5212 19450
rect 5080 18828 5132 18834
rect 5080 18770 5132 18776
rect 5172 18828 5224 18834
rect 5172 18770 5224 18776
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 4620 18216 4672 18222
rect 4620 18158 4672 18164
rect 4710 18184 4766 18193
rect 4710 18119 4766 18128
rect 4724 18086 4752 18119
rect 4436 18080 4488 18086
rect 4712 18080 4764 18086
rect 4488 18040 4660 18068
rect 4436 18022 4488 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17746 4660 18040
rect 4712 18022 4764 18028
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 3792 17264 3844 17270
rect 3792 17206 3844 17212
rect 3804 16522 3832 17206
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4816 16658 4844 18362
rect 5276 17746 5304 19654
rect 5368 18358 5396 20454
rect 5724 20402 5776 20408
rect 5448 20392 5500 20398
rect 5448 20334 5500 20340
rect 5460 19310 5488 20334
rect 5632 20256 5684 20262
rect 5632 20198 5684 20204
rect 5644 19854 5672 20198
rect 5828 20058 5856 21354
rect 6012 21026 6040 21814
rect 6092 21684 6144 21690
rect 6092 21626 6144 21632
rect 5920 20998 6040 21026
rect 5816 20052 5868 20058
rect 5816 19994 5868 20000
rect 5724 19984 5776 19990
rect 5724 19926 5776 19932
rect 5736 19854 5764 19926
rect 5632 19848 5684 19854
rect 5632 19790 5684 19796
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 5448 19304 5500 19310
rect 5448 19246 5500 19252
rect 5448 18692 5500 18698
rect 5448 18634 5500 18640
rect 5460 18426 5488 18634
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 5356 18352 5408 18358
rect 5356 18294 5408 18300
rect 5552 18222 5580 19314
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 5448 18148 5500 18154
rect 5448 18090 5500 18096
rect 5264 17740 5316 17746
rect 5264 17682 5316 17688
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 5276 17338 5304 17682
rect 5356 17536 5408 17542
rect 5356 17478 5408 17484
rect 5368 17338 5396 17478
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 5460 17218 5488 18090
rect 5368 17190 5488 17218
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 3792 16516 3844 16522
rect 3792 16458 3844 16464
rect 3804 16182 3832 16458
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 3240 16176 3292 16182
rect 3240 16118 3292 16124
rect 3792 16176 3844 16182
rect 3792 16118 3844 16124
rect 3252 12986 3280 16118
rect 3804 13258 3832 16118
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 5264 15564 5316 15570
rect 5264 15506 5316 15512
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 4632 15162 4660 15302
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 5276 15026 5304 15506
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4632 14550 4660 14894
rect 4620 14544 4672 14550
rect 4620 14486 4672 14492
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 4264 14074 4292 14418
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 4712 14408 4764 14414
rect 4712 14350 4764 14356
rect 4252 14068 4304 14074
rect 4252 14010 4304 14016
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 4172 13716 4200 13874
rect 4356 13802 4384 14350
rect 4724 13938 4752 14350
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4528 13932 4580 13938
rect 4712 13932 4764 13938
rect 4580 13892 4660 13920
rect 4528 13874 4580 13880
rect 4344 13796 4396 13802
rect 4344 13738 4396 13744
rect 4080 13688 4200 13716
rect 4080 13530 4108 13688
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4632 13530 4660 13892
rect 4712 13874 4764 13880
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4160 13456 4212 13462
rect 4160 13398 4212 13404
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 3792 13252 3844 13258
rect 3792 13194 3844 13200
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 3252 11694 3280 12922
rect 3804 12918 3832 13194
rect 3792 12912 3844 12918
rect 3792 12854 3844 12860
rect 3988 12238 4016 13262
rect 4172 13258 4200 13398
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4724 13308 4752 13874
rect 5172 13796 5224 13802
rect 5172 13738 5224 13744
rect 5184 13326 5212 13738
rect 4804 13320 4856 13326
rect 4724 13280 4804 13308
rect 4160 13252 4212 13258
rect 4160 13194 4212 13200
rect 4172 12730 4200 13194
rect 4632 12986 4660 13262
rect 4724 12986 4752 13280
rect 4804 13262 4856 13268
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 4620 12980 4672 12986
rect 4356 12940 4568 12968
rect 4356 12850 4384 12940
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 4436 12844 4488 12850
rect 4436 12786 4488 12792
rect 4080 12702 4200 12730
rect 4448 12714 4476 12786
rect 4540 12730 4568 12940
rect 4620 12922 4672 12928
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4632 12850 4752 12866
rect 4620 12844 4752 12850
rect 4672 12838 4752 12844
rect 4620 12786 4672 12792
rect 4436 12708 4488 12714
rect 4080 12434 4108 12702
rect 4540 12702 4660 12730
rect 4436 12650 4488 12656
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4080 12406 4200 12434
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3804 11830 3832 12038
rect 4172 11898 4200 12406
rect 4632 12374 4660 12702
rect 4724 12442 4752 12838
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4620 12368 4672 12374
rect 4816 12322 4844 13126
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4894 12880 4950 12889
rect 4894 12815 4896 12824
rect 4948 12815 4950 12824
rect 4896 12786 4948 12792
rect 5276 12714 5304 14962
rect 5368 13530 5396 17190
rect 5448 17128 5500 17134
rect 5448 17070 5500 17076
rect 5460 16266 5488 17070
rect 5460 16238 5580 16266
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5460 15706 5488 16050
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5552 15586 5580 16238
rect 5460 15558 5580 15586
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5264 12708 5316 12714
rect 5264 12650 5316 12656
rect 4620 12310 4672 12316
rect 4724 12306 4844 12322
rect 4712 12300 4844 12306
rect 4764 12294 4844 12300
rect 4712 12242 4764 12248
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 3792 11824 3844 11830
rect 3792 11766 3844 11772
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 3528 11150 3556 11630
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 1860 11008 1912 11014
rect 1858 10976 1860 10985
rect 1912 10976 1914 10985
rect 1858 10911 1914 10920
rect 3528 10130 3556 11086
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 4724 9994 4752 11834
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4712 9988 4764 9994
rect 4712 9930 4764 9936
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4724 8566 4752 9930
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5276 9042 5304 12650
rect 5460 12646 5488 15558
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5552 15162 5580 15438
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5552 12850 5580 13126
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 5460 12442 5488 12582
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5552 11898 5580 12242
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5644 8634 5672 19790
rect 5724 19440 5776 19446
rect 5724 19382 5776 19388
rect 5736 15162 5764 19382
rect 5920 19310 5948 20998
rect 6000 20936 6052 20942
rect 6104 20924 6132 21626
rect 6196 21078 6224 22578
rect 6288 22094 6316 22986
rect 6472 22166 6500 25094
rect 6564 24585 6592 25706
rect 6550 24576 6606 24585
rect 6550 24511 6606 24520
rect 6564 24206 6592 24511
rect 6552 24200 6604 24206
rect 6552 24142 6604 24148
rect 6550 23896 6606 23905
rect 6550 23831 6606 23840
rect 6564 23730 6592 23831
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 6460 22160 6512 22166
rect 6460 22102 6512 22108
rect 6288 22066 6408 22094
rect 6276 22024 6328 22030
rect 6276 21966 6328 21972
rect 6288 21146 6316 21966
rect 6276 21140 6328 21146
rect 6276 21082 6328 21088
rect 6184 21072 6236 21078
rect 6184 21014 6236 21020
rect 6184 20936 6236 20942
rect 6104 20896 6184 20924
rect 6000 20878 6052 20884
rect 6184 20878 6236 20884
rect 6012 20602 6040 20878
rect 6380 20602 6408 22066
rect 6460 22024 6512 22030
rect 6656 21978 6684 25860
rect 6748 24614 6776 26030
rect 6840 25906 6868 26318
rect 6828 25900 6880 25906
rect 6828 25842 6880 25848
rect 6932 25786 6960 27814
rect 7288 27056 7340 27062
rect 7288 26998 7340 27004
rect 7012 26512 7064 26518
rect 7012 26454 7064 26460
rect 7024 25906 7052 26454
rect 7300 26382 7328 26998
rect 7288 26376 7340 26382
rect 7288 26318 7340 26324
rect 7104 26308 7156 26314
rect 7104 26250 7156 26256
rect 7116 26042 7144 26250
rect 7104 26036 7156 26042
rect 7104 25978 7156 25984
rect 7012 25900 7064 25906
rect 7012 25842 7064 25848
rect 7196 25900 7248 25906
rect 7196 25842 7248 25848
rect 6840 25758 6960 25786
rect 6736 24608 6788 24614
rect 6736 24550 6788 24556
rect 6840 24426 6868 25758
rect 7012 25696 7064 25702
rect 7012 25638 7064 25644
rect 6920 25492 6972 25498
rect 6920 25434 6972 25440
rect 6748 24398 6868 24426
rect 6748 23866 6776 24398
rect 6828 24336 6880 24342
rect 6828 24278 6880 24284
rect 6736 23860 6788 23866
rect 6736 23802 6788 23808
rect 6840 23798 6868 24278
rect 6828 23792 6880 23798
rect 6828 23734 6880 23740
rect 6736 23112 6788 23118
rect 6736 23054 6788 23060
rect 6748 22778 6776 23054
rect 6736 22772 6788 22778
rect 6736 22714 6788 22720
rect 6736 22568 6788 22574
rect 6736 22510 6788 22516
rect 6460 21966 6512 21972
rect 6000 20596 6052 20602
rect 6000 20538 6052 20544
rect 6368 20596 6420 20602
rect 6368 20538 6420 20544
rect 6366 20496 6422 20505
rect 6366 20431 6422 20440
rect 5998 20360 6054 20369
rect 5998 20295 6054 20304
rect 5908 19304 5960 19310
rect 5908 19246 5960 19252
rect 6012 17134 6040 20295
rect 6380 19990 6408 20431
rect 6472 19990 6500 21966
rect 6564 21950 6684 21978
rect 6564 20262 6592 21950
rect 6644 21888 6696 21894
rect 6644 21830 6696 21836
rect 6656 21350 6684 21830
rect 6644 21344 6696 21350
rect 6644 21286 6696 21292
rect 6748 21185 6776 22510
rect 6828 21480 6880 21486
rect 6828 21422 6880 21428
rect 6734 21176 6790 21185
rect 6734 21111 6736 21120
rect 6788 21111 6790 21120
rect 6736 21082 6788 21088
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 6644 20324 6696 20330
rect 6644 20266 6696 20272
rect 6552 20256 6604 20262
rect 6552 20198 6604 20204
rect 6368 19984 6420 19990
rect 6182 19952 6238 19961
rect 6368 19926 6420 19932
rect 6460 19984 6512 19990
rect 6460 19926 6512 19932
rect 6182 19887 6238 19896
rect 6196 19854 6224 19887
rect 6380 19854 6408 19926
rect 6184 19848 6236 19854
rect 6184 19790 6236 19796
rect 6368 19848 6420 19854
rect 6368 19790 6420 19796
rect 6000 17128 6052 17134
rect 6000 17070 6052 17076
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 5816 16040 5868 16046
rect 5816 15982 5868 15988
rect 5828 15570 5856 15982
rect 6104 15706 6132 16594
rect 6092 15700 6144 15706
rect 6092 15642 6144 15648
rect 6000 15632 6052 15638
rect 6196 15586 6224 19790
rect 6656 19786 6684 20266
rect 6748 20058 6776 20878
rect 6736 20052 6788 20058
rect 6736 19994 6788 20000
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 6644 19780 6696 19786
rect 6644 19722 6696 19728
rect 6656 19378 6684 19722
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6748 19310 6776 19790
rect 6840 19514 6868 21422
rect 6828 19508 6880 19514
rect 6828 19450 6880 19456
rect 6736 19304 6788 19310
rect 6736 19246 6788 19252
rect 6552 17264 6604 17270
rect 6552 17206 6604 17212
rect 6564 16794 6592 17206
rect 6932 17202 6960 25434
rect 7024 25294 7052 25638
rect 7012 25288 7064 25294
rect 7012 25230 7064 25236
rect 7102 25256 7158 25265
rect 7102 25191 7104 25200
rect 7156 25191 7158 25200
rect 7104 25162 7156 25168
rect 7012 22024 7064 22030
rect 7012 21966 7064 21972
rect 7024 21078 7052 21966
rect 7104 21956 7156 21962
rect 7104 21898 7156 21904
rect 7116 21457 7144 21898
rect 7102 21448 7158 21457
rect 7102 21383 7158 21392
rect 7012 21072 7064 21078
rect 7012 21014 7064 21020
rect 7012 20868 7064 20874
rect 7012 20810 7064 20816
rect 7024 20505 7052 20810
rect 7116 20534 7144 21383
rect 7208 20942 7236 25842
rect 7300 25294 7328 26318
rect 7288 25288 7340 25294
rect 7288 25230 7340 25236
rect 7392 24614 7420 30194
rect 7668 30054 7696 30670
rect 7852 30394 7880 31214
rect 7840 30388 7892 30394
rect 7840 30330 7892 30336
rect 7840 30116 7892 30122
rect 7840 30058 7892 30064
rect 7656 30048 7708 30054
rect 7656 29990 7708 29996
rect 7564 27940 7616 27946
rect 7564 27882 7616 27888
rect 7472 25900 7524 25906
rect 7472 25842 7524 25848
rect 7484 25430 7512 25842
rect 7472 25424 7524 25430
rect 7472 25366 7524 25372
rect 7576 25242 7604 27882
rect 7484 25214 7604 25242
rect 7288 24608 7340 24614
rect 7288 24550 7340 24556
rect 7380 24608 7432 24614
rect 7380 24550 7432 24556
rect 7196 20936 7248 20942
rect 7196 20878 7248 20884
rect 7104 20528 7156 20534
rect 7010 20496 7066 20505
rect 7104 20470 7156 20476
rect 7010 20431 7066 20440
rect 7116 20058 7144 20470
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7116 19922 7144 19994
rect 7104 19916 7156 19922
rect 7104 19858 7156 19864
rect 7208 19802 7236 20878
rect 7116 19774 7236 19802
rect 7012 18828 7064 18834
rect 7012 18770 7064 18776
rect 7024 18222 7052 18770
rect 7012 18216 7064 18222
rect 7012 18158 7064 18164
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6000 15574 6052 15580
rect 5816 15564 5868 15570
rect 5816 15506 5868 15512
rect 5908 15564 5960 15570
rect 5908 15506 5960 15512
rect 5816 15428 5868 15434
rect 5816 15370 5868 15376
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5828 14618 5856 15370
rect 5920 15026 5948 15506
rect 6012 15026 6040 15574
rect 6104 15558 6224 15586
rect 5908 15020 5960 15026
rect 5908 14962 5960 14968
rect 6000 15020 6052 15026
rect 6000 14962 6052 14968
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5920 14414 5948 14962
rect 5908 14408 5960 14414
rect 5908 14350 5960 14356
rect 5920 14006 5948 14350
rect 6012 14278 6040 14962
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 6012 14074 6040 14214
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 5908 14000 5960 14006
rect 5908 13942 5960 13948
rect 5724 13796 5776 13802
rect 5724 13738 5776 13744
rect 5736 12782 5764 13738
rect 5920 13530 5948 13942
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5828 12646 5856 13262
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5920 12753 5948 12786
rect 5906 12744 5962 12753
rect 5906 12679 5962 12688
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5908 12368 5960 12374
rect 5908 12310 5960 12316
rect 5920 12170 5948 12310
rect 6104 12306 6132 15558
rect 6564 15502 6592 16730
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 6840 15502 6868 16594
rect 6932 16522 6960 16730
rect 7012 16720 7064 16726
rect 7012 16662 7064 16668
rect 6920 16516 6972 16522
rect 6920 16458 6972 16464
rect 7024 15502 7052 16662
rect 7116 16250 7144 19774
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7208 18630 7236 19654
rect 7196 18624 7248 18630
rect 7196 18566 7248 18572
rect 7300 17678 7328 24550
rect 7380 24132 7432 24138
rect 7380 24074 7432 24080
rect 7392 23730 7420 24074
rect 7484 23769 7512 25214
rect 7564 25152 7616 25158
rect 7564 25094 7616 25100
rect 7576 24886 7604 25094
rect 7564 24880 7616 24886
rect 7564 24822 7616 24828
rect 7668 24698 7696 29990
rect 7748 29232 7800 29238
rect 7748 29174 7800 29180
rect 7760 29102 7788 29174
rect 7748 29096 7800 29102
rect 7748 29038 7800 29044
rect 7760 27402 7788 29038
rect 7748 27396 7800 27402
rect 7748 27338 7800 27344
rect 7576 24670 7696 24698
rect 7470 23760 7526 23769
rect 7380 23724 7432 23730
rect 7470 23695 7526 23704
rect 7380 23666 7432 23672
rect 7288 17672 7340 17678
rect 7288 17614 7340 17620
rect 7288 17536 7340 17542
rect 7288 17478 7340 17484
rect 7300 16794 7328 17478
rect 7392 17270 7420 23666
rect 7470 21040 7526 21049
rect 7470 20975 7472 20984
rect 7524 20975 7526 20984
rect 7472 20946 7524 20952
rect 7472 19440 7524 19446
rect 7472 19382 7524 19388
rect 7484 18154 7512 19382
rect 7576 18154 7604 24670
rect 7656 24336 7708 24342
rect 7656 24278 7708 24284
rect 7668 21570 7696 24278
rect 7760 22982 7788 27338
rect 7852 24342 7880 30058
rect 7944 27062 7972 37284
rect 8024 37266 8076 37272
rect 8484 37324 8536 37330
rect 8484 37266 8536 37272
rect 8668 37324 8720 37330
rect 8668 37266 8720 37272
rect 8392 37256 8444 37262
rect 8392 37198 8444 37204
rect 8024 37188 8076 37194
rect 8024 37130 8076 37136
rect 8036 36718 8064 37130
rect 8404 36922 8432 37198
rect 8484 37188 8536 37194
rect 8484 37130 8536 37136
rect 8392 36916 8444 36922
rect 8392 36858 8444 36864
rect 8496 36786 8524 37130
rect 8300 36780 8352 36786
rect 8300 36722 8352 36728
rect 8484 36780 8536 36786
rect 8484 36722 8536 36728
rect 8024 36712 8076 36718
rect 8024 36654 8076 36660
rect 8312 36258 8340 36722
rect 8220 36230 8432 36258
rect 8220 36174 8248 36230
rect 8208 36168 8260 36174
rect 8208 36110 8260 36116
rect 8024 35760 8076 35766
rect 8024 35702 8076 35708
rect 8036 35086 8064 35702
rect 8404 35630 8432 36230
rect 8392 35624 8444 35630
rect 8392 35566 8444 35572
rect 8496 35170 8524 36722
rect 8576 36372 8628 36378
rect 8576 36314 8628 36320
rect 8588 36242 8616 36314
rect 8576 36236 8628 36242
rect 8576 36178 8628 36184
rect 8576 35760 8628 35766
rect 8576 35702 8628 35708
rect 8404 35154 8524 35170
rect 8392 35148 8524 35154
rect 8444 35142 8524 35148
rect 8392 35090 8444 35096
rect 8024 35080 8076 35086
rect 8024 35022 8076 35028
rect 8208 35080 8260 35086
rect 8208 35022 8260 35028
rect 8116 35012 8168 35018
rect 8116 34954 8168 34960
rect 8024 31884 8076 31890
rect 8024 31826 8076 31832
rect 8036 30938 8064 31826
rect 8024 30932 8076 30938
rect 8024 30874 8076 30880
rect 7932 27056 7984 27062
rect 7932 26998 7984 27004
rect 7944 25362 7972 26998
rect 8024 26376 8076 26382
rect 8024 26318 8076 26324
rect 7932 25356 7984 25362
rect 7932 25298 7984 25304
rect 7930 24440 7986 24449
rect 8036 24410 8064 26318
rect 8128 25498 8156 34954
rect 8220 34678 8248 35022
rect 8496 34678 8524 35142
rect 8208 34672 8260 34678
rect 8208 34614 8260 34620
rect 8484 34672 8536 34678
rect 8484 34614 8536 34620
rect 8220 34066 8248 34614
rect 8588 34610 8616 35702
rect 8576 34604 8628 34610
rect 8576 34546 8628 34552
rect 8484 34536 8536 34542
rect 8484 34478 8536 34484
rect 8392 34468 8444 34474
rect 8392 34410 8444 34416
rect 8208 34060 8260 34066
rect 8208 34002 8260 34008
rect 8404 33522 8432 34410
rect 8496 33998 8524 34478
rect 8484 33992 8536 33998
rect 8484 33934 8536 33940
rect 8680 33930 8708 37266
rect 8864 37262 8892 37402
rect 8852 37256 8904 37262
rect 8852 37198 8904 37204
rect 8852 36780 8904 36786
rect 8852 36722 8904 36728
rect 8864 35834 8892 36722
rect 9048 35834 9076 37862
rect 9312 37810 9364 37816
rect 9128 37664 9180 37670
rect 9128 37606 9180 37612
rect 9140 37262 9168 37606
rect 9128 37256 9180 37262
rect 9128 37198 9180 37204
rect 9404 37256 9456 37262
rect 9404 37198 9456 37204
rect 9140 36854 9168 37198
rect 9128 36848 9180 36854
rect 9128 36790 9180 36796
rect 9416 36786 9444 37198
rect 9772 36916 9824 36922
rect 9772 36858 9824 36864
rect 9404 36780 9456 36786
rect 9404 36722 9456 36728
rect 9220 36644 9272 36650
rect 9220 36586 9272 36592
rect 9128 36576 9180 36582
rect 9128 36518 9180 36524
rect 9140 36174 9168 36518
rect 9232 36174 9260 36586
rect 9128 36168 9180 36174
rect 9126 36136 9128 36145
rect 9220 36168 9272 36174
rect 9180 36136 9182 36145
rect 9220 36110 9272 36116
rect 9126 36071 9182 36080
rect 8852 35828 8904 35834
rect 8852 35770 8904 35776
rect 9036 35828 9088 35834
rect 9036 35770 9088 35776
rect 9048 35698 9076 35770
rect 9416 35698 9444 36722
rect 9496 36304 9548 36310
rect 9496 36246 9548 36252
rect 9036 35692 9088 35698
rect 9036 35634 9088 35640
rect 9312 35692 9364 35698
rect 9312 35634 9364 35640
rect 9404 35692 9456 35698
rect 9404 35634 9456 35640
rect 9128 35488 9180 35494
rect 9128 35430 9180 35436
rect 9036 35216 9088 35222
rect 9036 35158 9088 35164
rect 8760 35148 8812 35154
rect 8760 35090 8812 35096
rect 8772 34202 8800 35090
rect 9048 35086 9076 35158
rect 9140 35086 9168 35430
rect 9324 35290 9352 35634
rect 9312 35284 9364 35290
rect 9312 35226 9364 35232
rect 9508 35170 9536 36246
rect 9680 36168 9732 36174
rect 9680 36110 9732 36116
rect 9692 35698 9720 36110
rect 9680 35692 9732 35698
rect 9680 35634 9732 35640
rect 9324 35142 9536 35170
rect 9036 35080 9088 35086
rect 9036 35022 9088 35028
rect 9128 35080 9180 35086
rect 9128 35022 9180 35028
rect 8944 34604 8996 34610
rect 8944 34546 8996 34552
rect 8760 34196 8812 34202
rect 8760 34138 8812 34144
rect 8772 33998 8800 34138
rect 8956 34134 8984 34546
rect 9048 34202 9076 35022
rect 9128 34400 9180 34406
rect 9128 34342 9180 34348
rect 9036 34196 9088 34202
rect 9036 34138 9088 34144
rect 8944 34128 8996 34134
rect 8944 34070 8996 34076
rect 8760 33992 8812 33998
rect 8760 33934 8812 33940
rect 8668 33924 8720 33930
rect 8668 33866 8720 33872
rect 8392 33516 8444 33522
rect 8392 33458 8444 33464
rect 8484 33516 8536 33522
rect 8484 33458 8536 33464
rect 8404 33114 8432 33458
rect 8392 33108 8444 33114
rect 8392 33050 8444 33056
rect 8404 32978 8432 33050
rect 8392 32972 8444 32978
rect 8392 32914 8444 32920
rect 8496 32609 8524 33458
rect 8680 33454 8708 33866
rect 8956 33454 8984 34070
rect 9048 33522 9076 34138
rect 9140 33998 9168 34342
rect 9128 33992 9180 33998
rect 9128 33934 9180 33940
rect 9036 33516 9088 33522
rect 9036 33458 9088 33464
rect 8668 33448 8720 33454
rect 8668 33390 8720 33396
rect 8944 33448 8996 33454
rect 8944 33390 8996 33396
rect 8668 32972 8720 32978
rect 8668 32914 8720 32920
rect 8482 32600 8538 32609
rect 8482 32535 8538 32544
rect 8576 32428 8628 32434
rect 8576 32370 8628 32376
rect 8208 31748 8260 31754
rect 8208 31690 8260 31696
rect 8220 30734 8248 31690
rect 8300 31680 8352 31686
rect 8300 31622 8352 31628
rect 8312 30802 8340 31622
rect 8392 31476 8444 31482
rect 8392 31418 8444 31424
rect 8404 30870 8432 31418
rect 8588 31414 8616 32370
rect 8680 32026 8708 32914
rect 8852 32496 8904 32502
rect 8852 32438 8904 32444
rect 8668 32020 8720 32026
rect 8668 31962 8720 31968
rect 8576 31408 8628 31414
rect 8576 31350 8628 31356
rect 8576 31272 8628 31278
rect 8576 31214 8628 31220
rect 8588 30938 8616 31214
rect 8680 31210 8708 31962
rect 8760 31748 8812 31754
rect 8760 31690 8812 31696
rect 8668 31204 8720 31210
rect 8668 31146 8720 31152
rect 8576 30932 8628 30938
rect 8576 30874 8628 30880
rect 8772 30870 8800 31690
rect 8392 30864 8444 30870
rect 8392 30806 8444 30812
rect 8760 30864 8812 30870
rect 8760 30806 8812 30812
rect 8300 30796 8352 30802
rect 8300 30738 8352 30744
rect 8208 30728 8260 30734
rect 8208 30670 8260 30676
rect 8576 30388 8628 30394
rect 8576 30330 8628 30336
rect 8484 28620 8536 28626
rect 8484 28562 8536 28568
rect 8300 28416 8352 28422
rect 8300 28358 8352 28364
rect 8208 26240 8260 26246
rect 8208 26182 8260 26188
rect 8312 26194 8340 28358
rect 8496 28014 8524 28562
rect 8484 28008 8536 28014
rect 8484 27950 8536 27956
rect 8392 27668 8444 27674
rect 8392 27610 8444 27616
rect 8404 27130 8432 27610
rect 8392 27124 8444 27130
rect 8392 27066 8444 27072
rect 8390 27024 8446 27033
rect 8390 26959 8446 26968
rect 8404 26382 8432 26959
rect 8496 26926 8524 27950
rect 8484 26920 8536 26926
rect 8484 26862 8536 26868
rect 8392 26376 8444 26382
rect 8392 26318 8444 26324
rect 8484 26376 8536 26382
rect 8484 26318 8536 26324
rect 8116 25492 8168 25498
rect 8116 25434 8168 25440
rect 8220 25265 8248 26182
rect 8312 26166 8432 26194
rect 8300 25288 8352 25294
rect 8206 25256 8262 25265
rect 8300 25230 8352 25236
rect 8206 25191 8262 25200
rect 8116 24608 8168 24614
rect 8116 24550 8168 24556
rect 8128 24410 8156 24550
rect 7930 24375 7986 24384
rect 8024 24404 8076 24410
rect 7840 24336 7892 24342
rect 7840 24278 7892 24284
rect 7840 24200 7892 24206
rect 7840 24142 7892 24148
rect 7852 23866 7880 24142
rect 7840 23860 7892 23866
rect 7840 23802 7892 23808
rect 7944 23730 7972 24375
rect 8024 24346 8076 24352
rect 8116 24404 8168 24410
rect 8116 24346 8168 24352
rect 8114 24304 8170 24313
rect 8114 24239 8170 24248
rect 7932 23724 7984 23730
rect 7932 23666 7984 23672
rect 8128 23662 8156 24239
rect 8220 23730 8248 25191
rect 8312 24342 8340 25230
rect 8404 25158 8432 26166
rect 8496 25906 8524 26318
rect 8588 26194 8616 30330
rect 8760 29028 8812 29034
rect 8760 28970 8812 28976
rect 8668 28960 8720 28966
rect 8668 28902 8720 28908
rect 8680 28558 8708 28902
rect 8668 28552 8720 28558
rect 8668 28494 8720 28500
rect 8772 28234 8800 28970
rect 8864 28422 8892 32438
rect 8956 31872 8984 33390
rect 9036 33312 9088 33318
rect 9036 33254 9088 33260
rect 9048 32026 9076 33254
rect 9220 33108 9272 33114
rect 9220 33050 9272 33056
rect 9232 32366 9260 33050
rect 9220 32360 9272 32366
rect 9220 32302 9272 32308
rect 9036 32020 9088 32026
rect 9036 31962 9088 31968
rect 8956 31844 9076 31872
rect 8944 31748 8996 31754
rect 8944 31690 8996 31696
rect 8956 31414 8984 31690
rect 9048 31686 9076 31844
rect 9036 31680 9088 31686
rect 9036 31622 9088 31628
rect 8944 31408 8996 31414
rect 8944 31350 8996 31356
rect 9128 30864 9180 30870
rect 9128 30806 9180 30812
rect 8852 28416 8904 28422
rect 8852 28358 8904 28364
rect 8772 28206 8892 28234
rect 8864 28014 8892 28206
rect 8852 28008 8904 28014
rect 8852 27950 8904 27956
rect 8760 26920 8812 26926
rect 8760 26862 8812 26868
rect 8588 26166 8708 26194
rect 8484 25900 8536 25906
rect 8484 25842 8536 25848
rect 8484 25356 8536 25362
rect 8484 25298 8536 25304
rect 8392 25152 8444 25158
rect 8390 25120 8392 25129
rect 8444 25120 8446 25129
rect 8390 25055 8446 25064
rect 8496 24954 8524 25298
rect 8484 24948 8536 24954
rect 8484 24890 8536 24896
rect 8300 24336 8352 24342
rect 8300 24278 8352 24284
rect 8392 24132 8444 24138
rect 8392 24074 8444 24080
rect 8208 23724 8260 23730
rect 8208 23666 8260 23672
rect 8116 23656 8168 23662
rect 8116 23598 8168 23604
rect 8300 23588 8352 23594
rect 8300 23530 8352 23536
rect 7840 23112 7892 23118
rect 7840 23054 7892 23060
rect 7748 22976 7800 22982
rect 7748 22918 7800 22924
rect 7760 21894 7788 22918
rect 7852 22438 7880 23054
rect 8116 22772 8168 22778
rect 8116 22714 8168 22720
rect 8024 22704 8076 22710
rect 8024 22646 8076 22652
rect 7840 22432 7892 22438
rect 7840 22374 7892 22380
rect 7852 22030 7880 22374
rect 7840 22024 7892 22030
rect 7840 21966 7892 21972
rect 7748 21888 7800 21894
rect 7748 21830 7800 21836
rect 7668 21542 7972 21570
rect 7656 21480 7708 21486
rect 7656 21422 7708 21428
rect 7668 21146 7696 21422
rect 7656 21140 7708 21146
rect 7656 21082 7708 21088
rect 7840 20052 7892 20058
rect 7840 19994 7892 20000
rect 7852 19854 7880 19994
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7668 18970 7696 19246
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 7748 18624 7800 18630
rect 7748 18566 7800 18572
rect 7760 18290 7788 18566
rect 7840 18352 7892 18358
rect 7840 18294 7892 18300
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 7472 18148 7524 18154
rect 7472 18090 7524 18096
rect 7564 18148 7616 18154
rect 7564 18090 7616 18096
rect 7472 17604 7524 17610
rect 7472 17546 7524 17552
rect 7380 17264 7432 17270
rect 7380 17206 7432 17212
rect 7484 17202 7512 17546
rect 7852 17270 7880 18294
rect 7840 17264 7892 17270
rect 7840 17206 7892 17212
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7288 16584 7340 16590
rect 7288 16526 7340 16532
rect 7300 16454 7328 16526
rect 7392 16522 7420 16934
rect 7576 16658 7604 16934
rect 7668 16794 7696 17070
rect 7656 16788 7708 16794
rect 7656 16730 7708 16736
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 7380 16516 7432 16522
rect 7380 16458 7432 16464
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7300 16250 7328 16390
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 6196 14498 6224 15438
rect 6276 15360 6328 15366
rect 6276 15302 6328 15308
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6288 14618 6316 15302
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6276 14612 6328 14618
rect 6276 14554 6328 14560
rect 6196 14470 6316 14498
rect 6472 14482 6500 14758
rect 6564 14482 6592 15302
rect 6840 15094 6868 15438
rect 7024 15094 7052 15438
rect 6828 15088 6880 15094
rect 6828 15030 6880 15036
rect 7012 15088 7064 15094
rect 7012 15030 7064 15036
rect 6840 14482 6868 15030
rect 7576 15026 7604 16594
rect 7656 16448 7708 16454
rect 7656 16390 7708 16396
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6932 14498 6960 14894
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 7024 14618 7052 14826
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 6196 12238 6224 12582
rect 6288 12374 6316 14470
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6828 14476 6880 14482
rect 6932 14470 7052 14498
rect 6828 14418 6880 14424
rect 6840 14346 6868 14418
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6460 13184 6512 13190
rect 6460 13126 6512 13132
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6380 12442 6408 12582
rect 6472 12442 6500 13126
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 6276 12368 6328 12374
rect 6276 12310 6328 12316
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5908 12164 5960 12170
rect 5908 12106 5960 12112
rect 5736 11898 5764 12106
rect 6288 11914 6316 12310
rect 6656 12238 6684 13262
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 6932 12850 6960 12922
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6736 12776 6788 12782
rect 6736 12718 6788 12724
rect 6826 12744 6882 12753
rect 6748 12238 6776 12718
rect 6826 12679 6882 12688
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6736 12232 6788 12238
rect 6736 12174 6788 12180
rect 6288 11898 6592 11914
rect 5724 11892 5776 11898
rect 6288 11892 6604 11898
rect 6288 11886 6552 11892
rect 5724 11834 5776 11840
rect 6552 11834 6604 11840
rect 5724 10736 5776 10742
rect 5724 10678 5776 10684
rect 5736 10305 5764 10678
rect 6564 10674 6592 11834
rect 6748 11762 6776 12174
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 5722 10296 5778 10305
rect 6380 10266 6408 10406
rect 5722 10231 5778 10240
rect 6368 10260 6420 10266
rect 5736 10198 5764 10231
rect 6368 10202 6420 10208
rect 5724 10192 5776 10198
rect 5724 10134 5776 10140
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 4712 8560 4764 8566
rect 4712 8502 4764 8508
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4724 7342 4752 8502
rect 5644 7954 5672 8570
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5736 8090 5764 8366
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 6472 7886 6500 8230
rect 6564 7954 6592 10610
rect 6748 10266 6776 10610
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6840 10146 6868 12679
rect 7024 12306 7052 14470
rect 7208 14414 7236 14758
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7116 14006 7144 14350
rect 7104 14000 7156 14006
rect 7104 13942 7156 13948
rect 7116 13716 7144 13942
rect 7300 13870 7328 14758
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7116 13688 7328 13716
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7116 12850 7144 13262
rect 7300 12850 7328 13688
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7300 12306 7328 12786
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7104 11280 7156 11286
rect 7104 11222 7156 11228
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6748 10118 6868 10146
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6656 8498 6684 8774
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6748 8090 6776 10118
rect 6828 9988 6880 9994
rect 6828 9930 6880 9936
rect 6840 9586 6868 9930
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6840 8498 6868 8978
rect 6932 8634 6960 10610
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 7024 9586 7052 10406
rect 7116 10062 7144 11222
rect 7392 10810 7420 14214
rect 7484 13394 7512 14758
rect 7562 14512 7618 14521
rect 7562 14447 7564 14456
rect 7616 14447 7618 14456
rect 7564 14418 7616 14424
rect 7564 14340 7616 14346
rect 7564 14282 7616 14288
rect 7576 14074 7604 14282
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 7484 13258 7512 13330
rect 7472 13252 7524 13258
rect 7472 13194 7524 13200
rect 7472 12912 7524 12918
rect 7470 12880 7472 12889
rect 7524 12880 7526 12889
rect 7470 12815 7526 12824
rect 7564 12708 7616 12714
rect 7564 12650 7616 12656
rect 7576 12238 7604 12650
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7484 10674 7512 12038
rect 7668 11830 7696 16390
rect 7852 15162 7880 17206
rect 7944 16726 7972 21542
rect 8036 20058 8064 22646
rect 8128 22030 8156 22714
rect 8206 22400 8262 22409
rect 8206 22335 8262 22344
rect 8220 22166 8248 22335
rect 8208 22160 8260 22166
rect 8208 22102 8260 22108
rect 8116 22024 8168 22030
rect 8116 21966 8168 21972
rect 8128 20369 8156 21966
rect 8312 21962 8340 23530
rect 8404 23254 8432 24074
rect 8392 23248 8444 23254
rect 8392 23190 8444 23196
rect 8496 22094 8524 24890
rect 8680 24070 8708 26166
rect 8576 24064 8628 24070
rect 8668 24064 8720 24070
rect 8576 24006 8628 24012
rect 8666 24032 8668 24041
rect 8720 24032 8722 24041
rect 8588 23769 8616 24006
rect 8666 23967 8722 23976
rect 8666 23896 8722 23905
rect 8666 23831 8722 23840
rect 8574 23760 8630 23769
rect 8680 23730 8708 23831
rect 8574 23695 8630 23704
rect 8668 23724 8720 23730
rect 8668 23666 8720 23672
rect 8576 23520 8628 23526
rect 8576 23462 8628 23468
rect 8588 22642 8616 23462
rect 8576 22636 8628 22642
rect 8576 22578 8628 22584
rect 8576 22500 8628 22506
rect 8576 22442 8628 22448
rect 8588 22234 8616 22442
rect 8576 22228 8628 22234
rect 8576 22170 8628 22176
rect 8404 22066 8524 22094
rect 8300 21956 8352 21962
rect 8300 21898 8352 21904
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 8220 21554 8248 21830
rect 8208 21548 8260 21554
rect 8208 21490 8260 21496
rect 8206 21040 8262 21049
rect 8206 20975 8262 20984
rect 8220 20806 8248 20975
rect 8312 20806 8340 21898
rect 8404 21486 8432 22066
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 8392 21480 8444 21486
rect 8392 21422 8444 21428
rect 8496 21078 8524 21966
rect 8576 21956 8628 21962
rect 8576 21898 8628 21904
rect 8588 21690 8616 21898
rect 8576 21684 8628 21690
rect 8576 21626 8628 21632
rect 8588 21554 8616 21626
rect 8576 21548 8628 21554
rect 8576 21490 8628 21496
rect 8680 21434 8708 23666
rect 8772 22273 8800 26862
rect 8864 23730 8892 27950
rect 8942 26616 8998 26625
rect 8942 26551 8998 26560
rect 8956 26518 8984 26551
rect 8944 26512 8996 26518
rect 8944 26454 8996 26460
rect 9036 26308 9088 26314
rect 9036 26250 9088 26256
rect 9048 25294 9076 26250
rect 9140 25362 9168 30806
rect 9232 26042 9260 32302
rect 9324 26586 9352 35142
rect 9404 35080 9456 35086
rect 9404 35022 9456 35028
rect 9416 34746 9444 35022
rect 9404 34740 9456 34746
rect 9404 34682 9456 34688
rect 9588 34604 9640 34610
rect 9588 34546 9640 34552
rect 9600 33522 9628 34546
rect 9784 34474 9812 36858
rect 9968 36242 9996 38694
rect 10152 38332 10180 38694
rect 10244 38554 10272 38898
rect 10508 38888 10560 38894
rect 10508 38830 10560 38836
rect 10520 38554 10548 38830
rect 10600 38752 10652 38758
rect 10600 38694 10652 38700
rect 10232 38548 10284 38554
rect 10232 38490 10284 38496
rect 10508 38548 10560 38554
rect 10508 38490 10560 38496
rect 10232 38344 10284 38350
rect 10152 38304 10232 38332
rect 10232 38286 10284 38292
rect 9956 36236 10008 36242
rect 9956 36178 10008 36184
rect 10140 36100 10192 36106
rect 10140 36042 10192 36048
rect 10152 36009 10180 36042
rect 10138 36000 10194 36009
rect 10138 35935 10194 35944
rect 10140 35488 10192 35494
rect 10244 35476 10272 38286
rect 10612 36854 10640 38694
rect 10888 36922 10916 39034
rect 11072 38962 11100 39238
rect 11060 38956 11112 38962
rect 11060 38898 11112 38904
rect 11256 38214 11284 39374
rect 11532 38554 11560 39374
rect 11992 39302 12020 39578
rect 12072 39568 12124 39574
rect 12072 39510 12124 39516
rect 11612 39296 11664 39302
rect 11612 39238 11664 39244
rect 11980 39296 12032 39302
rect 11980 39238 12032 39244
rect 11624 39030 11652 39238
rect 11992 39098 12020 39238
rect 12084 39098 12112 39510
rect 12176 39438 12204 39782
rect 12164 39432 12216 39438
rect 12164 39374 12216 39380
rect 11980 39092 12032 39098
rect 11980 39034 12032 39040
rect 12072 39092 12124 39098
rect 12072 39034 12124 39040
rect 11612 39024 11664 39030
rect 11612 38966 11664 38972
rect 12268 38962 12296 39918
rect 12532 39840 12584 39846
rect 12532 39782 12584 39788
rect 12256 38956 12308 38962
rect 12256 38898 12308 38904
rect 11520 38548 11572 38554
rect 11520 38490 11572 38496
rect 12268 38350 12296 38898
rect 12440 38888 12492 38894
rect 12440 38830 12492 38836
rect 11336 38344 11388 38350
rect 11336 38286 11388 38292
rect 12256 38344 12308 38350
rect 12256 38286 12308 38292
rect 11244 38208 11296 38214
rect 11244 38150 11296 38156
rect 10876 36916 10928 36922
rect 10876 36858 10928 36864
rect 10600 36848 10652 36854
rect 10600 36790 10652 36796
rect 10692 36780 10744 36786
rect 10692 36722 10744 36728
rect 10600 36576 10652 36582
rect 10600 36518 10652 36524
rect 10612 36106 10640 36518
rect 10704 36394 10732 36722
rect 10704 36366 10824 36394
rect 10692 36236 10744 36242
rect 10692 36178 10744 36184
rect 10600 36100 10652 36106
rect 10600 36042 10652 36048
rect 10416 36032 10468 36038
rect 10416 35974 10468 35980
rect 10428 35630 10456 35974
rect 10600 35760 10652 35766
rect 10506 35728 10562 35737
rect 10600 35702 10652 35708
rect 10506 35663 10508 35672
rect 10560 35663 10562 35672
rect 10508 35634 10560 35640
rect 10416 35624 10468 35630
rect 10416 35566 10468 35572
rect 10612 35494 10640 35702
rect 10600 35488 10652 35494
rect 10244 35448 10456 35476
rect 10140 35430 10192 35436
rect 10152 35057 10180 35430
rect 10138 35048 10194 35057
rect 10138 34983 10194 34992
rect 10152 34610 10180 34983
rect 10140 34604 10192 34610
rect 10140 34546 10192 34552
rect 10324 34536 10376 34542
rect 10324 34478 10376 34484
rect 9772 34468 9824 34474
rect 9772 34410 9824 34416
rect 10140 34400 10192 34406
rect 10140 34342 10192 34348
rect 10232 34400 10284 34406
rect 10232 34342 10284 34348
rect 9680 34196 9732 34202
rect 9680 34138 9732 34144
rect 9692 33998 9720 34138
rect 9680 33992 9732 33998
rect 9680 33934 9732 33940
rect 9692 33658 9720 33934
rect 10048 33924 10100 33930
rect 10048 33866 10100 33872
rect 9772 33856 9824 33862
rect 9772 33798 9824 33804
rect 9680 33652 9732 33658
rect 9680 33594 9732 33600
rect 9588 33516 9640 33522
rect 9588 33458 9640 33464
rect 9600 33114 9628 33458
rect 9784 33386 9812 33798
rect 10060 33522 10088 33866
rect 10048 33516 10100 33522
rect 10048 33458 10100 33464
rect 10152 33454 10180 34342
rect 10244 33522 10272 34342
rect 10336 33998 10364 34478
rect 10324 33992 10376 33998
rect 10324 33934 10376 33940
rect 10336 33658 10364 33934
rect 10324 33652 10376 33658
rect 10324 33594 10376 33600
rect 10232 33516 10284 33522
rect 10232 33458 10284 33464
rect 10140 33448 10192 33454
rect 10140 33390 10192 33396
rect 9772 33380 9824 33386
rect 9772 33322 9824 33328
rect 9588 33108 9640 33114
rect 9588 33050 9640 33056
rect 9956 31340 10008 31346
rect 9956 31282 10008 31288
rect 9404 31272 9456 31278
rect 9404 31214 9456 31220
rect 9416 30326 9444 31214
rect 9864 31204 9916 31210
rect 9864 31146 9916 31152
rect 9588 31136 9640 31142
rect 9588 31078 9640 31084
rect 9404 30320 9456 30326
rect 9404 30262 9456 30268
rect 9416 29714 9444 30262
rect 9404 29708 9456 29714
rect 9404 29650 9456 29656
rect 9416 29084 9444 29650
rect 9496 29504 9548 29510
rect 9496 29446 9548 29452
rect 9508 29238 9536 29446
rect 9496 29232 9548 29238
rect 9496 29174 9548 29180
rect 9496 29096 9548 29102
rect 9416 29056 9496 29084
rect 9496 29038 9548 29044
rect 9496 28960 9548 28966
rect 9496 28902 9548 28908
rect 9508 27384 9536 28902
rect 9600 27538 9628 31078
rect 9680 30796 9732 30802
rect 9680 30738 9732 30744
rect 9692 29578 9720 30738
rect 9876 30190 9904 31146
rect 9968 31142 9996 31282
rect 9956 31136 10008 31142
rect 9956 31078 10008 31084
rect 10324 30592 10376 30598
rect 10324 30534 10376 30540
rect 9864 30184 9916 30190
rect 9864 30126 9916 30132
rect 9772 30048 9824 30054
rect 9772 29990 9824 29996
rect 9680 29572 9732 29578
rect 9680 29514 9732 29520
rect 9784 29238 9812 29990
rect 9956 29640 10008 29646
rect 9956 29582 10008 29588
rect 9772 29232 9824 29238
rect 9772 29174 9824 29180
rect 9968 29034 9996 29582
rect 9956 29028 10008 29034
rect 9956 28970 10008 28976
rect 9680 28960 9732 28966
rect 9680 28902 9732 28908
rect 9692 28558 9720 28902
rect 9864 28688 9916 28694
rect 9864 28630 9916 28636
rect 9680 28552 9732 28558
rect 9680 28494 9732 28500
rect 9876 28082 9904 28630
rect 9864 28076 9916 28082
rect 9864 28018 9916 28024
rect 9876 27985 9904 28018
rect 9862 27976 9918 27985
rect 9680 27940 9732 27946
rect 9862 27911 9918 27920
rect 9680 27882 9732 27888
rect 9588 27532 9640 27538
rect 9588 27474 9640 27480
rect 9508 27356 9628 27384
rect 9496 26852 9548 26858
rect 9496 26794 9548 26800
rect 9312 26580 9364 26586
rect 9312 26522 9364 26528
rect 9324 26382 9352 26522
rect 9508 26450 9536 26794
rect 9496 26444 9548 26450
rect 9496 26386 9548 26392
rect 9312 26376 9364 26382
rect 9312 26318 9364 26324
rect 9496 26308 9548 26314
rect 9496 26250 9548 26256
rect 9220 26036 9272 26042
rect 9220 25978 9272 25984
rect 9128 25356 9180 25362
rect 9128 25298 9180 25304
rect 9036 25288 9088 25294
rect 9036 25230 9088 25236
rect 9128 24608 9180 24614
rect 9034 24576 9090 24585
rect 9128 24550 9180 24556
rect 9034 24511 9090 24520
rect 9048 24342 9076 24511
rect 9036 24336 9088 24342
rect 9036 24278 9088 24284
rect 8942 24032 8998 24041
rect 8942 23967 8998 23976
rect 8852 23724 8904 23730
rect 8852 23666 8904 23672
rect 8956 23338 8984 23967
rect 9140 23769 9168 24550
rect 9232 24313 9260 25978
rect 9404 25288 9456 25294
rect 9404 25230 9456 25236
rect 9416 24886 9444 25230
rect 9404 24880 9456 24886
rect 9404 24822 9456 24828
rect 9312 24812 9364 24818
rect 9312 24754 9364 24760
rect 9324 24449 9352 24754
rect 9310 24440 9366 24449
rect 9310 24375 9366 24384
rect 9324 24342 9352 24375
rect 9312 24336 9364 24342
rect 9218 24304 9274 24313
rect 9312 24278 9364 24284
rect 9218 24239 9274 24248
rect 9220 24200 9272 24206
rect 9220 24142 9272 24148
rect 9126 23760 9182 23769
rect 9126 23695 9182 23704
rect 8864 23310 8984 23338
rect 9232 23322 9260 24142
rect 9312 24132 9364 24138
rect 9312 24074 9364 24080
rect 9220 23316 9272 23322
rect 8758 22264 8814 22273
rect 8758 22199 8814 22208
rect 8588 21406 8708 21434
rect 8484 21072 8536 21078
rect 8484 21014 8536 21020
rect 8588 20874 8616 21406
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8680 20942 8708 21286
rect 8668 20936 8720 20942
rect 8668 20878 8720 20884
rect 8576 20868 8628 20874
rect 8576 20810 8628 20816
rect 8208 20800 8260 20806
rect 8208 20742 8260 20748
rect 8300 20800 8352 20806
rect 8300 20742 8352 20748
rect 8114 20360 8170 20369
rect 8114 20295 8170 20304
rect 8024 20052 8076 20058
rect 8024 19994 8076 20000
rect 8116 19712 8168 19718
rect 8116 19654 8168 19660
rect 8128 18766 8156 19654
rect 8116 18760 8168 18766
rect 8116 18702 8168 18708
rect 8116 18624 8168 18630
rect 8220 18612 8248 20742
rect 8588 20641 8616 20810
rect 8574 20632 8630 20641
rect 8574 20567 8630 20576
rect 8576 20392 8628 20398
rect 8576 20334 8628 20340
rect 8588 19514 8616 20334
rect 8668 19916 8720 19922
rect 8668 19858 8720 19864
rect 8680 19514 8708 19858
rect 8576 19508 8628 19514
rect 8576 19450 8628 19456
rect 8668 19508 8720 19514
rect 8668 19450 8720 19456
rect 8588 19378 8616 19450
rect 8576 19372 8628 19378
rect 8864 19334 8892 23310
rect 9220 23258 9272 23264
rect 8944 23248 8996 23254
rect 8944 23190 8996 23196
rect 8956 23118 8984 23190
rect 8944 23112 8996 23118
rect 8944 23054 8996 23060
rect 9324 22778 9352 24074
rect 9416 23730 9444 24822
rect 9508 24818 9536 26250
rect 9496 24812 9548 24818
rect 9496 24754 9548 24760
rect 9496 24676 9548 24682
rect 9496 24618 9548 24624
rect 9404 23724 9456 23730
rect 9404 23666 9456 23672
rect 9508 23322 9536 24618
rect 9496 23316 9548 23322
rect 9496 23258 9548 23264
rect 9508 22982 9536 23258
rect 9496 22976 9548 22982
rect 9496 22918 9548 22924
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 9496 22568 9548 22574
rect 9496 22510 9548 22516
rect 8944 22432 8996 22438
rect 9036 22432 9088 22438
rect 8944 22374 8996 22380
rect 9034 22400 9036 22409
rect 9088 22400 9090 22409
rect 8956 22234 8984 22374
rect 9034 22335 9090 22344
rect 8944 22228 8996 22234
rect 8944 22170 8996 22176
rect 9508 21894 9536 22510
rect 9600 22438 9628 27356
rect 9692 27130 9720 27882
rect 9864 27464 9916 27470
rect 9864 27406 9916 27412
rect 9772 27396 9824 27402
rect 9772 27338 9824 27344
rect 9784 27130 9812 27338
rect 9680 27124 9732 27130
rect 9680 27066 9732 27072
rect 9772 27124 9824 27130
rect 9772 27066 9824 27072
rect 9692 25242 9720 27066
rect 9772 26920 9824 26926
rect 9876 26908 9904 27406
rect 9824 26880 9904 26908
rect 9772 26862 9824 26868
rect 9772 26784 9824 26790
rect 9772 26726 9824 26732
rect 9784 26246 9812 26726
rect 9772 26240 9824 26246
rect 9772 26182 9824 26188
rect 9692 25214 9904 25242
rect 9772 25152 9824 25158
rect 9772 25094 9824 25100
rect 9784 24818 9812 25094
rect 9680 24812 9732 24818
rect 9680 24754 9732 24760
rect 9772 24812 9824 24818
rect 9772 24754 9824 24760
rect 9692 24410 9720 24754
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 9678 24304 9734 24313
rect 9678 24239 9734 24248
rect 9588 22432 9640 22438
rect 9588 22374 9640 22380
rect 9586 22264 9642 22273
rect 9586 22199 9642 22208
rect 9496 21888 9548 21894
rect 9496 21830 9548 21836
rect 9496 20528 9548 20534
rect 9496 20470 9548 20476
rect 9312 20392 9364 20398
rect 9312 20334 9364 20340
rect 9324 20058 9352 20334
rect 9312 20052 9364 20058
rect 9312 19994 9364 20000
rect 9508 19446 9536 20470
rect 9496 19440 9548 19446
rect 9496 19382 9548 19388
rect 8576 19314 8628 19320
rect 8772 19306 8892 19334
rect 8772 18766 8800 19306
rect 9496 19304 9548 19310
rect 9496 19246 9548 19252
rect 9508 18970 9536 19246
rect 9496 18964 9548 18970
rect 9496 18906 9548 18912
rect 8760 18760 8812 18766
rect 8760 18702 8812 18708
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 8168 18584 8248 18612
rect 8116 18566 8168 18572
rect 8128 18426 8156 18566
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 8758 17912 8814 17921
rect 8758 17847 8814 17856
rect 8024 17740 8076 17746
rect 8024 17682 8076 17688
rect 8036 17202 8064 17682
rect 8772 17678 8800 17847
rect 9232 17678 9260 18022
rect 8760 17672 8812 17678
rect 8760 17614 8812 17620
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 9416 17542 9444 18702
rect 9600 17814 9628 22199
rect 9588 17808 9640 17814
rect 9588 17750 9640 17756
rect 9692 17678 9720 24239
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 9784 23186 9812 23666
rect 9772 23180 9824 23186
rect 9772 23122 9824 23128
rect 9770 23080 9826 23089
rect 9770 23015 9772 23024
rect 9824 23015 9826 23024
rect 9772 22986 9824 22992
rect 9876 21486 9904 25214
rect 9968 22982 9996 28970
rect 10232 28416 10284 28422
rect 10232 28358 10284 28364
rect 10244 27130 10272 28358
rect 10232 27124 10284 27130
rect 10232 27066 10284 27072
rect 10232 26988 10284 26994
rect 10232 26930 10284 26936
rect 10140 26852 10192 26858
rect 10140 26794 10192 26800
rect 10048 26308 10100 26314
rect 10048 26250 10100 26256
rect 10060 25906 10088 26250
rect 10048 25900 10100 25906
rect 10048 25842 10100 25848
rect 9956 22976 10008 22982
rect 9956 22918 10008 22924
rect 10048 22432 10100 22438
rect 10048 22374 10100 22380
rect 10060 21690 10088 22374
rect 10048 21684 10100 21690
rect 10048 21626 10100 21632
rect 9864 21480 9916 21486
rect 9784 21440 9864 21468
rect 9784 19922 9812 21440
rect 9864 21422 9916 21428
rect 10152 21010 10180 26794
rect 10244 26518 10272 26930
rect 10232 26512 10284 26518
rect 10232 26454 10284 26460
rect 10336 26466 10364 30534
rect 10428 29050 10456 35448
rect 10600 35430 10652 35436
rect 10600 34604 10652 34610
rect 10600 34546 10652 34552
rect 10612 34202 10640 34546
rect 10704 34542 10732 36178
rect 10796 34950 10824 36366
rect 10888 36106 10916 36858
rect 11152 36780 11204 36786
rect 11152 36722 11204 36728
rect 10876 36100 10928 36106
rect 10876 36042 10928 36048
rect 11058 36000 11114 36009
rect 11058 35935 11114 35944
rect 11072 35834 11100 35935
rect 11060 35828 11112 35834
rect 11060 35770 11112 35776
rect 10966 35728 11022 35737
rect 10966 35663 10968 35672
rect 11020 35663 11022 35672
rect 10968 35634 11020 35640
rect 11164 35562 11192 36722
rect 11348 36718 11376 38286
rect 12452 38282 12480 38830
rect 12440 38276 12492 38282
rect 12440 38218 12492 38224
rect 12164 37324 12216 37330
rect 12164 37266 12216 37272
rect 12440 37324 12492 37330
rect 12440 37266 12492 37272
rect 11704 36916 11756 36922
rect 11704 36858 11756 36864
rect 11336 36712 11388 36718
rect 11336 36654 11388 36660
rect 11520 36576 11572 36582
rect 11520 36518 11572 36524
rect 11532 36258 11560 36518
rect 11532 36242 11652 36258
rect 11532 36236 11664 36242
rect 11532 36230 11612 36236
rect 11532 35766 11560 36230
rect 11612 36178 11664 36184
rect 11612 36032 11664 36038
rect 11716 35986 11744 36858
rect 11980 36712 12032 36718
rect 11980 36654 12032 36660
rect 11888 36236 11940 36242
rect 11888 36178 11940 36184
rect 11664 35980 11744 35986
rect 11612 35974 11744 35980
rect 11624 35958 11744 35974
rect 11520 35760 11572 35766
rect 11520 35702 11572 35708
rect 11716 35698 11744 35958
rect 11900 35834 11928 36178
rect 11992 36174 12020 36654
rect 12176 36378 12204 37266
rect 12348 37256 12400 37262
rect 12348 37198 12400 37204
rect 12256 37120 12308 37126
rect 12256 37062 12308 37068
rect 12268 36718 12296 37062
rect 12360 36922 12388 37198
rect 12348 36916 12400 36922
rect 12348 36858 12400 36864
rect 12256 36712 12308 36718
rect 12256 36654 12308 36660
rect 12164 36372 12216 36378
rect 12164 36314 12216 36320
rect 12452 36258 12480 37266
rect 12544 37262 12572 39782
rect 12992 39296 13044 39302
rect 12992 39238 13044 39244
rect 13004 38418 13032 39238
rect 13464 38554 13492 40054
rect 15028 40050 15056 40530
rect 15752 40520 15804 40526
rect 15752 40462 15804 40468
rect 16396 40520 16448 40526
rect 16396 40462 16448 40468
rect 16580 40520 16632 40526
rect 16580 40462 16632 40468
rect 15476 40180 15528 40186
rect 15476 40122 15528 40128
rect 13636 40044 13688 40050
rect 13636 39986 13688 39992
rect 15016 40044 15068 40050
rect 15016 39986 15068 39992
rect 13648 39506 13676 39986
rect 14464 39976 14516 39982
rect 14464 39918 14516 39924
rect 14280 39908 14332 39914
rect 14280 39850 14332 39856
rect 13636 39500 13688 39506
rect 13636 39442 13688 39448
rect 13452 38548 13504 38554
rect 13452 38490 13504 38496
rect 13464 38418 13492 38490
rect 12992 38412 13044 38418
rect 12992 38354 13044 38360
rect 13452 38412 13504 38418
rect 13452 38354 13504 38360
rect 12624 38344 12676 38350
rect 12624 38286 12676 38292
rect 13176 38344 13228 38350
rect 13176 38286 13228 38292
rect 12636 37466 12664 38286
rect 12808 38208 12860 38214
rect 12808 38150 12860 38156
rect 12820 38010 12848 38150
rect 13188 38010 13216 38286
rect 13268 38208 13320 38214
rect 13268 38150 13320 38156
rect 12808 38004 12860 38010
rect 12808 37946 12860 37952
rect 13176 38004 13228 38010
rect 13176 37946 13228 37952
rect 13280 37942 13308 38150
rect 13268 37936 13320 37942
rect 13268 37878 13320 37884
rect 13728 37664 13780 37670
rect 13728 37606 13780 37612
rect 12624 37460 12676 37466
rect 12624 37402 12676 37408
rect 13740 37380 13768 37606
rect 13740 37352 13860 37380
rect 12532 37256 12584 37262
rect 12532 37198 12584 37204
rect 12624 37256 12676 37262
rect 12624 37198 12676 37204
rect 12636 36922 12664 37198
rect 13832 37194 13860 37352
rect 14188 37256 14240 37262
rect 14188 37198 14240 37204
rect 13820 37188 13872 37194
rect 13820 37130 13872 37136
rect 12624 36916 12676 36922
rect 12624 36858 12676 36864
rect 12716 36848 12768 36854
rect 12716 36790 12768 36796
rect 13176 36848 13228 36854
rect 13176 36790 13228 36796
rect 12452 36230 12572 36258
rect 11980 36168 12032 36174
rect 11980 36110 12032 36116
rect 12440 36100 12492 36106
rect 12440 36042 12492 36048
rect 11888 35828 11940 35834
rect 11888 35770 11940 35776
rect 12452 35698 12480 36042
rect 12544 35834 12572 36230
rect 12728 36174 12756 36790
rect 13084 36780 13136 36786
rect 13084 36722 13136 36728
rect 12900 36644 12952 36650
rect 12900 36586 12952 36592
rect 12716 36168 12768 36174
rect 12716 36110 12768 36116
rect 12532 35828 12584 35834
rect 12532 35770 12584 35776
rect 11704 35692 11756 35698
rect 11704 35634 11756 35640
rect 12440 35692 12492 35698
rect 12440 35634 12492 35640
rect 12808 35692 12860 35698
rect 12808 35634 12860 35640
rect 11152 35556 11204 35562
rect 11152 35498 11204 35504
rect 11244 35488 11296 35494
rect 11244 35430 11296 35436
rect 11256 35222 11284 35430
rect 11244 35216 11296 35222
rect 11244 35158 11296 35164
rect 10784 34944 10836 34950
rect 10784 34886 10836 34892
rect 10796 34610 10824 34886
rect 11256 34610 11284 35158
rect 12256 35080 12308 35086
rect 12256 35022 12308 35028
rect 12440 35080 12492 35086
rect 12440 35022 12492 35028
rect 11888 35012 11940 35018
rect 11888 34954 11940 34960
rect 11336 34944 11388 34950
rect 11336 34886 11388 34892
rect 11348 34610 11376 34886
rect 11428 34672 11480 34678
rect 11428 34614 11480 34620
rect 10784 34604 10836 34610
rect 10784 34546 10836 34552
rect 11060 34604 11112 34610
rect 11060 34546 11112 34552
rect 11244 34604 11296 34610
rect 11244 34546 11296 34552
rect 11336 34604 11388 34610
rect 11336 34546 11388 34552
rect 10692 34536 10744 34542
rect 10692 34478 10744 34484
rect 10968 34468 11020 34474
rect 10968 34410 11020 34416
rect 10980 34202 11008 34410
rect 10600 34196 10652 34202
rect 10600 34138 10652 34144
rect 10968 34196 11020 34202
rect 10968 34138 11020 34144
rect 10600 32904 10652 32910
rect 11072 32892 11100 34546
rect 11440 34490 11468 34614
rect 11900 34610 11928 34954
rect 11888 34604 11940 34610
rect 11888 34546 11940 34552
rect 11348 34462 11468 34490
rect 11348 33998 11376 34462
rect 11704 34400 11756 34406
rect 11704 34342 11756 34348
rect 12072 34400 12124 34406
rect 12072 34342 12124 34348
rect 11716 33998 11744 34342
rect 12084 34066 12112 34342
rect 12268 34202 12296 35022
rect 12348 34944 12400 34950
rect 12348 34886 12400 34892
rect 12256 34196 12308 34202
rect 12256 34138 12308 34144
rect 12360 34066 12388 34886
rect 12452 34202 12480 35022
rect 12440 34196 12492 34202
rect 12440 34138 12492 34144
rect 12072 34060 12124 34066
rect 12072 34002 12124 34008
rect 12348 34060 12400 34066
rect 12348 34002 12400 34008
rect 11152 33992 11204 33998
rect 11152 33934 11204 33940
rect 11336 33992 11388 33998
rect 11336 33934 11388 33940
rect 11704 33992 11756 33998
rect 11704 33934 11756 33940
rect 11164 33386 11192 33934
rect 11152 33380 11204 33386
rect 11152 33322 11204 33328
rect 11072 32864 11192 32892
rect 10600 32846 10652 32852
rect 10508 31680 10560 31686
rect 10508 31622 10560 31628
rect 10520 30870 10548 31622
rect 10508 30864 10560 30870
rect 10508 30806 10560 30812
rect 10612 30598 10640 32846
rect 11060 32768 11112 32774
rect 11060 32710 11112 32716
rect 10968 32360 11020 32366
rect 10968 32302 11020 32308
rect 10980 32026 11008 32302
rect 11072 32026 11100 32710
rect 10968 32020 11020 32026
rect 10968 31962 11020 31968
rect 11060 32020 11112 32026
rect 11060 31962 11112 31968
rect 11164 31906 11192 32864
rect 10888 31878 11192 31906
rect 10888 31482 10916 31878
rect 11244 31816 11296 31822
rect 10966 31784 11022 31793
rect 11244 31758 11296 31764
rect 10966 31719 11022 31728
rect 11152 31748 11204 31754
rect 10980 31482 11008 31719
rect 11152 31690 11204 31696
rect 11164 31657 11192 31690
rect 11150 31648 11206 31657
rect 11150 31583 11206 31592
rect 10876 31476 10928 31482
rect 10876 31418 10928 31424
rect 10968 31476 11020 31482
rect 10968 31418 11020 31424
rect 10784 31340 10836 31346
rect 10784 31282 10836 31288
rect 10876 31340 10928 31346
rect 10876 31282 10928 31288
rect 10692 31272 10744 31278
rect 10692 31214 10744 31220
rect 10704 30734 10732 31214
rect 10796 30938 10824 31282
rect 10784 30932 10836 30938
rect 10784 30874 10836 30880
rect 10692 30728 10744 30734
rect 10692 30670 10744 30676
rect 10600 30592 10652 30598
rect 10600 30534 10652 30540
rect 10704 30394 10732 30670
rect 10692 30388 10744 30394
rect 10888 30376 10916 31282
rect 10980 31278 11008 31418
rect 11152 31408 11204 31414
rect 11152 31350 11204 31356
rect 10968 31272 11020 31278
rect 10968 31214 11020 31220
rect 11060 31272 11112 31278
rect 11060 31214 11112 31220
rect 10968 30864 11020 30870
rect 10968 30806 11020 30812
rect 10692 30330 10744 30336
rect 10796 30348 10916 30376
rect 10704 29782 10732 30330
rect 10692 29776 10744 29782
rect 10796 29753 10824 30348
rect 10876 30252 10928 30258
rect 10876 30194 10928 30200
rect 10692 29718 10744 29724
rect 10782 29744 10838 29753
rect 10782 29679 10784 29688
rect 10836 29679 10838 29688
rect 10784 29650 10836 29656
rect 10692 29640 10744 29646
rect 10690 29608 10692 29617
rect 10744 29608 10746 29617
rect 10690 29543 10746 29552
rect 10784 29096 10836 29102
rect 10428 29022 10548 29050
rect 10784 29038 10836 29044
rect 10416 28960 10468 28966
rect 10416 28902 10468 28908
rect 10428 28558 10456 28902
rect 10416 28552 10468 28558
rect 10416 28494 10468 28500
rect 10520 26994 10548 29022
rect 10692 28960 10744 28966
rect 10692 28902 10744 28908
rect 10704 28558 10732 28902
rect 10692 28552 10744 28558
rect 10692 28494 10744 28500
rect 10796 28490 10824 29038
rect 10784 28484 10836 28490
rect 10784 28426 10836 28432
rect 10692 27464 10744 27470
rect 10692 27406 10744 27412
rect 10704 27305 10732 27406
rect 10690 27296 10746 27305
rect 10690 27231 10746 27240
rect 10690 27160 10746 27169
rect 10690 27095 10746 27104
rect 10704 27062 10732 27095
rect 10692 27056 10744 27062
rect 10692 26998 10744 27004
rect 10508 26988 10560 26994
rect 10508 26930 10560 26936
rect 10520 26586 10548 26930
rect 10600 26920 10652 26926
rect 10652 26880 10732 26908
rect 10600 26862 10652 26868
rect 10600 26784 10652 26790
rect 10600 26726 10652 26732
rect 10612 26586 10640 26726
rect 10508 26580 10560 26586
rect 10508 26522 10560 26528
rect 10600 26580 10652 26586
rect 10600 26522 10652 26528
rect 10244 23361 10272 26454
rect 10336 26438 10548 26466
rect 10324 26376 10376 26382
rect 10324 26318 10376 26324
rect 10336 25702 10364 26318
rect 10324 25696 10376 25702
rect 10324 25638 10376 25644
rect 10230 23352 10286 23361
rect 10336 23322 10364 25638
rect 10414 24848 10470 24857
rect 10414 24783 10416 24792
rect 10468 24783 10470 24792
rect 10416 24754 10468 24760
rect 10416 24200 10468 24206
rect 10416 24142 10468 24148
rect 10428 23866 10456 24142
rect 10520 23866 10548 26438
rect 10600 24812 10652 24818
rect 10600 24754 10652 24760
rect 10612 24206 10640 24754
rect 10600 24200 10652 24206
rect 10600 24142 10652 24148
rect 10416 23860 10468 23866
rect 10416 23802 10468 23808
rect 10508 23860 10560 23866
rect 10508 23802 10560 23808
rect 10520 23730 10548 23802
rect 10704 23730 10732 26880
rect 10796 26586 10824 28426
rect 10888 27470 10916 30194
rect 10876 27464 10928 27470
rect 10876 27406 10928 27412
rect 10784 26580 10836 26586
rect 10784 26522 10836 26528
rect 10888 26518 10916 27406
rect 10980 27062 11008 30806
rect 11072 30734 11100 31214
rect 11060 30728 11112 30734
rect 11060 30670 11112 30676
rect 11060 29844 11112 29850
rect 11060 29786 11112 29792
rect 11072 29238 11100 29786
rect 11060 29232 11112 29238
rect 11060 29174 11112 29180
rect 11164 28082 11192 31350
rect 11256 31142 11284 31758
rect 11348 31414 11376 33934
rect 11716 33862 11744 33934
rect 11704 33856 11756 33862
rect 11704 33798 11756 33804
rect 12440 33040 12492 33046
rect 12440 32982 12492 32988
rect 11612 32428 11664 32434
rect 11612 32370 11664 32376
rect 11428 31748 11480 31754
rect 11428 31690 11480 31696
rect 11336 31408 11388 31414
rect 11336 31350 11388 31356
rect 11336 31272 11388 31278
rect 11336 31214 11388 31220
rect 11244 31136 11296 31142
rect 11244 31078 11296 31084
rect 11152 28076 11204 28082
rect 11152 28018 11204 28024
rect 11152 27464 11204 27470
rect 11152 27406 11204 27412
rect 11164 27334 11192 27406
rect 11152 27328 11204 27334
rect 11152 27270 11204 27276
rect 11256 27130 11284 31078
rect 11348 30938 11376 31214
rect 11336 30932 11388 30938
rect 11336 30874 11388 30880
rect 11348 30326 11376 30874
rect 11440 30734 11468 31690
rect 11624 31482 11652 32370
rect 11888 32360 11940 32366
rect 11888 32302 11940 32308
rect 11704 32020 11756 32026
rect 11704 31962 11756 31968
rect 11612 31476 11664 31482
rect 11612 31418 11664 31424
rect 11520 31136 11572 31142
rect 11520 31078 11572 31084
rect 11532 30802 11560 31078
rect 11520 30796 11572 30802
rect 11520 30738 11572 30744
rect 11428 30728 11480 30734
rect 11428 30670 11480 30676
rect 11624 30546 11652 31418
rect 11716 31346 11744 31962
rect 11900 31890 11928 32302
rect 12072 32292 12124 32298
rect 12072 32234 12124 32240
rect 11888 31884 11940 31890
rect 11888 31826 11940 31832
rect 11888 31680 11940 31686
rect 11888 31622 11940 31628
rect 11900 31414 11928 31622
rect 11888 31408 11940 31414
rect 11888 31350 11940 31356
rect 11704 31340 11756 31346
rect 11704 31282 11756 31288
rect 11900 30938 11928 31350
rect 12084 31346 12112 32234
rect 12452 32230 12480 32982
rect 12532 32904 12584 32910
rect 12532 32846 12584 32852
rect 12544 32570 12572 32846
rect 12532 32564 12584 32570
rect 12532 32506 12584 32512
rect 12544 32366 12572 32506
rect 12532 32360 12584 32366
rect 12532 32302 12584 32308
rect 12624 32360 12676 32366
rect 12624 32302 12676 32308
rect 12440 32224 12492 32230
rect 12440 32166 12492 32172
rect 12544 31958 12572 32302
rect 12532 31952 12584 31958
rect 12532 31894 12584 31900
rect 12256 31884 12308 31890
rect 12256 31826 12308 31832
rect 12164 31816 12216 31822
rect 12268 31793 12296 31826
rect 12164 31758 12216 31764
rect 12254 31784 12310 31793
rect 12176 31634 12204 31758
rect 12254 31719 12310 31728
rect 12254 31648 12310 31657
rect 12176 31606 12254 31634
rect 12254 31583 12310 31592
rect 12544 31414 12572 31894
rect 12532 31408 12584 31414
rect 12532 31350 12584 31356
rect 12072 31340 12124 31346
rect 12072 31282 12124 31288
rect 11888 30932 11940 30938
rect 11888 30874 11940 30880
rect 12164 30660 12216 30666
rect 12164 30602 12216 30608
rect 11440 30518 11652 30546
rect 11336 30320 11388 30326
rect 11336 30262 11388 30268
rect 11336 29640 11388 29646
rect 11336 29582 11388 29588
rect 11348 29306 11376 29582
rect 11336 29300 11388 29306
rect 11336 29242 11388 29248
rect 11336 29164 11388 29170
rect 11336 29106 11388 29112
rect 11348 29034 11376 29106
rect 11336 29028 11388 29034
rect 11336 28970 11388 28976
rect 11336 28076 11388 28082
rect 11336 28018 11388 28024
rect 11060 27124 11112 27130
rect 11060 27066 11112 27072
rect 11244 27124 11296 27130
rect 11244 27066 11296 27072
rect 10968 27056 11020 27062
rect 10968 26998 11020 27004
rect 10876 26512 10928 26518
rect 10876 26454 10928 26460
rect 10966 26480 11022 26489
rect 10966 26415 10968 26424
rect 11020 26415 11022 26424
rect 10968 26386 11020 26392
rect 11072 26314 11100 27066
rect 11348 27010 11376 28018
rect 11256 26982 11376 27010
rect 11152 26920 11204 26926
rect 11152 26862 11204 26868
rect 11164 26382 11192 26862
rect 11152 26376 11204 26382
rect 11152 26318 11204 26324
rect 11060 26308 11112 26314
rect 11060 26250 11112 26256
rect 11256 25294 11284 26982
rect 11336 26920 11388 26926
rect 11336 26862 11388 26868
rect 11348 26450 11376 26862
rect 11336 26444 11388 26450
rect 11336 26386 11388 26392
rect 11336 25492 11388 25498
rect 11336 25434 11388 25440
rect 11060 25288 11112 25294
rect 11060 25230 11112 25236
rect 11244 25288 11296 25294
rect 11244 25230 11296 25236
rect 10968 24880 11020 24886
rect 10968 24822 11020 24828
rect 10876 24812 10928 24818
rect 10876 24754 10928 24760
rect 10784 24676 10836 24682
rect 10784 24618 10836 24624
rect 10508 23724 10560 23730
rect 10508 23666 10560 23672
rect 10692 23724 10744 23730
rect 10692 23666 10744 23672
rect 10692 23588 10744 23594
rect 10692 23530 10744 23536
rect 10230 23287 10286 23296
rect 10324 23316 10376 23322
rect 10324 23258 10376 23264
rect 10508 23112 10560 23118
rect 10230 23080 10286 23089
rect 10230 23015 10286 23024
rect 10414 23080 10470 23089
rect 10704 23089 10732 23530
rect 10508 23054 10560 23060
rect 10690 23080 10746 23089
rect 10414 23015 10416 23024
rect 10244 22642 10272 23015
rect 10468 23015 10470 23024
rect 10416 22986 10468 22992
rect 10520 22710 10548 23054
rect 10690 23015 10746 23024
rect 10692 22976 10744 22982
rect 10692 22918 10744 22924
rect 10508 22704 10560 22710
rect 10508 22646 10560 22652
rect 10232 22636 10284 22642
rect 10232 22578 10284 22584
rect 10232 22500 10284 22506
rect 10232 22442 10284 22448
rect 10244 21146 10272 22442
rect 10506 22128 10562 22137
rect 10416 22092 10468 22098
rect 10468 22072 10506 22080
rect 10468 22063 10562 22072
rect 10468 22052 10548 22063
rect 10416 22034 10468 22040
rect 10520 21962 10548 22052
rect 10416 21956 10468 21962
rect 10416 21898 10468 21904
rect 10508 21956 10560 21962
rect 10508 21898 10560 21904
rect 10428 21690 10456 21898
rect 10416 21684 10468 21690
rect 10416 21626 10468 21632
rect 10506 21584 10562 21593
rect 10506 21519 10508 21528
rect 10560 21519 10562 21528
rect 10508 21490 10560 21496
rect 10232 21140 10284 21146
rect 10232 21082 10284 21088
rect 10508 21140 10560 21146
rect 10508 21082 10560 21088
rect 9864 21004 9916 21010
rect 9864 20946 9916 20952
rect 10140 21004 10192 21010
rect 10140 20946 10192 20952
rect 9876 20330 9904 20946
rect 10232 20936 10284 20942
rect 10232 20878 10284 20884
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 9864 20324 9916 20330
rect 9864 20266 9916 20272
rect 9876 19922 9904 20266
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9784 19334 9812 19858
rect 9968 19854 9996 20198
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 10060 19718 10088 20742
rect 10244 20058 10272 20878
rect 10232 20052 10284 20058
rect 10232 19994 10284 20000
rect 10416 19780 10468 19786
rect 10416 19722 10468 19728
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 10428 19514 10456 19722
rect 10416 19508 10468 19514
rect 10416 19450 10468 19456
rect 9784 19306 9996 19334
rect 9968 18630 9996 19306
rect 9864 18624 9916 18630
rect 9864 18566 9916 18572
rect 9956 18624 10008 18630
rect 9956 18566 10008 18572
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8852 17536 8904 17542
rect 8852 17478 8904 17484
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 8680 17202 8708 17478
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 7932 16720 7984 16726
rect 7932 16662 7984 16668
rect 8036 15502 8064 17138
rect 8116 16992 8168 16998
rect 8116 16934 8168 16940
rect 8128 16658 8156 16934
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8220 16522 8248 16730
rect 8208 16516 8260 16522
rect 8208 16458 8260 16464
rect 8220 16250 8248 16458
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 7932 15360 7984 15366
rect 7932 15302 7984 15308
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7944 15026 7972 15302
rect 8036 15026 8064 15438
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 8024 15020 8076 15026
rect 8024 14962 8076 14968
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 8022 14512 8078 14521
rect 8022 14447 8078 14456
rect 8036 13326 8064 14447
rect 8128 13462 8156 14758
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8116 13456 8168 13462
rect 8116 13398 8168 13404
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 8128 13274 8156 13398
rect 8220 13394 8248 14214
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 7760 13190 7788 13262
rect 8128 13258 8248 13274
rect 8128 13252 8260 13258
rect 8128 13246 8208 13252
rect 8208 13194 8260 13200
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 7760 12986 7788 13126
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 8312 12850 8340 13126
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 7852 12442 7880 12786
rect 8036 12646 8064 12786
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 8116 12640 8168 12646
rect 8116 12582 8168 12588
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7656 11824 7708 11830
rect 7656 11766 7708 11772
rect 7668 11150 7696 11766
rect 7760 11694 7788 12174
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7656 10736 7708 10742
rect 7656 10678 7708 10684
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7392 10062 7420 10406
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7380 10056 7432 10062
rect 7484 10044 7512 10610
rect 7668 10062 7696 10678
rect 7564 10056 7616 10062
rect 7484 10016 7564 10044
rect 7380 9998 7432 10004
rect 7564 9998 7616 10004
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7760 9926 7788 11630
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 7944 10674 7972 11018
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 7944 10062 7972 10610
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7116 8974 7144 9318
rect 7300 8974 7328 9862
rect 7668 9586 7696 9862
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7104 8968 7156 8974
rect 7010 8936 7066 8945
rect 7104 8910 7156 8916
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7010 8871 7012 8880
rect 7064 8871 7066 8880
rect 7012 8842 7064 8848
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 7116 8498 7144 8774
rect 7484 8498 7512 8774
rect 7576 8634 7604 9318
rect 8036 9110 8064 12582
rect 8128 12170 8156 12582
rect 8116 12164 8168 12170
rect 8116 12106 8168 12112
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 8220 10674 8248 11018
rect 8312 11014 8340 11698
rect 8404 11150 8432 16390
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8496 14414 8524 15098
rect 8576 15020 8628 15026
rect 8576 14962 8628 14968
rect 8588 14414 8616 14962
rect 8758 14512 8814 14521
rect 8758 14447 8760 14456
rect 8812 14447 8814 14456
rect 8760 14418 8812 14424
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8680 14278 8708 14350
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8680 14006 8708 14214
rect 8668 14000 8720 14006
rect 8668 13942 8720 13948
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8588 12102 8616 12786
rect 8680 12714 8708 13126
rect 8668 12708 8720 12714
rect 8668 12650 8720 12656
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8772 11762 8800 13262
rect 8864 11830 8892 17478
rect 9416 17270 9444 17478
rect 9404 17264 9456 17270
rect 9404 17206 9456 17212
rect 8944 16448 8996 16454
rect 8944 16390 8996 16396
rect 8956 15162 8984 16390
rect 9416 16114 9444 17206
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9508 16250 9536 16594
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 8944 15156 8996 15162
rect 8944 15098 8996 15104
rect 9220 15088 9272 15094
rect 9140 15048 9220 15076
rect 9140 14550 9168 15048
rect 9220 15030 9272 15036
rect 9404 15020 9456 15026
rect 9404 14962 9456 14968
rect 9416 14618 9444 14962
rect 9496 14952 9548 14958
rect 9496 14894 9548 14900
rect 9508 14618 9536 14894
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9128 14544 9180 14550
rect 9508 14498 9536 14554
rect 9128 14486 9180 14492
rect 9416 14470 9536 14498
rect 9416 14278 9444 14470
rect 9496 14408 9548 14414
rect 9496 14350 9548 14356
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 9232 13530 9260 13670
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 8942 12744 8998 12753
rect 8942 12679 8944 12688
rect 8996 12679 8998 12688
rect 8944 12650 8996 12656
rect 9508 12102 9536 14350
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9600 11830 9628 16934
rect 9876 15706 9904 18566
rect 9968 17678 9996 18566
rect 10060 18426 10088 18566
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 9956 17672 10008 17678
rect 9956 17614 10008 17620
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 10060 15502 10088 17478
rect 10520 16697 10548 21082
rect 10600 20868 10652 20874
rect 10600 20810 10652 20816
rect 10612 20602 10640 20810
rect 10600 20596 10652 20602
rect 10600 20538 10652 20544
rect 10704 19990 10732 22918
rect 10692 19984 10744 19990
rect 10692 19926 10744 19932
rect 10692 19848 10744 19854
rect 10796 19836 10824 24618
rect 10888 24274 10916 24754
rect 10876 24268 10928 24274
rect 10876 24210 10928 24216
rect 10888 24070 10916 24210
rect 10876 24064 10928 24070
rect 10876 24006 10928 24012
rect 10876 23180 10928 23186
rect 10876 23122 10928 23128
rect 10888 22642 10916 23122
rect 10980 23066 11008 24822
rect 11072 23798 11100 25230
rect 11244 25152 11296 25158
rect 11244 25094 11296 25100
rect 11256 24206 11284 25094
rect 11348 24274 11376 25434
rect 11336 24268 11388 24274
rect 11336 24210 11388 24216
rect 11244 24200 11296 24206
rect 11244 24142 11296 24148
rect 11060 23792 11112 23798
rect 11060 23734 11112 23740
rect 11336 23656 11388 23662
rect 11336 23598 11388 23604
rect 11152 23520 11204 23526
rect 11152 23462 11204 23468
rect 11244 23520 11296 23526
rect 11244 23462 11296 23468
rect 10980 23038 11100 23066
rect 10968 22976 11020 22982
rect 10968 22918 11020 22924
rect 10876 22636 10928 22642
rect 10876 22578 10928 22584
rect 10876 22024 10928 22030
rect 10876 21966 10928 21972
rect 10888 21146 10916 21966
rect 10876 21140 10928 21146
rect 10876 21082 10928 21088
rect 10876 19984 10928 19990
rect 10876 19926 10928 19932
rect 10744 19808 10824 19836
rect 10692 19790 10744 19796
rect 10600 19168 10652 19174
rect 10600 19110 10652 19116
rect 10612 18766 10640 19110
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 10704 18136 10732 19790
rect 10612 18108 10732 18136
rect 10506 16688 10562 16697
rect 10506 16623 10508 16632
rect 10560 16623 10562 16632
rect 10508 16594 10560 16600
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 10508 15428 10560 15434
rect 10508 15370 10560 15376
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 10416 15360 10468 15366
rect 10416 15302 10468 15308
rect 9864 15020 9916 15026
rect 9864 14962 9916 14968
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9692 12782 9720 14350
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 9784 13394 9812 13874
rect 9876 13802 9904 14962
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 9968 14414 9996 14554
rect 10060 14414 10088 15302
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10244 14958 10272 15098
rect 10232 14952 10284 14958
rect 10232 14894 10284 14900
rect 10324 14952 10376 14958
rect 10324 14894 10376 14900
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 10152 14618 10180 14758
rect 10336 14618 10364 14894
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 10428 14498 10456 15302
rect 10152 14482 10456 14498
rect 10140 14476 10456 14482
rect 10192 14470 10456 14476
rect 10140 14418 10192 14424
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 10048 14408 10100 14414
rect 10048 14350 10100 14356
rect 10152 14074 10180 14418
rect 10428 14414 10456 14470
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 9864 13796 9916 13802
rect 9864 13738 9916 13744
rect 9876 13462 9904 13738
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9968 13326 9996 13942
rect 10428 13938 10456 14214
rect 10520 13938 10548 15370
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 10244 12850 10272 13670
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10520 11898 10548 12106
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 8852 11824 8904 11830
rect 8852 11766 8904 11772
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8864 11626 8892 11766
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 8852 11620 8904 11626
rect 8852 11562 8904 11568
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8680 11354 8708 11494
rect 9324 11354 9352 11698
rect 9588 11688 9640 11694
rect 9864 11688 9916 11694
rect 9588 11630 9640 11636
rect 9784 11648 9864 11676
rect 9600 11558 9628 11630
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9600 11218 9628 11494
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 8392 11144 8444 11150
rect 9312 11144 9364 11150
rect 8444 11104 8524 11132
rect 8392 11086 8444 11092
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8392 10736 8444 10742
rect 8392 10678 8444 10684
rect 8496 10690 8524 11104
rect 9312 11086 9364 11092
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 8760 10736 8812 10742
rect 8496 10684 8760 10690
rect 8496 10678 8812 10684
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8128 10130 8156 10406
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 7748 9104 7800 9110
rect 7748 9046 7800 9052
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7012 8424 7064 8430
rect 7010 8392 7012 8401
rect 7064 8392 7066 8401
rect 7010 8327 7066 8336
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 6748 7886 6776 8026
rect 7208 8022 7236 8434
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7196 8016 7248 8022
rect 7196 7958 7248 7964
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 7300 7546 7328 8366
rect 7576 7886 7604 8570
rect 7760 8498 7788 9046
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 8036 8922 8064 9046
rect 8116 9036 8168 9042
rect 8168 8996 8248 9024
rect 8116 8978 8168 8984
rect 8220 8945 8248 8996
rect 8206 8936 8262 8945
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7852 7886 7880 8910
rect 8036 8894 8156 8922
rect 7932 8424 7984 8430
rect 7930 8392 7932 8401
rect 7984 8392 7986 8401
rect 7930 8327 7986 8336
rect 8128 8294 8156 8894
rect 8206 8871 8262 8880
rect 8220 8498 8248 8871
rect 8312 8566 8340 9998
rect 8404 9450 8432 10678
rect 8496 10662 8800 10678
rect 8496 10470 8524 10662
rect 9324 10538 9352 11086
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9312 10532 9364 10538
rect 9312 10474 9364 10480
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8496 9722 8524 10406
rect 8772 10266 8800 10406
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8680 9722 8708 10202
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 9048 9926 9076 10066
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8496 9450 8524 9658
rect 9324 9654 9352 9862
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9416 9586 9444 11018
rect 9508 11014 9536 11086
rect 9784 11014 9812 11648
rect 9864 11630 9916 11636
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10060 11234 10088 11494
rect 9968 11206 10088 11234
rect 9968 11150 9996 11206
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9784 10606 9812 10950
rect 9864 10668 9916 10674
rect 9968 10656 9996 11086
rect 10060 10810 10088 11086
rect 10336 11082 10364 11630
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 9916 10628 9996 10656
rect 10140 10668 10192 10674
rect 9864 10610 9916 10616
rect 10140 10610 10192 10616
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9588 10192 9640 10198
rect 9588 10134 9640 10140
rect 9600 9994 9628 10134
rect 10152 10062 10180 10610
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10244 10062 10272 10406
rect 10324 10192 10376 10198
rect 10324 10134 10376 10140
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 9588 9988 9640 9994
rect 9588 9930 9640 9936
rect 10244 9654 10272 9998
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8484 9444 8536 9450
rect 8484 9386 8536 9392
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 8956 9042 8984 9318
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 8220 8090 8248 8434
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 7944 7954 7972 8026
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 8220 7410 8248 8026
rect 8312 7954 8340 8366
rect 8404 8294 8432 8774
rect 8956 8634 8984 8978
rect 9048 8974 9076 9318
rect 9140 9178 9168 9522
rect 10336 9178 10364 10134
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 9864 9172 9916 9178
rect 9864 9114 9916 9120
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8496 8498 8524 8570
rect 9048 8498 9076 8910
rect 9876 8566 9904 9114
rect 10428 8974 10456 10746
rect 10520 8974 10548 11834
rect 10612 8974 10640 18108
rect 10888 17746 10916 19926
rect 10876 17740 10928 17746
rect 10876 17682 10928 17688
rect 10874 17096 10930 17105
rect 10874 17031 10876 17040
rect 10928 17031 10930 17040
rect 10876 17002 10928 17008
rect 10980 16810 11008 22918
rect 11072 22030 11100 23038
rect 11164 22030 11192 23462
rect 11256 22166 11284 23462
rect 11348 23118 11376 23598
rect 11336 23112 11388 23118
rect 11336 23054 11388 23060
rect 11348 22710 11376 23054
rect 11440 22982 11468 30518
rect 11612 30320 11664 30326
rect 11612 30262 11664 30268
rect 11704 30320 11756 30326
rect 11704 30262 11756 30268
rect 11520 29572 11572 29578
rect 11520 29514 11572 29520
rect 11532 29481 11560 29514
rect 11518 29472 11574 29481
rect 11518 29407 11574 29416
rect 11624 28626 11652 30262
rect 11716 29617 11744 30262
rect 11888 30184 11940 30190
rect 11888 30126 11940 30132
rect 11796 29640 11848 29646
rect 11702 29608 11758 29617
rect 11796 29582 11848 29588
rect 11702 29543 11758 29552
rect 11716 29306 11744 29543
rect 11704 29300 11756 29306
rect 11704 29242 11756 29248
rect 11704 29164 11756 29170
rect 11704 29106 11756 29112
rect 11716 28966 11744 29106
rect 11704 28960 11756 28966
rect 11704 28902 11756 28908
rect 11808 28762 11836 29582
rect 11900 28762 11928 30126
rect 11980 30116 12032 30122
rect 11980 30058 12032 30064
rect 11992 29238 12020 30058
rect 12176 29594 12204 30602
rect 12440 30252 12492 30258
rect 12440 30194 12492 30200
rect 12348 30048 12400 30054
rect 12348 29990 12400 29996
rect 12256 29844 12308 29850
rect 12256 29786 12308 29792
rect 12084 29566 12204 29594
rect 11980 29232 12032 29238
rect 11980 29174 12032 29180
rect 11796 28756 11848 28762
rect 11796 28698 11848 28704
rect 11888 28756 11940 28762
rect 11888 28698 11940 28704
rect 11612 28620 11664 28626
rect 11612 28562 11664 28568
rect 11704 28552 11756 28558
rect 11756 28500 11836 28506
rect 11704 28494 11836 28500
rect 11716 28478 11836 28494
rect 11808 28422 11836 28478
rect 11704 28416 11756 28422
rect 11704 28358 11756 28364
rect 11796 28416 11848 28422
rect 11796 28358 11848 28364
rect 11716 28082 11744 28358
rect 11808 28082 11836 28358
rect 11704 28076 11756 28082
rect 11704 28018 11756 28024
rect 11796 28076 11848 28082
rect 11796 28018 11848 28024
rect 11808 27674 11836 28018
rect 11520 27668 11572 27674
rect 11520 27610 11572 27616
rect 11796 27668 11848 27674
rect 11796 27610 11848 27616
rect 11532 26994 11560 27610
rect 11900 27554 11928 28698
rect 12084 28422 12112 29566
rect 12164 29504 12216 29510
rect 12164 29446 12216 29452
rect 12176 29170 12204 29446
rect 12268 29322 12296 29786
rect 12360 29646 12388 29990
rect 12348 29640 12400 29646
rect 12348 29582 12400 29588
rect 12348 29504 12400 29510
rect 12348 29446 12400 29452
rect 12360 29322 12388 29446
rect 12268 29294 12388 29322
rect 12452 29306 12480 30194
rect 12636 30138 12664 32302
rect 12716 31816 12768 31822
rect 12716 31758 12768 31764
rect 12728 31482 12756 31758
rect 12716 31476 12768 31482
rect 12716 31418 12768 31424
rect 12544 30122 12664 30138
rect 12532 30116 12664 30122
rect 12584 30110 12664 30116
rect 12532 30058 12584 30064
rect 12532 29640 12584 29646
rect 12532 29582 12584 29588
rect 12440 29300 12492 29306
rect 12164 29164 12216 29170
rect 12164 29106 12216 29112
rect 12268 28558 12296 29294
rect 12440 29242 12492 29248
rect 12348 29232 12400 29238
rect 12348 29174 12400 29180
rect 12256 28552 12308 28558
rect 12256 28494 12308 28500
rect 12072 28416 12124 28422
rect 12072 28358 12124 28364
rect 11624 27526 11928 27554
rect 12256 27532 12308 27538
rect 11520 26988 11572 26994
rect 11520 26930 11572 26936
rect 11520 23724 11572 23730
rect 11520 23666 11572 23672
rect 11532 23322 11560 23666
rect 11520 23316 11572 23322
rect 11520 23258 11572 23264
rect 11532 23186 11560 23258
rect 11520 23180 11572 23186
rect 11520 23122 11572 23128
rect 11428 22976 11480 22982
rect 11428 22918 11480 22924
rect 11520 22976 11572 22982
rect 11624 22964 11652 27526
rect 12256 27474 12308 27480
rect 11980 26852 12032 26858
rect 11980 26794 12032 26800
rect 11888 26784 11940 26790
rect 11888 26726 11940 26732
rect 11704 26512 11756 26518
rect 11704 26454 11756 26460
rect 11716 25906 11744 26454
rect 11900 26042 11928 26726
rect 11992 26314 12020 26794
rect 12072 26784 12124 26790
rect 12072 26726 12124 26732
rect 12268 26738 12296 27474
rect 12360 27044 12388 29174
rect 12440 29164 12492 29170
rect 12440 29106 12492 29112
rect 12452 28490 12480 29106
rect 12544 29102 12572 29582
rect 12624 29232 12676 29238
rect 12624 29174 12676 29180
rect 12532 29096 12584 29102
rect 12532 29038 12584 29044
rect 12440 28484 12492 28490
rect 12440 28426 12492 28432
rect 12636 28082 12664 29174
rect 12624 28076 12676 28082
rect 12624 28018 12676 28024
rect 12716 28076 12768 28082
rect 12716 28018 12768 28024
rect 12532 27872 12584 27878
rect 12530 27840 12532 27849
rect 12584 27840 12586 27849
rect 12530 27775 12586 27784
rect 12440 27056 12492 27062
rect 12360 27016 12440 27044
rect 12440 26998 12492 27004
rect 12084 26586 12112 26726
rect 12268 26710 12388 26738
rect 12072 26580 12124 26586
rect 12072 26522 12124 26528
rect 12256 26580 12308 26586
rect 12256 26522 12308 26528
rect 11980 26308 12032 26314
rect 11980 26250 12032 26256
rect 11888 26036 11940 26042
rect 11888 25978 11940 25984
rect 11900 25906 11928 25978
rect 11992 25906 12020 26250
rect 11704 25900 11756 25906
rect 11704 25842 11756 25848
rect 11888 25900 11940 25906
rect 11888 25842 11940 25848
rect 11980 25900 12032 25906
rect 11980 25842 12032 25848
rect 11716 23662 11744 25842
rect 11796 24812 11848 24818
rect 11796 24754 11848 24760
rect 11808 24585 11836 24754
rect 11794 24576 11850 24585
rect 11794 24511 11850 24520
rect 11900 23730 11928 25842
rect 11980 25288 12032 25294
rect 11980 25230 12032 25236
rect 11992 24954 12020 25230
rect 11980 24948 12032 24954
rect 11980 24890 12032 24896
rect 11978 24848 12034 24857
rect 11978 24783 11980 24792
rect 12032 24783 12034 24792
rect 11980 24754 12032 24760
rect 11888 23724 11940 23730
rect 11888 23666 11940 23672
rect 11704 23656 11756 23662
rect 11704 23598 11756 23604
rect 11980 23248 12032 23254
rect 11980 23190 12032 23196
rect 11992 23089 12020 23190
rect 12084 23186 12112 26522
rect 12164 26376 12216 26382
rect 12164 26318 12216 26324
rect 12176 25702 12204 26318
rect 12268 26042 12296 26522
rect 12256 26036 12308 26042
rect 12256 25978 12308 25984
rect 12164 25696 12216 25702
rect 12164 25638 12216 25644
rect 12176 23322 12204 25638
rect 12256 24948 12308 24954
rect 12256 24890 12308 24896
rect 12268 24138 12296 24890
rect 12256 24132 12308 24138
rect 12256 24074 12308 24080
rect 12164 23316 12216 23322
rect 12164 23258 12216 23264
rect 12072 23180 12124 23186
rect 12072 23122 12124 23128
rect 11978 23080 12034 23089
rect 11704 23044 11756 23050
rect 11978 23015 12034 23024
rect 12164 23044 12216 23050
rect 11704 22986 11756 22992
rect 12164 22986 12216 22992
rect 11572 22936 11652 22964
rect 11520 22918 11572 22924
rect 11336 22704 11388 22710
rect 11336 22646 11388 22652
rect 11244 22160 11296 22166
rect 11244 22102 11296 22108
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 11152 22024 11204 22030
rect 11152 21966 11204 21972
rect 11164 21622 11192 21966
rect 11152 21616 11204 21622
rect 11152 21558 11204 21564
rect 11256 21010 11284 22102
rect 11440 21418 11468 22918
rect 11532 22166 11560 22918
rect 11612 22568 11664 22574
rect 11612 22510 11664 22516
rect 11520 22160 11572 22166
rect 11520 22102 11572 22108
rect 11624 22030 11652 22510
rect 11612 22024 11664 22030
rect 11612 21966 11664 21972
rect 11428 21412 11480 21418
rect 11428 21354 11480 21360
rect 11244 21004 11296 21010
rect 11244 20946 11296 20952
rect 11072 18834 11192 18850
rect 11256 18834 11284 20946
rect 11520 20868 11572 20874
rect 11520 20810 11572 20816
rect 11532 20602 11560 20810
rect 11520 20596 11572 20602
rect 11520 20538 11572 20544
rect 11072 18828 11204 18834
rect 11072 18822 11152 18828
rect 11072 18222 11100 18822
rect 11152 18770 11204 18776
rect 11244 18828 11296 18834
rect 11244 18770 11296 18776
rect 11152 18692 11204 18698
rect 11152 18634 11204 18640
rect 11164 18426 11192 18634
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 11060 17264 11112 17270
rect 11060 17206 11112 17212
rect 10888 16782 11008 16810
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10704 16182 10732 16390
rect 10692 16176 10744 16182
rect 10692 16118 10744 16124
rect 10888 15978 10916 16782
rect 11072 16522 11100 17206
rect 11060 16516 11112 16522
rect 11060 16458 11112 16464
rect 11072 16250 11100 16458
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 10876 15972 10928 15978
rect 10876 15914 10928 15920
rect 10888 15881 10916 15914
rect 10874 15872 10930 15881
rect 10874 15807 10930 15816
rect 11072 15502 11100 16186
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 10796 14618 10824 14962
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10980 12850 11008 13806
rect 11072 13802 11100 13874
rect 11060 13796 11112 13802
rect 11060 13738 11112 13744
rect 11072 13462 11100 13738
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 11060 12776 11112 12782
rect 10980 12724 11060 12730
rect 10980 12718 11112 12724
rect 10980 12702 11100 12718
rect 10980 11830 11008 12702
rect 10968 11824 11020 11830
rect 10968 11766 11020 11772
rect 10980 11694 11008 11766
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 11164 11150 11192 17478
rect 11244 17332 11296 17338
rect 11244 17274 11296 17280
rect 11256 16590 11284 17274
rect 11716 16697 11744 22986
rect 11978 22672 12034 22681
rect 11978 22607 11980 22616
rect 12032 22607 12034 22616
rect 11980 22578 12032 22584
rect 11992 21690 12020 22578
rect 12176 22574 12204 22986
rect 12360 22778 12388 26710
rect 12452 26382 12480 26998
rect 12532 26920 12584 26926
rect 12532 26862 12584 26868
rect 12440 26376 12492 26382
rect 12440 26318 12492 26324
rect 12440 25900 12492 25906
rect 12440 25842 12492 25848
rect 12452 24614 12480 25842
rect 12544 25838 12572 26862
rect 12636 26586 12664 28018
rect 12728 27674 12756 28018
rect 12716 27668 12768 27674
rect 12716 27610 12768 27616
rect 12624 26580 12676 26586
rect 12624 26522 12676 26528
rect 12624 26308 12676 26314
rect 12624 26250 12676 26256
rect 12636 26217 12664 26250
rect 12622 26208 12678 26217
rect 12622 26143 12678 26152
rect 12532 25832 12584 25838
rect 12532 25774 12584 25780
rect 12820 24970 12848 35634
rect 12912 35086 12940 36586
rect 13096 36310 13124 36722
rect 13084 36304 13136 36310
rect 13084 36246 13136 36252
rect 13084 35148 13136 35154
rect 13084 35090 13136 35096
rect 12900 35080 12952 35086
rect 12898 35048 12900 35057
rect 12952 35048 12954 35057
rect 12898 34983 12954 34992
rect 13096 33998 13124 35090
rect 13084 33992 13136 33998
rect 13084 33934 13136 33940
rect 13096 33522 13124 33934
rect 13084 33516 13136 33522
rect 13084 33458 13136 33464
rect 13084 32428 13136 32434
rect 13084 32370 13136 32376
rect 12992 32292 13044 32298
rect 12992 32234 13044 32240
rect 13004 31686 13032 32234
rect 12992 31680 13044 31686
rect 12992 31622 13044 31628
rect 12900 31340 12952 31346
rect 12900 31282 12952 31288
rect 12992 31340 13044 31346
rect 12992 31282 13044 31288
rect 12912 30598 12940 31282
rect 12900 30592 12952 30598
rect 12900 30534 12952 30540
rect 12900 30116 12952 30122
rect 12900 30058 12952 30064
rect 12912 29646 12940 30058
rect 12900 29640 12952 29646
rect 12900 29582 12952 29588
rect 12544 24942 12848 24970
rect 12544 24614 12572 24942
rect 12440 24608 12492 24614
rect 12440 24550 12492 24556
rect 12532 24608 12584 24614
rect 12532 24550 12584 24556
rect 12624 24608 12676 24614
rect 12624 24550 12676 24556
rect 12440 23656 12492 23662
rect 12440 23598 12492 23604
rect 12452 23322 12480 23598
rect 12440 23316 12492 23322
rect 12440 23258 12492 23264
rect 12544 23202 12572 24550
rect 12636 24206 12664 24550
rect 12624 24200 12676 24206
rect 12624 24142 12676 24148
rect 12452 23174 12572 23202
rect 12348 22772 12400 22778
rect 12348 22714 12400 22720
rect 12164 22568 12216 22574
rect 12164 22510 12216 22516
rect 12164 22432 12216 22438
rect 12164 22374 12216 22380
rect 12072 22228 12124 22234
rect 12072 22170 12124 22176
rect 12084 22030 12112 22170
rect 12072 22024 12124 22030
rect 12072 21966 12124 21972
rect 11980 21684 12032 21690
rect 11980 21626 12032 21632
rect 11888 17128 11940 17134
rect 11888 17070 11940 17076
rect 11702 16688 11758 16697
rect 11702 16623 11704 16632
rect 11756 16623 11758 16632
rect 11704 16594 11756 16600
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 11256 16182 11284 16526
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11716 16250 11744 16390
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11244 16176 11296 16182
rect 11244 16118 11296 16124
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11336 13252 11388 13258
rect 11336 13194 11388 13200
rect 11348 12714 11376 13194
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11440 11150 11468 15846
rect 11808 15502 11836 15846
rect 11900 15502 11928 17070
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 11992 16114 12020 16934
rect 12176 16726 12204 22374
rect 12256 20868 12308 20874
rect 12256 20810 12308 20816
rect 12268 18766 12296 20810
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 12452 18272 12480 23174
rect 12624 22772 12676 22778
rect 12624 22714 12676 22720
rect 12636 22166 12664 22714
rect 12624 22160 12676 22166
rect 12624 22102 12676 22108
rect 12806 22128 12862 22137
rect 12912 22098 12940 29582
rect 13004 27606 13032 31282
rect 13096 30734 13124 32370
rect 13084 30728 13136 30734
rect 13084 30670 13136 30676
rect 13096 30394 13124 30670
rect 13084 30388 13136 30394
rect 13084 30330 13136 30336
rect 13096 29714 13124 30330
rect 13188 30190 13216 36790
rect 13544 36780 13596 36786
rect 13544 36722 13596 36728
rect 13556 36106 13584 36722
rect 13544 36100 13596 36106
rect 13544 36042 13596 36048
rect 13360 36032 13412 36038
rect 13360 35974 13412 35980
rect 13728 36032 13780 36038
rect 13728 35974 13780 35980
rect 13268 30592 13320 30598
rect 13268 30534 13320 30540
rect 13280 30326 13308 30534
rect 13268 30320 13320 30326
rect 13268 30262 13320 30268
rect 13176 30184 13228 30190
rect 13176 30126 13228 30132
rect 13084 29708 13136 29714
rect 13084 29650 13136 29656
rect 13372 29617 13400 35974
rect 13740 35630 13768 35974
rect 13832 35766 13860 37130
rect 14004 37120 14056 37126
rect 14004 37062 14056 37068
rect 14016 36786 14044 37062
rect 14004 36780 14056 36786
rect 14004 36722 14056 36728
rect 14200 36718 14228 37198
rect 14292 36854 14320 39850
rect 14476 39438 14504 39918
rect 14464 39432 14516 39438
rect 14464 39374 14516 39380
rect 14648 39296 14700 39302
rect 14648 39238 14700 39244
rect 14660 39098 14688 39238
rect 15028 39098 15056 39986
rect 15200 39840 15252 39846
rect 15200 39782 15252 39788
rect 15212 39438 15240 39782
rect 15292 39636 15344 39642
rect 15292 39578 15344 39584
rect 15200 39432 15252 39438
rect 15200 39374 15252 39380
rect 15304 39250 15332 39578
rect 15488 39370 15516 40122
rect 15568 40044 15620 40050
rect 15568 39986 15620 39992
rect 15580 39574 15608 39986
rect 15764 39914 15792 40462
rect 15936 40384 15988 40390
rect 15936 40326 15988 40332
rect 15752 39908 15804 39914
rect 15752 39850 15804 39856
rect 15568 39568 15620 39574
rect 15568 39510 15620 39516
rect 15476 39364 15528 39370
rect 15476 39306 15528 39312
rect 15212 39222 15332 39250
rect 14648 39092 14700 39098
rect 14648 39034 14700 39040
rect 15016 39092 15068 39098
rect 15016 39034 15068 39040
rect 15212 38554 15240 39222
rect 15200 38548 15252 38554
rect 15200 38490 15252 38496
rect 14832 38208 14884 38214
rect 14832 38150 14884 38156
rect 14844 37874 14872 38150
rect 15016 37936 15068 37942
rect 15016 37878 15068 37884
rect 14832 37868 14884 37874
rect 14832 37810 14884 37816
rect 14844 37398 14872 37810
rect 14832 37392 14884 37398
rect 14832 37334 14884 37340
rect 14648 37256 14700 37262
rect 14648 37198 14700 37204
rect 14740 37256 14792 37262
rect 14740 37198 14792 37204
rect 14280 36848 14332 36854
rect 14280 36790 14332 36796
rect 14188 36712 14240 36718
rect 14188 36654 14240 36660
rect 14200 36281 14228 36654
rect 14556 36576 14608 36582
rect 14556 36518 14608 36524
rect 14186 36272 14242 36281
rect 14568 36242 14596 36518
rect 14186 36207 14242 36216
rect 14556 36236 14608 36242
rect 14556 36178 14608 36184
rect 13820 35760 13872 35766
rect 13820 35702 13872 35708
rect 13728 35624 13780 35630
rect 13728 35566 13780 35572
rect 13544 35488 13596 35494
rect 13544 35430 13596 35436
rect 13452 35148 13504 35154
rect 13452 35090 13504 35096
rect 13464 29782 13492 35090
rect 13452 29776 13504 29782
rect 13452 29718 13504 29724
rect 13082 29608 13138 29617
rect 13082 29543 13138 29552
rect 13358 29608 13414 29617
rect 13358 29543 13414 29552
rect 12992 27600 13044 27606
rect 12992 27542 13044 27548
rect 13096 25906 13124 29543
rect 13176 29504 13228 29510
rect 13556 29481 13584 35430
rect 13832 34746 13860 35702
rect 14660 35476 14688 37198
rect 14752 36378 14780 37198
rect 14740 36372 14792 36378
rect 14740 36314 14792 36320
rect 14844 36242 14872 37334
rect 15028 36582 15056 37878
rect 15212 37806 15240 38490
rect 15384 37868 15436 37874
rect 15384 37810 15436 37816
rect 15200 37800 15252 37806
rect 15200 37742 15252 37748
rect 15212 37210 15240 37742
rect 15292 37664 15344 37670
rect 15292 37606 15344 37612
rect 15304 37330 15332 37606
rect 15396 37466 15424 37810
rect 15384 37460 15436 37466
rect 15384 37402 15436 37408
rect 15292 37324 15344 37330
rect 15292 37266 15344 37272
rect 15212 37182 15424 37210
rect 15200 36916 15252 36922
rect 15200 36858 15252 36864
rect 15212 36786 15240 36858
rect 15200 36780 15252 36786
rect 15200 36722 15252 36728
rect 15292 36780 15344 36786
rect 15292 36722 15344 36728
rect 15016 36576 15068 36582
rect 15016 36518 15068 36524
rect 14832 36236 14884 36242
rect 14832 36178 14884 36184
rect 15028 35766 15056 36518
rect 15212 36394 15240 36722
rect 15120 36366 15240 36394
rect 15016 35760 15068 35766
rect 15016 35702 15068 35708
rect 14740 35488 14792 35494
rect 14660 35448 14740 35476
rect 14740 35430 14792 35436
rect 13820 34740 13872 34746
rect 13820 34682 13872 34688
rect 13832 34066 13860 34682
rect 15028 34678 15056 35702
rect 15120 35698 15148 36366
rect 15304 36310 15332 36722
rect 15292 36304 15344 36310
rect 15292 36246 15344 36252
rect 15200 36236 15252 36242
rect 15200 36178 15252 36184
rect 15108 35692 15160 35698
rect 15108 35634 15160 35640
rect 15016 34672 15068 34678
rect 15016 34614 15068 34620
rect 14280 34536 14332 34542
rect 14280 34478 14332 34484
rect 13820 34060 13872 34066
rect 13820 34002 13872 34008
rect 14292 33658 14320 34478
rect 14740 34400 14792 34406
rect 14740 34342 14792 34348
rect 14752 34066 14780 34342
rect 14740 34060 14792 34066
rect 14740 34002 14792 34008
rect 15028 33930 15056 34614
rect 15016 33924 15068 33930
rect 15016 33866 15068 33872
rect 14280 33652 14332 33658
rect 14280 33594 14332 33600
rect 14740 33652 14792 33658
rect 14740 33594 14792 33600
rect 14752 33454 14780 33594
rect 14740 33448 14792 33454
rect 14740 33390 14792 33396
rect 13912 32428 13964 32434
rect 13912 32370 13964 32376
rect 14188 32428 14240 32434
rect 14188 32370 14240 32376
rect 14648 32428 14700 32434
rect 14648 32370 14700 32376
rect 13820 32360 13872 32366
rect 13820 32302 13872 32308
rect 13728 31816 13780 31822
rect 13728 31758 13780 31764
rect 13636 31680 13688 31686
rect 13636 31622 13688 31628
rect 13648 31346 13676 31622
rect 13740 31346 13768 31758
rect 13832 31482 13860 32302
rect 13924 31822 13952 32370
rect 13912 31816 13964 31822
rect 13912 31758 13964 31764
rect 14200 31482 14228 32370
rect 14556 32224 14608 32230
rect 14556 32166 14608 32172
rect 14568 32026 14596 32166
rect 14556 32020 14608 32026
rect 14556 31962 14608 31968
rect 13820 31476 13872 31482
rect 13820 31418 13872 31424
rect 14188 31476 14240 31482
rect 14188 31418 14240 31424
rect 13636 31340 13688 31346
rect 13636 31282 13688 31288
rect 13728 31340 13780 31346
rect 13728 31282 13780 31288
rect 13912 31340 13964 31346
rect 13912 31282 13964 31288
rect 14188 31340 14240 31346
rect 14188 31282 14240 31288
rect 14464 31340 14516 31346
rect 14464 31282 14516 31288
rect 13176 29446 13228 29452
rect 13542 29472 13598 29481
rect 13084 25900 13136 25906
rect 13084 25842 13136 25848
rect 13188 23186 13216 29446
rect 13542 29407 13598 29416
rect 13360 28552 13412 28558
rect 13360 28494 13412 28500
rect 13372 28082 13400 28494
rect 13360 28076 13412 28082
rect 13360 28018 13412 28024
rect 13544 28076 13596 28082
rect 13544 28018 13596 28024
rect 13556 27606 13584 28018
rect 13544 27600 13596 27606
rect 13372 27560 13544 27588
rect 13268 27464 13320 27470
rect 13268 27406 13320 27412
rect 13280 26858 13308 27406
rect 13372 26994 13400 27560
rect 13544 27542 13596 27548
rect 13452 27464 13504 27470
rect 13648 27418 13676 31282
rect 13924 31142 13952 31282
rect 13912 31136 13964 31142
rect 13912 31078 13964 31084
rect 14200 30734 14228 31282
rect 14188 30728 14240 30734
rect 14108 30688 14188 30716
rect 14108 29646 14136 30688
rect 14188 30670 14240 30676
rect 14280 30388 14332 30394
rect 14280 30330 14332 30336
rect 14188 30252 14240 30258
rect 14188 30194 14240 30200
rect 14096 29640 14148 29646
rect 14096 29582 14148 29588
rect 14200 29578 14228 30194
rect 14292 30054 14320 30330
rect 14372 30252 14424 30258
rect 14372 30194 14424 30200
rect 14280 30048 14332 30054
rect 14280 29990 14332 29996
rect 14384 29646 14412 30194
rect 14372 29640 14424 29646
rect 14372 29582 14424 29588
rect 14188 29572 14240 29578
rect 14188 29514 14240 29520
rect 13820 29504 13872 29510
rect 13820 29446 13872 29452
rect 13832 29034 13860 29446
rect 13820 29028 13872 29034
rect 13820 28970 13872 28976
rect 13912 28688 13964 28694
rect 13912 28630 13964 28636
rect 13924 28150 13952 28630
rect 14096 28416 14148 28422
rect 14096 28358 14148 28364
rect 13912 28144 13964 28150
rect 13912 28086 13964 28092
rect 13820 28076 13872 28082
rect 13820 28018 13872 28024
rect 13832 27946 13860 28018
rect 13820 27940 13872 27946
rect 13820 27882 13872 27888
rect 13912 27940 13964 27946
rect 13912 27882 13964 27888
rect 13832 27674 13860 27882
rect 13820 27668 13872 27674
rect 13820 27610 13872 27616
rect 13452 27406 13504 27412
rect 13360 26988 13412 26994
rect 13360 26930 13412 26936
rect 13268 26852 13320 26858
rect 13268 26794 13320 26800
rect 13360 25900 13412 25906
rect 13464 25888 13492 27406
rect 13412 25860 13492 25888
rect 13556 27390 13676 27418
rect 13726 27432 13782 27441
rect 13360 25842 13412 25848
rect 13372 25498 13400 25842
rect 13360 25492 13412 25498
rect 13360 25434 13412 25440
rect 13556 24290 13584 27390
rect 13726 27367 13782 27376
rect 13740 27130 13768 27367
rect 13728 27124 13780 27130
rect 13728 27066 13780 27072
rect 13634 25936 13690 25945
rect 13634 25871 13636 25880
rect 13688 25871 13690 25880
rect 13636 25842 13688 25848
rect 13648 24410 13676 25842
rect 13740 25770 13768 27066
rect 13820 26988 13872 26994
rect 13820 26930 13872 26936
rect 13832 25906 13860 26930
rect 13924 26926 13952 27882
rect 14004 27872 14056 27878
rect 14004 27814 14056 27820
rect 13912 26920 13964 26926
rect 13912 26862 13964 26868
rect 14016 26058 14044 27814
rect 14108 27402 14136 28358
rect 14096 27396 14148 27402
rect 14096 27338 14148 27344
rect 14200 26790 14228 29514
rect 14384 29306 14412 29582
rect 14372 29300 14424 29306
rect 14372 29242 14424 29248
rect 14372 28756 14424 28762
rect 14372 28698 14424 28704
rect 14280 28552 14332 28558
rect 14280 28494 14332 28500
rect 14292 28082 14320 28494
rect 14280 28076 14332 28082
rect 14280 28018 14332 28024
rect 14384 28014 14412 28698
rect 14372 28008 14424 28014
rect 14372 27950 14424 27956
rect 14280 27872 14332 27878
rect 14372 27872 14424 27878
rect 14280 27814 14332 27820
rect 14370 27840 14372 27849
rect 14424 27840 14426 27849
rect 14188 26784 14240 26790
rect 14188 26726 14240 26732
rect 14096 26512 14148 26518
rect 14094 26480 14096 26489
rect 14148 26480 14150 26489
rect 14094 26415 14150 26424
rect 14016 26030 14136 26058
rect 14108 25906 14136 26030
rect 14200 25945 14228 26726
rect 14292 26586 14320 27814
rect 14370 27775 14426 27784
rect 14372 27328 14424 27334
rect 14372 27270 14424 27276
rect 14280 26580 14332 26586
rect 14280 26522 14332 26528
rect 14384 26450 14412 27270
rect 14372 26444 14424 26450
rect 14372 26386 14424 26392
rect 14280 26240 14332 26246
rect 14280 26182 14332 26188
rect 14186 25936 14242 25945
rect 13820 25900 13872 25906
rect 13820 25842 13872 25848
rect 13912 25900 13964 25906
rect 13912 25842 13964 25848
rect 14004 25900 14056 25906
rect 14004 25842 14056 25848
rect 14096 25900 14148 25906
rect 14186 25871 14242 25880
rect 14096 25842 14148 25848
rect 13728 25764 13780 25770
rect 13728 25706 13780 25712
rect 13728 25356 13780 25362
rect 13728 25298 13780 25304
rect 13636 24404 13688 24410
rect 13636 24346 13688 24352
rect 13556 24262 13676 24290
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 13556 23594 13584 23666
rect 13544 23588 13596 23594
rect 13544 23530 13596 23536
rect 13176 23180 13228 23186
rect 13176 23122 13228 23128
rect 13452 23180 13504 23186
rect 13452 23122 13504 23128
rect 12992 22568 13044 22574
rect 12992 22510 13044 22516
rect 12806 22063 12862 22072
rect 12900 22092 12952 22098
rect 12624 22024 12676 22030
rect 12624 21966 12676 21972
rect 12716 22024 12768 22030
rect 12716 21966 12768 21972
rect 12636 21622 12664 21966
rect 12728 21894 12756 21966
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12624 21616 12676 21622
rect 12624 21558 12676 21564
rect 12728 21418 12756 21830
rect 12716 21412 12768 21418
rect 12716 21354 12768 21360
rect 12820 20890 12848 22063
rect 12900 22034 12952 22040
rect 13004 22030 13032 22510
rect 12992 22024 13044 22030
rect 12992 21966 13044 21972
rect 13084 22024 13136 22030
rect 13084 21966 13136 21972
rect 13096 21690 13124 21966
rect 13084 21684 13136 21690
rect 13084 21626 13136 21632
rect 12900 21548 12952 21554
rect 12900 21490 12952 21496
rect 12992 21548 13044 21554
rect 12992 21490 13044 21496
rect 12912 21010 12940 21490
rect 13004 21350 13032 21490
rect 12992 21344 13044 21350
rect 12992 21286 13044 21292
rect 12900 21004 12952 21010
rect 12900 20946 12952 20952
rect 12728 20862 12848 20890
rect 12900 20868 12952 20874
rect 12728 19922 12756 20862
rect 12900 20810 12952 20816
rect 12808 20800 12860 20806
rect 12808 20742 12860 20748
rect 12820 20602 12848 20742
rect 12808 20596 12860 20602
rect 12808 20538 12860 20544
rect 12808 20460 12860 20466
rect 12808 20402 12860 20408
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 12544 19514 12572 19858
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12532 19508 12584 19514
rect 12532 19450 12584 19456
rect 12636 18970 12664 19790
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 12636 18766 12664 18906
rect 12624 18760 12676 18766
rect 12624 18702 12676 18708
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12636 18306 12664 18566
rect 12728 18426 12756 18566
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12820 18358 12848 20402
rect 12912 19854 12940 20810
rect 13004 20262 13032 21286
rect 13084 20528 13136 20534
rect 13188 20516 13216 23122
rect 13360 21956 13412 21962
rect 13360 21898 13412 21904
rect 13372 21554 13400 21898
rect 13464 21593 13492 23122
rect 13556 23050 13584 23530
rect 13544 23044 13596 23050
rect 13544 22986 13596 22992
rect 13648 22778 13676 24262
rect 13740 23730 13768 25298
rect 13924 24993 13952 25842
rect 14016 25786 14044 25842
rect 14292 25786 14320 26182
rect 14016 25758 14320 25786
rect 14476 25702 14504 31282
rect 14660 31278 14688 32370
rect 14740 32360 14792 32366
rect 14740 32302 14792 32308
rect 14752 31890 14780 32302
rect 15212 32298 15240 36178
rect 15292 34604 15344 34610
rect 15292 34546 15344 34552
rect 15304 33590 15332 34546
rect 15292 33584 15344 33590
rect 15292 33526 15344 33532
rect 15304 33114 15332 33526
rect 15292 33108 15344 33114
rect 15292 33050 15344 33056
rect 15396 32366 15424 37182
rect 15488 36038 15516 39306
rect 15580 37738 15608 39510
rect 15948 39506 15976 40326
rect 16408 40050 16436 40462
rect 16488 40384 16540 40390
rect 16488 40326 16540 40332
rect 16396 40044 16448 40050
rect 16396 39986 16448 39992
rect 16304 39976 16356 39982
rect 16224 39936 16304 39964
rect 15936 39500 15988 39506
rect 15936 39442 15988 39448
rect 16224 39438 16252 39936
rect 16304 39918 16356 39924
rect 16396 39840 16448 39846
rect 16396 39782 16448 39788
rect 16408 39642 16436 39782
rect 16396 39636 16448 39642
rect 16396 39578 16448 39584
rect 16500 39574 16528 40326
rect 16488 39568 16540 39574
rect 16488 39510 16540 39516
rect 16592 39438 16620 40462
rect 16856 39908 16908 39914
rect 16856 39850 16908 39856
rect 15844 39432 15896 39438
rect 16212 39432 16264 39438
rect 15896 39380 15976 39386
rect 15844 39374 15976 39380
rect 16212 39374 16264 39380
rect 16580 39432 16632 39438
rect 16580 39374 16632 39380
rect 15856 39358 15976 39374
rect 15948 39302 15976 39358
rect 15844 39296 15896 39302
rect 15844 39238 15896 39244
rect 15936 39296 15988 39302
rect 15936 39238 15988 39244
rect 15856 37874 15884 39238
rect 15844 37868 15896 37874
rect 15844 37810 15896 37816
rect 15568 37732 15620 37738
rect 15568 37674 15620 37680
rect 15580 37346 15608 37674
rect 15580 37330 15700 37346
rect 15580 37324 15712 37330
rect 15580 37318 15660 37324
rect 15580 36156 15608 37318
rect 15660 37266 15712 37272
rect 15660 37120 15712 37126
rect 15660 37062 15712 37068
rect 15672 36922 15700 37062
rect 15660 36916 15712 36922
rect 15660 36858 15712 36864
rect 15672 36310 15700 36858
rect 15660 36304 15712 36310
rect 15660 36246 15712 36252
rect 15842 36272 15898 36281
rect 15842 36207 15844 36216
rect 15896 36207 15898 36216
rect 15844 36178 15896 36184
rect 15580 36128 15792 36156
rect 15476 36032 15528 36038
rect 15476 35974 15528 35980
rect 15488 35630 15516 35974
rect 15476 35624 15528 35630
rect 15476 35566 15528 35572
rect 15660 35012 15712 35018
rect 15660 34954 15712 34960
rect 15672 34542 15700 34954
rect 15660 34536 15712 34542
rect 15660 34478 15712 34484
rect 15672 33658 15700 34478
rect 15660 33652 15712 33658
rect 15660 33594 15712 33600
rect 15566 33008 15622 33017
rect 15566 32943 15622 32952
rect 15580 32910 15608 32943
rect 15568 32904 15620 32910
rect 15568 32846 15620 32852
rect 15384 32360 15436 32366
rect 15384 32302 15436 32308
rect 15200 32292 15252 32298
rect 15200 32234 15252 32240
rect 14924 32020 14976 32026
rect 14924 31962 14976 31968
rect 14740 31884 14792 31890
rect 14740 31826 14792 31832
rect 14648 31272 14700 31278
rect 14648 31214 14700 31220
rect 14660 30258 14688 31214
rect 14830 30696 14886 30705
rect 14830 30631 14886 30640
rect 14648 30252 14700 30258
rect 14648 30194 14700 30200
rect 14660 30025 14688 30194
rect 14646 30016 14702 30025
rect 14646 29951 14702 29960
rect 14556 29844 14608 29850
rect 14556 29786 14608 29792
rect 14568 28098 14596 29786
rect 14740 29776 14792 29782
rect 14738 29744 14740 29753
rect 14792 29744 14794 29753
rect 14738 29679 14794 29688
rect 14648 29640 14700 29646
rect 14648 29582 14700 29588
rect 14660 29238 14688 29582
rect 14648 29232 14700 29238
rect 14648 29174 14700 29180
rect 14740 28620 14792 28626
rect 14740 28562 14792 28568
rect 14648 28552 14700 28558
rect 14648 28494 14700 28500
rect 14660 28218 14688 28494
rect 14648 28212 14700 28218
rect 14648 28154 14700 28160
rect 14568 28070 14688 28098
rect 14752 28082 14780 28562
rect 14844 28218 14872 30631
rect 14936 29646 14964 31962
rect 15292 31816 15344 31822
rect 15292 31758 15344 31764
rect 15476 31816 15528 31822
rect 15476 31758 15528 31764
rect 15304 31414 15332 31758
rect 15292 31408 15344 31414
rect 15292 31350 15344 31356
rect 15488 31346 15516 31758
rect 15476 31340 15528 31346
rect 15476 31282 15528 31288
rect 15016 31272 15068 31278
rect 15016 31214 15068 31220
rect 15384 31272 15436 31278
rect 15384 31214 15436 31220
rect 15028 30734 15056 31214
rect 15016 30728 15068 30734
rect 15016 30670 15068 30676
rect 15028 30258 15056 30670
rect 15292 30592 15344 30598
rect 15292 30534 15344 30540
rect 15016 30252 15068 30258
rect 15016 30194 15068 30200
rect 15108 30252 15160 30258
rect 15108 30194 15160 30200
rect 15028 29646 15056 30194
rect 14924 29640 14976 29646
rect 14924 29582 14976 29588
rect 15016 29640 15068 29646
rect 15016 29582 15068 29588
rect 15028 29102 15056 29582
rect 15016 29096 15068 29102
rect 15016 29038 15068 29044
rect 15016 28484 15068 28490
rect 15016 28426 15068 28432
rect 15028 28218 15056 28426
rect 14832 28212 14884 28218
rect 14832 28154 14884 28160
rect 15016 28212 15068 28218
rect 15016 28154 15068 28160
rect 14556 28008 14608 28014
rect 14556 27950 14608 27956
rect 14568 27674 14596 27950
rect 14556 27668 14608 27674
rect 14556 27610 14608 27616
rect 14568 27470 14596 27610
rect 14660 27470 14688 28070
rect 14740 28076 14792 28082
rect 14740 28018 14792 28024
rect 15028 28014 15056 28154
rect 15016 28008 15068 28014
rect 15016 27950 15068 27956
rect 14740 27940 14792 27946
rect 14740 27882 14792 27888
rect 14752 27674 14780 27882
rect 14740 27668 14792 27674
rect 14740 27610 14792 27616
rect 14752 27470 14780 27610
rect 15016 27532 15068 27538
rect 15016 27474 15068 27480
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 14648 27464 14700 27470
rect 14648 27406 14700 27412
rect 14740 27464 14792 27470
rect 14740 27406 14792 27412
rect 14832 27396 14884 27402
rect 14832 27338 14884 27344
rect 14844 27305 14872 27338
rect 14924 27328 14976 27334
rect 14830 27296 14886 27305
rect 14924 27270 14976 27276
rect 14830 27231 14886 27240
rect 14648 27124 14700 27130
rect 14648 27066 14700 27072
rect 14556 26988 14608 26994
rect 14556 26930 14608 26936
rect 14568 26586 14596 26930
rect 14660 26625 14688 27066
rect 14936 26994 14964 27270
rect 14924 26988 14976 26994
rect 14924 26930 14976 26936
rect 14740 26920 14792 26926
rect 14740 26862 14792 26868
rect 14832 26920 14884 26926
rect 14832 26862 14884 26868
rect 14646 26616 14702 26625
rect 14556 26580 14608 26586
rect 14646 26551 14702 26560
rect 14556 26522 14608 26528
rect 14554 26480 14610 26489
rect 14554 26415 14610 26424
rect 14568 26058 14596 26415
rect 14660 26382 14688 26551
rect 14752 26382 14780 26862
rect 14844 26586 14872 26862
rect 14924 26784 14976 26790
rect 14924 26726 14976 26732
rect 14832 26580 14884 26586
rect 14832 26522 14884 26528
rect 14648 26376 14700 26382
rect 14648 26318 14700 26324
rect 14740 26376 14792 26382
rect 14740 26318 14792 26324
rect 14832 26308 14884 26314
rect 14832 26250 14884 26256
rect 14568 26030 14688 26058
rect 14556 25900 14608 25906
rect 14556 25842 14608 25848
rect 14464 25696 14516 25702
rect 14186 25664 14242 25673
rect 14186 25599 14242 25608
rect 14384 25656 14464 25684
rect 13910 24984 13966 24993
rect 13910 24919 13966 24928
rect 14096 24812 14148 24818
rect 14096 24754 14148 24760
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 13728 23724 13780 23730
rect 13728 23666 13780 23672
rect 13924 23662 13952 24142
rect 13912 23656 13964 23662
rect 13912 23598 13964 23604
rect 13924 23526 13952 23598
rect 13912 23520 13964 23526
rect 13912 23462 13964 23468
rect 14004 23520 14056 23526
rect 14004 23462 14056 23468
rect 13820 23044 13872 23050
rect 13820 22986 13872 22992
rect 13832 22953 13860 22986
rect 13818 22944 13874 22953
rect 13818 22879 13874 22888
rect 13636 22772 13688 22778
rect 13636 22714 13688 22720
rect 13544 22024 13596 22030
rect 13544 21966 13596 21972
rect 13450 21584 13506 21593
rect 13360 21548 13412 21554
rect 13450 21519 13506 21528
rect 13360 21490 13412 21496
rect 13268 21480 13320 21486
rect 13268 21422 13320 21428
rect 13280 21146 13308 21422
rect 13268 21140 13320 21146
rect 13268 21082 13320 21088
rect 13136 20488 13216 20516
rect 13084 20470 13136 20476
rect 13280 20330 13308 21082
rect 13268 20324 13320 20330
rect 13268 20266 13320 20272
rect 12992 20256 13044 20262
rect 12992 20198 13044 20204
rect 13372 19990 13400 21490
rect 13360 19984 13412 19990
rect 13360 19926 13412 19932
rect 12900 19848 12952 19854
rect 12992 19848 13044 19854
rect 12900 19790 12952 19796
rect 12990 19816 12992 19825
rect 13044 19816 13046 19825
rect 12990 19751 13046 19760
rect 12808 18352 12860 18358
rect 12636 18278 12756 18306
rect 12860 18300 12940 18306
rect 12808 18294 12940 18300
rect 12820 18278 12940 18294
rect 12452 18244 12572 18272
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 12164 16720 12216 16726
rect 12084 16680 12164 16708
rect 11980 16108 12032 16114
rect 11980 16050 12032 16056
rect 12084 15994 12112 16680
rect 12164 16662 12216 16668
rect 12164 16516 12216 16522
rect 12164 16458 12216 16464
rect 11992 15966 12112 15994
rect 12176 15978 12204 16458
rect 12268 16250 12296 18158
rect 12440 18148 12492 18154
rect 12440 18090 12492 18096
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 12164 15972 12216 15978
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11612 14952 11664 14958
rect 11612 14894 11664 14900
rect 11624 14414 11652 14894
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11520 13932 11572 13938
rect 11520 13874 11572 13880
rect 11532 13394 11560 13874
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11532 13258 11560 13330
rect 11520 13252 11572 13258
rect 11520 13194 11572 13200
rect 11532 12918 11560 13194
rect 11520 12912 11572 12918
rect 11520 12854 11572 12860
rect 11624 12646 11652 14350
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10704 10062 10732 10950
rect 10888 10742 10916 11086
rect 10876 10736 10928 10742
rect 10876 10678 10928 10684
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 10704 9178 10732 9998
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8404 7954 8432 8230
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8312 7834 8340 7890
rect 8496 7834 8524 8298
rect 8312 7806 8524 7834
rect 8312 7410 8340 7806
rect 8680 7546 8708 8366
rect 9048 8022 9076 8434
rect 9140 8294 9168 8434
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9036 8016 9088 8022
rect 9036 7958 9088 7964
rect 9876 7954 9904 8502
rect 10336 7954 10364 8774
rect 10428 8498 10456 8774
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 9864 7948 9916 7954
rect 9864 7890 9916 7896
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 9508 7478 9536 7686
rect 10612 7528 10640 8910
rect 10704 7954 10732 9114
rect 10796 9110 10824 9454
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10784 9104 10836 9110
rect 10784 9046 10836 9052
rect 10888 8498 10916 9318
rect 10980 8786 11008 9590
rect 11072 9586 11100 9862
rect 11532 9722 11560 9998
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11716 9586 11744 14758
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11808 12850 11836 13670
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11900 12434 11928 14214
rect 11808 12406 11928 12434
rect 11808 10198 11836 12406
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11900 10674 11928 11630
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11900 10538 11928 10610
rect 11888 10532 11940 10538
rect 11888 10474 11940 10480
rect 11796 10192 11848 10198
rect 11796 10134 11848 10140
rect 11900 9994 11928 10474
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11072 8906 11100 9522
rect 11164 8974 11192 9522
rect 11440 9450 11468 9522
rect 11428 9444 11480 9450
rect 11428 9386 11480 9392
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11624 9058 11652 9318
rect 11348 9042 11652 9058
rect 11336 9036 11652 9042
rect 11388 9030 11652 9036
rect 11336 8978 11388 8984
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 11886 8936 11942 8945
rect 11060 8900 11112 8906
rect 11060 8842 11112 8848
rect 11152 8832 11204 8838
rect 10980 8780 11152 8786
rect 10980 8774 11204 8780
rect 10980 8758 11192 8774
rect 11440 8634 11468 8910
rect 11886 8871 11942 8880
rect 11900 8838 11928 8871
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 10980 8022 11008 8366
rect 11440 8022 11468 8570
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11610 8256 11666 8265
rect 11610 8191 11666 8200
rect 10968 8016 11020 8022
rect 10968 7958 11020 7964
rect 11428 8016 11480 8022
rect 11428 7958 11480 7964
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 11624 7818 11652 8191
rect 11900 8090 11928 8434
rect 11992 8090 12020 15966
rect 12164 15914 12216 15920
rect 12164 15428 12216 15434
rect 12164 15370 12216 15376
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 12084 14278 12112 14894
rect 12072 14272 12124 14278
rect 12072 14214 12124 14220
rect 12176 12434 12204 15370
rect 12360 13938 12388 16730
rect 12452 16436 12480 18090
rect 12544 17202 12572 18244
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12532 16448 12584 16454
rect 12452 16408 12532 16436
rect 12532 16390 12584 16396
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12544 15094 12572 15438
rect 12532 15088 12584 15094
rect 12532 15030 12584 15036
rect 12728 15026 12756 18278
rect 12808 18216 12860 18222
rect 12808 18158 12860 18164
rect 12820 17882 12848 18158
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 12820 16114 12848 17682
rect 12912 17610 12940 18278
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 13280 17678 13308 18158
rect 13464 17882 13492 21519
rect 13556 20058 13584 21966
rect 13728 21888 13780 21894
rect 13728 21830 13780 21836
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13556 19718 13584 19994
rect 13648 19961 13676 19994
rect 13634 19952 13690 19961
rect 13634 19887 13690 19896
rect 13544 19712 13596 19718
rect 13544 19654 13596 19660
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 13268 17672 13320 17678
rect 13188 17632 13268 17660
rect 12900 17604 12952 17610
rect 12900 17546 12952 17552
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12820 16017 12848 16050
rect 12806 16008 12862 16017
rect 12806 15943 12862 15952
rect 12912 15026 12940 17546
rect 12992 16652 13044 16658
rect 12992 16594 13044 16600
rect 13004 16182 13032 16594
rect 12992 16176 13044 16182
rect 12992 16118 13044 16124
rect 13188 15502 13216 17632
rect 13268 17614 13320 17620
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 13648 16114 13676 16934
rect 13740 16538 13768 21830
rect 13924 21622 13952 23462
rect 14016 23118 14044 23462
rect 14004 23112 14056 23118
rect 14004 23054 14056 23060
rect 14004 22976 14056 22982
rect 14004 22918 14056 22924
rect 14016 22642 14044 22918
rect 14004 22636 14056 22642
rect 14004 22578 14056 22584
rect 14108 22094 14136 24754
rect 14200 22710 14228 25599
rect 14384 23118 14412 25656
rect 14464 25638 14516 25644
rect 14568 25226 14596 25842
rect 14556 25220 14608 25226
rect 14556 25162 14608 25168
rect 14660 24818 14688 26030
rect 14464 24812 14516 24818
rect 14464 24754 14516 24760
rect 14648 24812 14700 24818
rect 14648 24754 14700 24760
rect 14740 24812 14792 24818
rect 14740 24754 14792 24760
rect 14476 24410 14504 24754
rect 14556 24608 14608 24614
rect 14752 24585 14780 24754
rect 14556 24550 14608 24556
rect 14738 24576 14794 24585
rect 14464 24404 14516 24410
rect 14464 24346 14516 24352
rect 14568 24206 14596 24550
rect 14738 24511 14794 24520
rect 14752 24274 14780 24511
rect 14740 24268 14792 24274
rect 14740 24210 14792 24216
rect 14556 24200 14608 24206
rect 14556 24142 14608 24148
rect 14648 23724 14700 23730
rect 14648 23666 14700 23672
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14280 22976 14332 22982
rect 14280 22918 14332 22924
rect 14292 22778 14320 22918
rect 14280 22772 14332 22778
rect 14280 22714 14332 22720
rect 14188 22704 14240 22710
rect 14188 22646 14240 22652
rect 14556 22432 14608 22438
rect 14556 22374 14608 22380
rect 14016 22066 14136 22094
rect 14370 22128 14426 22137
rect 14016 22030 14044 22066
rect 14370 22063 14426 22072
rect 14384 22030 14412 22063
rect 14004 22024 14056 22030
rect 14004 21966 14056 21972
rect 14372 22024 14424 22030
rect 14372 21966 14424 21972
rect 13912 21616 13964 21622
rect 13912 21558 13964 21564
rect 13820 20936 13872 20942
rect 13820 20878 13872 20884
rect 13832 20466 13860 20878
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 13924 20534 13952 20742
rect 13912 20528 13964 20534
rect 13912 20470 13964 20476
rect 13820 20460 13872 20466
rect 13820 20402 13872 20408
rect 13924 19802 13952 20470
rect 13832 19786 13952 19802
rect 13820 19780 13952 19786
rect 13872 19774 13952 19780
rect 13820 19722 13872 19728
rect 14016 18170 14044 21966
rect 14384 21554 14412 21966
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 14372 20800 14424 20806
rect 14372 20742 14424 20748
rect 14280 20528 14332 20534
rect 14280 20470 14332 20476
rect 14188 20392 14240 20398
rect 14188 20334 14240 20340
rect 14096 20256 14148 20262
rect 14096 20198 14148 20204
rect 14108 19378 14136 20198
rect 14200 20058 14228 20334
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 14186 19816 14242 19825
rect 14186 19751 14242 19760
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 14200 19242 14228 19751
rect 14292 19718 14320 20470
rect 14384 20466 14412 20742
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 14464 20460 14516 20466
rect 14464 20402 14516 20408
rect 14476 20058 14504 20402
rect 14464 20052 14516 20058
rect 14464 19994 14516 20000
rect 14370 19816 14426 19825
rect 14370 19751 14372 19760
rect 14424 19751 14426 19760
rect 14464 19780 14516 19786
rect 14372 19722 14424 19728
rect 14464 19722 14516 19728
rect 14280 19712 14332 19718
rect 14280 19654 14332 19660
rect 14292 19514 14320 19654
rect 14280 19508 14332 19514
rect 14280 19450 14332 19456
rect 14372 19372 14424 19378
rect 14476 19360 14504 19722
rect 14424 19332 14504 19360
rect 14372 19314 14424 19320
rect 14188 19236 14240 19242
rect 14188 19178 14240 19184
rect 14096 18692 14148 18698
rect 14096 18634 14148 18640
rect 14108 18358 14136 18634
rect 14200 18426 14228 19178
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14096 18352 14148 18358
rect 14096 18294 14148 18300
rect 13924 18142 14044 18170
rect 13818 17096 13874 17105
rect 13818 17031 13874 17040
rect 13832 16658 13860 17031
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13740 16510 13860 16538
rect 13832 16454 13860 16510
rect 13728 16448 13780 16454
rect 13728 16390 13780 16396
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13740 16266 13768 16390
rect 13740 16238 13860 16266
rect 13832 16114 13860 16238
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 13188 15026 13216 15438
rect 13280 15026 13308 15846
rect 13360 15360 13412 15366
rect 13360 15302 13412 15308
rect 13372 15162 13400 15302
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13452 15088 13504 15094
rect 13452 15030 13504 15036
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 13176 15020 13228 15026
rect 13176 14962 13228 14968
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 12084 12406 12204 12434
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 11612 7812 11664 7818
rect 11612 7754 11664 7760
rect 11796 7812 11848 7818
rect 11796 7754 11848 7760
rect 10612 7500 10732 7528
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 10612 5574 10640 7346
rect 10704 7342 10732 7500
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10704 5642 10732 6054
rect 10980 5794 11008 7414
rect 11518 6896 11574 6905
rect 11518 6831 11574 6840
rect 11532 6798 11560 6831
rect 11808 6798 11836 7754
rect 12084 7546 12112 12406
rect 12268 11694 12296 13330
rect 12360 13326 12388 13874
rect 12452 13870 12480 14962
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12360 12782 12388 13262
rect 12452 13190 12480 13670
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12452 12986 12480 13126
rect 12544 12986 12572 13942
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12808 13932 12860 13938
rect 12912 13920 12940 14758
rect 13464 14362 13492 15030
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 12992 14340 13044 14346
rect 12992 14282 13044 14288
rect 13280 14334 13492 14362
rect 13004 13938 13032 14282
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 13188 14074 13216 14214
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 12860 13892 12940 13920
rect 12808 13874 12860 13880
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 12360 11626 12388 12582
rect 12636 12238 12664 13874
rect 12716 13796 12768 13802
rect 12716 13738 12768 13744
rect 12728 13326 12756 13738
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 12820 13326 12848 13670
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12912 12238 12940 13892
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 13084 13728 13136 13734
rect 13004 13676 13084 13682
rect 13004 13670 13136 13676
rect 13004 13654 13124 13670
rect 13004 13190 13032 13654
rect 13188 13394 13216 14010
rect 13280 13938 13308 14334
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 13004 12850 13032 13126
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 13096 12442 13124 13262
rect 13176 13252 13228 13258
rect 13176 13194 13228 13200
rect 13188 12986 13216 13194
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 13280 12646 13308 13874
rect 13372 12714 13400 13874
rect 13360 12708 13412 12714
rect 13360 12650 13412 12656
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12898 12064 12954 12073
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 12348 11620 12400 11626
rect 12348 11562 12400 11568
rect 12176 11354 12204 11562
rect 12256 11552 12308 11558
rect 12308 11500 12388 11506
rect 12256 11494 12388 11500
rect 12268 11478 12388 11494
rect 12360 11354 12388 11478
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12440 11280 12492 11286
rect 12440 11222 12492 11228
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 12268 9654 12296 11018
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 12360 10742 12388 10950
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 12360 9722 12388 10678
rect 12452 10674 12480 11222
rect 12544 11150 12572 11630
rect 12820 11286 12848 12038
rect 12898 11999 12954 12008
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12636 10266 12664 10610
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12544 10118 12848 10146
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12256 9648 12308 9654
rect 12256 9590 12308 9596
rect 12268 9450 12296 9590
rect 12256 9444 12308 9450
rect 12256 9386 12308 9392
rect 12268 8974 12296 9386
rect 12360 8974 12388 9658
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 12268 6798 12296 8774
rect 12452 7546 12480 10066
rect 12544 9994 12572 10118
rect 12820 10062 12848 10118
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12532 9988 12584 9994
rect 12532 9930 12584 9936
rect 12544 9110 12572 9930
rect 12728 9518 12756 9998
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12820 9586 12848 9862
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 12544 8906 12572 9046
rect 12728 9042 12756 9454
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12912 8922 12940 11999
rect 12992 11824 13044 11830
rect 12992 11766 13044 11772
rect 13004 10674 13032 11766
rect 13096 11762 13124 12378
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 13464 11694 13492 14214
rect 13648 13870 13676 14758
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13740 12850 13768 13126
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13464 11150 13492 11494
rect 13832 11354 13860 13126
rect 13924 12238 13952 18142
rect 14200 17542 14228 18362
rect 14188 17536 14240 17542
rect 14188 17478 14240 17484
rect 14568 16674 14596 22374
rect 14660 17270 14688 23666
rect 14740 23248 14792 23254
rect 14740 23190 14792 23196
rect 14752 22409 14780 23190
rect 14738 22400 14794 22409
rect 14738 22335 14794 22344
rect 14740 22024 14792 22030
rect 14740 21966 14792 21972
rect 14752 21554 14780 21966
rect 14740 21548 14792 21554
rect 14740 21490 14792 21496
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 14752 19242 14780 21286
rect 14740 19236 14792 19242
rect 14740 19178 14792 19184
rect 14648 17264 14700 17270
rect 14648 17206 14700 17212
rect 14844 17218 14872 26250
rect 14936 25906 14964 26726
rect 14924 25900 14976 25906
rect 14924 25842 14976 25848
rect 14924 24336 14976 24342
rect 14924 24278 14976 24284
rect 14936 24138 14964 24278
rect 14924 24132 14976 24138
rect 14924 24074 14976 24080
rect 15028 21350 15056 27474
rect 15120 27130 15148 30194
rect 15304 29186 15332 30534
rect 15396 29322 15424 31214
rect 15488 30938 15516 31282
rect 15660 31272 15712 31278
rect 15660 31214 15712 31220
rect 15476 30932 15528 30938
rect 15476 30874 15528 30880
rect 15488 30190 15516 30874
rect 15672 30734 15700 31214
rect 15568 30728 15620 30734
rect 15566 30696 15568 30705
rect 15660 30728 15712 30734
rect 15620 30696 15622 30705
rect 15660 30670 15712 30676
rect 15566 30631 15622 30640
rect 15672 30326 15700 30670
rect 15660 30320 15712 30326
rect 15660 30262 15712 30268
rect 15568 30252 15620 30258
rect 15568 30194 15620 30200
rect 15476 30184 15528 30190
rect 15476 30126 15528 30132
rect 15580 30054 15608 30194
rect 15658 30152 15714 30161
rect 15658 30087 15714 30096
rect 15568 30048 15620 30054
rect 15568 29990 15620 29996
rect 15474 29744 15530 29753
rect 15474 29679 15476 29688
rect 15528 29679 15530 29688
rect 15476 29650 15528 29656
rect 15396 29294 15516 29322
rect 15304 29158 15424 29186
rect 15292 29096 15344 29102
rect 15292 29038 15344 29044
rect 15200 28076 15252 28082
rect 15200 28018 15252 28024
rect 15212 27606 15240 28018
rect 15200 27600 15252 27606
rect 15200 27542 15252 27548
rect 15108 27124 15160 27130
rect 15108 27066 15160 27072
rect 15108 26920 15160 26926
rect 15108 26862 15160 26868
rect 15120 25838 15148 26862
rect 15108 25832 15160 25838
rect 15108 25774 15160 25780
rect 15120 25498 15148 25774
rect 15212 25770 15240 27542
rect 15304 27130 15332 29038
rect 15292 27124 15344 27130
rect 15292 27066 15344 27072
rect 15292 26988 15344 26994
rect 15396 26976 15424 29158
rect 15488 28370 15516 29294
rect 15580 28694 15608 29990
rect 15568 28688 15620 28694
rect 15568 28630 15620 28636
rect 15488 28342 15608 28370
rect 15476 28212 15528 28218
rect 15476 28154 15528 28160
rect 15488 27470 15516 28154
rect 15476 27464 15528 27470
rect 15580 27441 15608 28342
rect 15476 27406 15528 27412
rect 15566 27432 15622 27441
rect 15566 27367 15622 27376
rect 15344 26948 15424 26976
rect 15292 26930 15344 26936
rect 15200 25764 15252 25770
rect 15200 25706 15252 25712
rect 15108 25492 15160 25498
rect 15108 25434 15160 25440
rect 15200 24744 15252 24750
rect 15200 24686 15252 24692
rect 15212 23730 15240 24686
rect 15304 24206 15332 26930
rect 15476 26512 15528 26518
rect 15672 26489 15700 30087
rect 15764 29646 15792 36128
rect 15844 36032 15896 36038
rect 15844 35974 15896 35980
rect 15856 35698 15884 35974
rect 15844 35692 15896 35698
rect 15844 35634 15896 35640
rect 15856 35494 15884 35634
rect 15844 35488 15896 35494
rect 15844 35430 15896 35436
rect 15844 35012 15896 35018
rect 15844 34954 15896 34960
rect 15856 33046 15884 34954
rect 15844 33040 15896 33046
rect 15844 32982 15896 32988
rect 15844 32564 15896 32570
rect 15844 32506 15896 32512
rect 15752 29640 15804 29646
rect 15752 29582 15804 29588
rect 15764 28150 15792 29582
rect 15856 29170 15884 32506
rect 15948 30054 15976 39238
rect 16592 38418 16620 39374
rect 16672 39296 16724 39302
rect 16672 39238 16724 39244
rect 16684 39030 16712 39238
rect 16672 39024 16724 39030
rect 16672 38966 16724 38972
rect 16580 38412 16632 38418
rect 16580 38354 16632 38360
rect 16764 37732 16816 37738
rect 16764 37674 16816 37680
rect 16028 37120 16080 37126
rect 16028 37062 16080 37068
rect 16040 36786 16068 37062
rect 16120 36916 16172 36922
rect 16120 36858 16172 36864
rect 16132 36786 16160 36858
rect 16028 36780 16080 36786
rect 16028 36722 16080 36728
rect 16120 36780 16172 36786
rect 16120 36722 16172 36728
rect 16132 36106 16160 36722
rect 16396 36168 16448 36174
rect 16396 36110 16448 36116
rect 16120 36100 16172 36106
rect 16120 36042 16172 36048
rect 16304 36100 16356 36106
rect 16304 36042 16356 36048
rect 16132 35714 16160 36042
rect 16316 35834 16344 36042
rect 16304 35828 16356 35834
rect 16304 35770 16356 35776
rect 16040 35698 16160 35714
rect 16028 35692 16160 35698
rect 16080 35686 16160 35692
rect 16028 35634 16080 35640
rect 16120 35624 16172 35630
rect 16120 35566 16172 35572
rect 16132 35290 16160 35566
rect 16212 35556 16264 35562
rect 16212 35498 16264 35504
rect 16304 35556 16356 35562
rect 16304 35498 16356 35504
rect 16120 35284 16172 35290
rect 16120 35226 16172 35232
rect 16028 34604 16080 34610
rect 16028 34546 16080 34552
rect 16040 32774 16068 34546
rect 16120 33584 16172 33590
rect 16120 33526 16172 33532
rect 16132 32910 16160 33526
rect 16120 32904 16172 32910
rect 16120 32846 16172 32852
rect 16028 32768 16080 32774
rect 16028 32710 16080 32716
rect 16120 32496 16172 32502
rect 16120 32438 16172 32444
rect 16224 32450 16252 35498
rect 16316 35154 16344 35498
rect 16304 35148 16356 35154
rect 16304 35090 16356 35096
rect 16408 35018 16436 36110
rect 16672 35624 16724 35630
rect 16672 35566 16724 35572
rect 16684 35290 16712 35566
rect 16672 35284 16724 35290
rect 16672 35226 16724 35232
rect 16684 35018 16712 35226
rect 16396 35012 16448 35018
rect 16396 34954 16448 34960
rect 16672 35012 16724 35018
rect 16672 34954 16724 34960
rect 16580 34128 16632 34134
rect 16580 34070 16632 34076
rect 16304 33856 16356 33862
rect 16304 33798 16356 33804
rect 16316 33454 16344 33798
rect 16396 33652 16448 33658
rect 16396 33594 16448 33600
rect 16304 33448 16356 33454
rect 16304 33390 16356 33396
rect 16316 32586 16344 33390
rect 16408 32774 16436 33594
rect 16486 33008 16542 33017
rect 16486 32943 16542 32952
rect 16500 32910 16528 32943
rect 16488 32904 16540 32910
rect 16488 32846 16540 32852
rect 16396 32768 16448 32774
rect 16396 32710 16448 32716
rect 16316 32558 16528 32586
rect 16132 31890 16160 32438
rect 16224 32422 16436 32450
rect 16212 32360 16264 32366
rect 16212 32302 16264 32308
rect 16120 31884 16172 31890
rect 16120 31826 16172 31832
rect 16132 31793 16160 31826
rect 16118 31784 16174 31793
rect 16118 31719 16174 31728
rect 16028 31340 16080 31346
rect 16028 31282 16080 31288
rect 16040 31142 16068 31282
rect 16028 31136 16080 31142
rect 16080 31096 16160 31124
rect 16028 31078 16080 31084
rect 16028 30252 16080 30258
rect 16028 30194 16080 30200
rect 16040 30161 16068 30194
rect 16026 30152 16082 30161
rect 16026 30087 16082 30096
rect 15936 30048 15988 30054
rect 15936 29990 15988 29996
rect 16028 30048 16080 30054
rect 16028 29990 16080 29996
rect 16040 29238 16068 29990
rect 16028 29232 16080 29238
rect 16028 29174 16080 29180
rect 15844 29164 15896 29170
rect 15844 29106 15896 29112
rect 15752 28144 15804 28150
rect 15752 28086 15804 28092
rect 15752 28008 15804 28014
rect 15752 27950 15804 27956
rect 15764 27674 15792 27950
rect 15752 27668 15804 27674
rect 15752 27610 15804 27616
rect 15764 27470 15792 27610
rect 15856 27538 15884 29106
rect 16028 28960 16080 28966
rect 16028 28902 16080 28908
rect 16040 28150 16068 28902
rect 16132 28422 16160 31096
rect 16224 30240 16252 32302
rect 16408 31822 16436 32422
rect 16304 31816 16356 31822
rect 16304 31758 16356 31764
rect 16396 31816 16448 31822
rect 16396 31758 16448 31764
rect 16316 31210 16344 31758
rect 16304 31204 16356 31210
rect 16304 31146 16356 31152
rect 16304 30252 16356 30258
rect 16224 30212 16304 30240
rect 16304 30194 16356 30200
rect 16316 29850 16344 30194
rect 16304 29844 16356 29850
rect 16304 29786 16356 29792
rect 16302 29744 16358 29753
rect 16302 29679 16358 29688
rect 16120 28416 16172 28422
rect 16120 28358 16172 28364
rect 16028 28144 16080 28150
rect 16028 28086 16080 28092
rect 16120 27872 16172 27878
rect 16120 27814 16172 27820
rect 15844 27532 15896 27538
rect 15844 27474 15896 27480
rect 15936 27532 15988 27538
rect 15936 27474 15988 27480
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 15844 27124 15896 27130
rect 15948 27112 15976 27474
rect 16028 27328 16080 27334
rect 16028 27270 16080 27276
rect 15896 27084 15976 27112
rect 15844 27066 15896 27072
rect 15476 26454 15528 26460
rect 15658 26480 15714 26489
rect 15488 26246 15516 26454
rect 15658 26415 15714 26424
rect 15856 26382 15884 27066
rect 16040 26382 16068 27270
rect 16132 26382 16160 27814
rect 16212 27328 16264 27334
rect 16212 27270 16264 27276
rect 16224 26994 16252 27270
rect 16212 26988 16264 26994
rect 16212 26930 16264 26936
rect 16316 26382 16344 29679
rect 16408 28762 16436 31758
rect 16500 30598 16528 32558
rect 16488 30592 16540 30598
rect 16488 30534 16540 30540
rect 16592 30054 16620 34070
rect 16672 33652 16724 33658
rect 16672 33594 16724 33600
rect 16684 32842 16712 33594
rect 16672 32836 16724 32842
rect 16672 32778 16724 32784
rect 16776 31906 16804 37674
rect 16868 35086 16896 39850
rect 16948 39840 17000 39846
rect 16948 39782 17000 39788
rect 16960 38962 16988 39782
rect 17052 39506 17080 40598
rect 17132 40044 17184 40050
rect 17132 39986 17184 39992
rect 17040 39500 17092 39506
rect 17040 39442 17092 39448
rect 17144 39438 17172 39986
rect 17868 39908 17920 39914
rect 17868 39850 17920 39856
rect 17880 39506 17908 39850
rect 17868 39500 17920 39506
rect 17868 39442 17920 39448
rect 17132 39432 17184 39438
rect 17132 39374 17184 39380
rect 18052 39364 18104 39370
rect 18052 39306 18104 39312
rect 17960 39296 18012 39302
rect 17960 39238 18012 39244
rect 16948 38956 17000 38962
rect 16948 38898 17000 38904
rect 17972 38350 18000 39238
rect 18064 39030 18092 39306
rect 20720 39092 20772 39098
rect 20720 39034 20772 39040
rect 18052 39024 18104 39030
rect 18052 38966 18104 38972
rect 18328 39024 18380 39030
rect 18328 38966 18380 38972
rect 18340 38350 18368 38966
rect 19800 38888 19852 38894
rect 19800 38830 19852 38836
rect 20076 38888 20128 38894
rect 20076 38830 20128 38836
rect 19064 38752 19116 38758
rect 19064 38694 19116 38700
rect 17776 38344 17828 38350
rect 17776 38286 17828 38292
rect 17960 38344 18012 38350
rect 17960 38286 18012 38292
rect 18052 38344 18104 38350
rect 18052 38286 18104 38292
rect 18328 38344 18380 38350
rect 18328 38286 18380 38292
rect 17788 38010 17816 38286
rect 17776 38004 17828 38010
rect 17776 37946 17828 37952
rect 17408 37868 17460 37874
rect 17408 37810 17460 37816
rect 17684 37868 17736 37874
rect 17684 37810 17736 37816
rect 17316 37800 17368 37806
rect 17316 37742 17368 37748
rect 17328 37466 17356 37742
rect 17316 37460 17368 37466
rect 17316 37402 17368 37408
rect 17420 37398 17448 37810
rect 17696 37466 17724 37810
rect 18064 37806 18092 38286
rect 18512 38276 18564 38282
rect 18512 38218 18564 38224
rect 18328 38208 18380 38214
rect 18328 38150 18380 38156
rect 18144 37868 18196 37874
rect 18144 37810 18196 37816
rect 18052 37800 18104 37806
rect 18052 37742 18104 37748
rect 17684 37460 17736 37466
rect 17684 37402 17736 37408
rect 17408 37392 17460 37398
rect 17408 37334 17460 37340
rect 17224 37324 17276 37330
rect 17224 37266 17276 37272
rect 17132 36780 17184 36786
rect 17132 36722 17184 36728
rect 17144 36038 17172 36722
rect 17236 36242 17264 37266
rect 17224 36236 17276 36242
rect 17276 36196 17356 36224
rect 17224 36178 17276 36184
rect 17132 36032 17184 36038
rect 17132 35974 17184 35980
rect 17328 35834 17356 36196
rect 17316 35828 17368 35834
rect 17144 35788 17316 35816
rect 17040 35216 17092 35222
rect 17040 35158 17092 35164
rect 16856 35080 16908 35086
rect 16856 35022 16908 35028
rect 17052 32434 17080 35158
rect 17144 34066 17172 35788
rect 17316 35770 17368 35776
rect 17420 35562 17448 37334
rect 17696 37262 17724 37402
rect 18052 37392 18104 37398
rect 18156 37380 18184 37810
rect 18104 37352 18184 37380
rect 18052 37334 18104 37340
rect 17684 37256 17736 37262
rect 17684 37198 17736 37204
rect 17776 37256 17828 37262
rect 17776 37198 17828 37204
rect 17960 37256 18012 37262
rect 17960 37198 18012 37204
rect 17788 36718 17816 37198
rect 17868 37188 17920 37194
rect 17868 37130 17920 37136
rect 17776 36712 17828 36718
rect 17776 36654 17828 36660
rect 17880 36666 17908 37130
rect 17972 36786 18000 37198
rect 18064 36786 18092 37334
rect 18236 37256 18288 37262
rect 18236 37198 18288 37204
rect 18248 36922 18276 37198
rect 18236 36916 18288 36922
rect 18236 36858 18288 36864
rect 17960 36780 18012 36786
rect 17960 36722 18012 36728
rect 18052 36780 18104 36786
rect 18052 36722 18104 36728
rect 17880 36650 18000 36666
rect 17880 36644 18012 36650
rect 17880 36638 17960 36644
rect 17960 36586 18012 36592
rect 18052 36372 18104 36378
rect 18052 36314 18104 36320
rect 17960 36032 18012 36038
rect 17960 35974 18012 35980
rect 17972 35766 18000 35974
rect 17960 35760 18012 35766
rect 17960 35702 18012 35708
rect 17500 35692 17552 35698
rect 17500 35634 17552 35640
rect 17512 35601 17540 35634
rect 17972 35630 18000 35702
rect 18064 35630 18092 36314
rect 18248 36174 18276 36858
rect 18236 36168 18288 36174
rect 18236 36110 18288 36116
rect 17960 35624 18012 35630
rect 17498 35592 17554 35601
rect 17408 35556 17460 35562
rect 18052 35624 18104 35630
rect 17960 35566 18012 35572
rect 18050 35592 18052 35601
rect 18104 35592 18106 35601
rect 17498 35527 17554 35536
rect 17408 35498 17460 35504
rect 17408 35216 17460 35222
rect 17408 35158 17460 35164
rect 17512 35170 17540 35527
rect 17316 35012 17368 35018
rect 17316 34954 17368 34960
rect 17328 34610 17356 34954
rect 17420 34746 17448 35158
rect 17512 35154 17724 35170
rect 17500 35148 17724 35154
rect 17552 35142 17724 35148
rect 17500 35090 17552 35096
rect 17696 35086 17724 35142
rect 17972 35086 18000 35566
rect 18050 35527 18106 35536
rect 18236 35488 18288 35494
rect 18236 35430 18288 35436
rect 17684 35080 17736 35086
rect 17684 35022 17736 35028
rect 17960 35080 18012 35086
rect 17960 35022 18012 35028
rect 17776 35012 17828 35018
rect 17776 34954 17828 34960
rect 17500 34944 17552 34950
rect 17500 34886 17552 34892
rect 17512 34746 17540 34886
rect 17408 34740 17460 34746
rect 17408 34682 17460 34688
rect 17500 34740 17552 34746
rect 17500 34682 17552 34688
rect 17788 34678 17816 34954
rect 17776 34672 17828 34678
rect 17776 34614 17828 34620
rect 18248 34610 18276 35430
rect 17316 34604 17368 34610
rect 17316 34546 17368 34552
rect 18236 34604 18288 34610
rect 18236 34546 18288 34552
rect 17684 34468 17736 34474
rect 17684 34410 17736 34416
rect 17408 34400 17460 34406
rect 17408 34342 17460 34348
rect 17132 34060 17184 34066
rect 17132 34002 17184 34008
rect 17144 33590 17172 34002
rect 17420 33998 17448 34342
rect 17408 33992 17460 33998
rect 17408 33934 17460 33940
rect 17592 33856 17644 33862
rect 17592 33798 17644 33804
rect 17132 33584 17184 33590
rect 17132 33526 17184 33532
rect 17224 33448 17276 33454
rect 17224 33390 17276 33396
rect 17040 32428 17092 32434
rect 17040 32370 17092 32376
rect 17236 32026 17264 33390
rect 17604 32910 17632 33798
rect 17696 33454 17724 34410
rect 18144 34400 18196 34406
rect 18144 34342 18196 34348
rect 18156 33998 18184 34342
rect 18248 34134 18276 34546
rect 18340 34202 18368 38150
rect 18524 35834 18552 38218
rect 18972 37868 19024 37874
rect 18972 37810 19024 37816
rect 18604 37664 18656 37670
rect 18604 37606 18656 37612
rect 18616 37330 18644 37606
rect 18604 37324 18656 37330
rect 18604 37266 18656 37272
rect 18696 37120 18748 37126
rect 18696 37062 18748 37068
rect 18708 36786 18736 37062
rect 18984 36922 19012 37810
rect 19076 37330 19104 38694
rect 19812 38554 19840 38830
rect 19800 38548 19852 38554
rect 19800 38490 19852 38496
rect 19892 38548 19944 38554
rect 19892 38490 19944 38496
rect 19248 38344 19300 38350
rect 19248 38286 19300 38292
rect 19260 37942 19288 38286
rect 19340 38208 19392 38214
rect 19340 38150 19392 38156
rect 19248 37936 19300 37942
rect 19248 37878 19300 37884
rect 19352 37874 19380 38150
rect 19156 37868 19208 37874
rect 19156 37810 19208 37816
rect 19340 37868 19392 37874
rect 19340 37810 19392 37816
rect 19168 37466 19196 37810
rect 19248 37800 19300 37806
rect 19248 37742 19300 37748
rect 19156 37460 19208 37466
rect 19156 37402 19208 37408
rect 19260 37346 19288 37742
rect 19064 37324 19116 37330
rect 19064 37266 19116 37272
rect 19168 37318 19288 37346
rect 18972 36916 19024 36922
rect 18972 36858 19024 36864
rect 18696 36780 18748 36786
rect 18696 36722 18748 36728
rect 18788 36576 18840 36582
rect 18788 36518 18840 36524
rect 18800 36242 18828 36518
rect 18788 36236 18840 36242
rect 18788 36178 18840 36184
rect 18512 35828 18564 35834
rect 18512 35770 18564 35776
rect 19064 35828 19116 35834
rect 19064 35770 19116 35776
rect 18512 35692 18564 35698
rect 18512 35634 18564 35640
rect 18524 35222 18552 35634
rect 18512 35216 18564 35222
rect 18512 35158 18564 35164
rect 18880 35216 18932 35222
rect 18880 35158 18932 35164
rect 18694 35048 18750 35057
rect 18694 34983 18696 34992
rect 18748 34983 18750 34992
rect 18696 34954 18748 34960
rect 18512 34944 18564 34950
rect 18512 34886 18564 34892
rect 18788 34944 18840 34950
rect 18788 34886 18840 34892
rect 18524 34746 18552 34886
rect 18800 34746 18828 34886
rect 18512 34740 18564 34746
rect 18512 34682 18564 34688
rect 18788 34740 18840 34746
rect 18788 34682 18840 34688
rect 18328 34196 18380 34202
rect 18328 34138 18380 34144
rect 18236 34128 18288 34134
rect 18236 34070 18288 34076
rect 18144 33992 18196 33998
rect 18340 33946 18368 34138
rect 18524 33998 18552 34682
rect 18604 34604 18656 34610
rect 18604 34546 18656 34552
rect 18616 34202 18644 34546
rect 18604 34196 18656 34202
rect 18604 34138 18656 34144
rect 18892 34066 18920 35158
rect 19076 34678 19104 35770
rect 19168 35630 19196 37318
rect 19340 37256 19392 37262
rect 19340 37198 19392 37204
rect 19708 37256 19760 37262
rect 19708 37198 19760 37204
rect 19352 36582 19380 37198
rect 19432 37120 19484 37126
rect 19432 37062 19484 37068
rect 19444 36718 19472 37062
rect 19432 36712 19484 36718
rect 19432 36654 19484 36660
rect 19340 36576 19392 36582
rect 19340 36518 19392 36524
rect 19248 36236 19300 36242
rect 19248 36178 19300 36184
rect 19260 35698 19288 36178
rect 19616 36168 19668 36174
rect 19616 36110 19668 36116
rect 19432 35828 19484 35834
rect 19432 35770 19484 35776
rect 19444 35698 19472 35770
rect 19248 35692 19300 35698
rect 19248 35634 19300 35640
rect 19432 35692 19484 35698
rect 19432 35634 19484 35640
rect 19524 35692 19576 35698
rect 19524 35634 19576 35640
rect 19156 35624 19208 35630
rect 19156 35566 19208 35572
rect 19248 35284 19300 35290
rect 19248 35226 19300 35232
rect 19064 34672 19116 34678
rect 19064 34614 19116 34620
rect 19076 34406 19104 34614
rect 19260 34610 19288 35226
rect 19248 34604 19300 34610
rect 19168 34564 19248 34592
rect 19064 34400 19116 34406
rect 19064 34342 19116 34348
rect 18880 34060 18932 34066
rect 18880 34002 18932 34008
rect 18144 33934 18196 33940
rect 18156 33658 18184 33934
rect 18248 33918 18368 33946
rect 18512 33992 18564 33998
rect 18512 33934 18564 33940
rect 18248 33658 18276 33918
rect 18328 33856 18380 33862
rect 18328 33798 18380 33804
rect 18144 33652 18196 33658
rect 18144 33594 18196 33600
rect 18236 33652 18288 33658
rect 18236 33594 18288 33600
rect 17684 33448 17736 33454
rect 17684 33390 17736 33396
rect 17960 33448 18012 33454
rect 17960 33390 18012 33396
rect 17972 33114 18000 33390
rect 18144 33312 18196 33318
rect 18144 33254 18196 33260
rect 17960 33108 18012 33114
rect 17960 33050 18012 33056
rect 18156 32910 18184 33254
rect 18340 32978 18368 33798
rect 18604 33652 18656 33658
rect 18604 33594 18656 33600
rect 18512 33448 18564 33454
rect 18512 33390 18564 33396
rect 18328 32972 18380 32978
rect 18328 32914 18380 32920
rect 17592 32904 17644 32910
rect 17592 32846 17644 32852
rect 18144 32904 18196 32910
rect 18144 32846 18196 32852
rect 18236 32904 18288 32910
rect 18236 32846 18288 32852
rect 18156 32570 18184 32846
rect 18144 32564 18196 32570
rect 18144 32506 18196 32512
rect 18248 32502 18276 32846
rect 18236 32496 18288 32502
rect 18236 32438 18288 32444
rect 17224 32020 17276 32026
rect 17224 31962 17276 31968
rect 16684 31878 16804 31906
rect 17236 31890 17264 31962
rect 17224 31884 17276 31890
rect 16684 30802 16712 31878
rect 17224 31826 17276 31832
rect 18052 31884 18104 31890
rect 18052 31826 18104 31832
rect 16764 31748 16816 31754
rect 16764 31690 16816 31696
rect 17960 31748 18012 31754
rect 17960 31690 18012 31696
rect 16776 31482 16804 31690
rect 16764 31476 16816 31482
rect 16764 31418 16816 31424
rect 16948 31340 17000 31346
rect 16948 31282 17000 31288
rect 17500 31340 17552 31346
rect 17500 31282 17552 31288
rect 16672 30796 16724 30802
rect 16672 30738 16724 30744
rect 16764 30252 16816 30258
rect 16684 30212 16764 30240
rect 16580 30048 16632 30054
rect 16580 29990 16632 29996
rect 16488 29640 16540 29646
rect 16684 29628 16712 30212
rect 16764 30194 16816 30200
rect 16960 30122 16988 31282
rect 17224 31272 17276 31278
rect 17224 31214 17276 31220
rect 17132 30252 17184 30258
rect 17132 30194 17184 30200
rect 16948 30116 17000 30122
rect 16948 30058 17000 30064
rect 16764 30048 16816 30054
rect 16764 29990 16816 29996
rect 16540 29600 16712 29628
rect 16488 29582 16540 29588
rect 16500 29170 16528 29582
rect 16776 29578 16804 29990
rect 16960 29646 16988 30058
rect 17040 30048 17092 30054
rect 17040 29990 17092 29996
rect 16948 29640 17000 29646
rect 16948 29582 17000 29588
rect 16764 29572 16816 29578
rect 16764 29514 16816 29520
rect 16764 29300 16816 29306
rect 16764 29242 16816 29248
rect 16488 29164 16540 29170
rect 16488 29106 16540 29112
rect 16776 29102 16804 29242
rect 16764 29096 16816 29102
rect 16764 29038 16816 29044
rect 16960 29034 16988 29582
rect 17052 29170 17080 29990
rect 17144 29646 17172 30194
rect 17132 29640 17184 29646
rect 17132 29582 17184 29588
rect 17040 29164 17092 29170
rect 17040 29106 17092 29112
rect 16948 29028 17000 29034
rect 16948 28970 17000 28976
rect 16396 28756 16448 28762
rect 16396 28698 16448 28704
rect 16960 28626 16988 28970
rect 16948 28620 17000 28626
rect 16948 28562 17000 28568
rect 16672 28076 16724 28082
rect 16672 28018 16724 28024
rect 16684 27606 16712 28018
rect 16672 27600 16724 27606
rect 16672 27542 16724 27548
rect 16486 27160 16542 27169
rect 16486 27095 16488 27104
rect 16540 27095 16542 27104
rect 16488 27066 16540 27072
rect 16764 26988 16816 26994
rect 16764 26930 16816 26936
rect 16948 26988 17000 26994
rect 16948 26930 17000 26936
rect 16396 26920 16448 26926
rect 16396 26862 16448 26868
rect 16408 26382 16436 26862
rect 16776 26382 16804 26930
rect 16854 26480 16910 26489
rect 16854 26415 16910 26424
rect 15844 26376 15896 26382
rect 15658 26344 15714 26353
rect 15844 26318 15896 26324
rect 16028 26376 16080 26382
rect 16028 26318 16080 26324
rect 16120 26376 16172 26382
rect 16120 26318 16172 26324
rect 16304 26376 16356 26382
rect 16304 26318 16356 26324
rect 16396 26376 16448 26382
rect 16396 26318 16448 26324
rect 16764 26376 16816 26382
rect 16764 26318 16816 26324
rect 15658 26279 15660 26288
rect 15712 26279 15714 26288
rect 15660 26250 15712 26256
rect 15384 26240 15436 26246
rect 15384 26182 15436 26188
rect 15476 26240 15528 26246
rect 15476 26182 15528 26188
rect 15396 25974 15424 26182
rect 15384 25968 15436 25974
rect 15384 25910 15436 25916
rect 15660 25492 15712 25498
rect 15660 25434 15712 25440
rect 15476 25152 15528 25158
rect 15476 25094 15528 25100
rect 15488 24818 15516 25094
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 15488 24342 15516 24754
rect 15672 24750 15700 25434
rect 15856 25362 15884 26318
rect 16212 26240 16264 26246
rect 16212 26182 16264 26188
rect 16028 25832 16080 25838
rect 16028 25774 16080 25780
rect 15844 25356 15896 25362
rect 15844 25298 15896 25304
rect 15752 24948 15804 24954
rect 15752 24890 15804 24896
rect 15660 24744 15712 24750
rect 15660 24686 15712 24692
rect 15672 24410 15700 24686
rect 15660 24404 15712 24410
rect 15660 24346 15712 24352
rect 15476 24336 15528 24342
rect 15476 24278 15528 24284
rect 15292 24200 15344 24206
rect 15292 24142 15344 24148
rect 15476 24200 15528 24206
rect 15476 24142 15528 24148
rect 15488 23730 15516 24142
rect 15672 23730 15700 24346
rect 15764 24342 15792 24890
rect 15936 24676 15988 24682
rect 15936 24618 15988 24624
rect 15752 24336 15804 24342
rect 15752 24278 15804 24284
rect 15948 24070 15976 24618
rect 15936 24064 15988 24070
rect 15936 24006 15988 24012
rect 15200 23724 15252 23730
rect 15200 23666 15252 23672
rect 15476 23724 15528 23730
rect 15476 23666 15528 23672
rect 15660 23724 15712 23730
rect 15660 23666 15712 23672
rect 15488 23526 15516 23666
rect 15948 23526 15976 24006
rect 15476 23520 15528 23526
rect 15476 23462 15528 23468
rect 15936 23520 15988 23526
rect 15936 23462 15988 23468
rect 15382 23352 15438 23361
rect 15382 23287 15438 23296
rect 15108 21412 15160 21418
rect 15108 21354 15160 21360
rect 15016 21344 15068 21350
rect 15016 21286 15068 21292
rect 15120 20398 15148 21354
rect 15016 20392 15068 20398
rect 15016 20334 15068 20340
rect 15108 20392 15160 20398
rect 15108 20334 15160 20340
rect 14922 19952 14978 19961
rect 14922 19887 14978 19896
rect 14936 19854 14964 19887
rect 14924 19848 14976 19854
rect 14924 19790 14976 19796
rect 15028 19718 15056 20334
rect 15396 20058 15424 23287
rect 15476 21140 15528 21146
rect 15476 21082 15528 21088
rect 15488 21010 15516 21082
rect 15476 21004 15528 21010
rect 15476 20946 15528 20952
rect 15488 20466 15516 20946
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15476 20460 15528 20466
rect 15476 20402 15528 20408
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 15396 19854 15424 19994
rect 15488 19990 15516 20402
rect 15476 19984 15528 19990
rect 15580 19961 15608 20402
rect 15672 20330 15700 20878
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15660 20324 15712 20330
rect 15660 20266 15712 20272
rect 15476 19926 15528 19932
rect 15566 19952 15622 19961
rect 15566 19887 15622 19896
rect 15292 19848 15344 19854
rect 15290 19816 15292 19825
rect 15384 19848 15436 19854
rect 15344 19816 15346 19825
rect 15384 19790 15436 19796
rect 15290 19751 15346 19760
rect 15304 19718 15332 19751
rect 15016 19712 15068 19718
rect 15016 19654 15068 19660
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 15028 19514 15056 19654
rect 15304 19514 15332 19654
rect 15016 19508 15068 19514
rect 15016 19450 15068 19456
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 15292 19372 15344 19378
rect 15396 19360 15424 19790
rect 15580 19514 15608 19887
rect 15672 19854 15700 20266
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15568 19508 15620 19514
rect 15568 19450 15620 19456
rect 15764 19446 15792 20402
rect 15752 19440 15804 19446
rect 15752 19382 15804 19388
rect 15344 19332 15424 19360
rect 15292 19314 15344 19320
rect 15764 18850 15792 19382
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 15856 18970 15884 19314
rect 15936 19168 15988 19174
rect 15936 19110 15988 19116
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 15764 18822 15884 18850
rect 15566 18320 15622 18329
rect 15566 18255 15568 18264
rect 15620 18255 15622 18264
rect 15568 18226 15620 18232
rect 15476 18148 15528 18154
rect 15476 18090 15528 18096
rect 14844 17190 14964 17218
rect 14004 16652 14056 16658
rect 14004 16594 14056 16600
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 14476 16646 14596 16674
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 13924 11694 13952 12174
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13464 9586 13492 10406
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13188 9178 13216 9454
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 12636 8894 12940 8922
rect 12544 8498 12572 8842
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 11888 6724 11940 6730
rect 11888 6666 11940 6672
rect 11900 6458 11928 6666
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11992 6338 12020 6734
rect 10796 5778 11008 5794
rect 10784 5772 11008 5778
rect 10836 5766 11008 5772
rect 10784 5714 10836 5720
rect 10692 5636 10744 5642
rect 10692 5578 10744 5584
rect 10600 5568 10652 5574
rect 10600 5510 10652 5516
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 10612 3398 10640 5510
rect 10980 5234 11008 5766
rect 11900 6310 12020 6338
rect 11336 5568 11388 5574
rect 11336 5510 11388 5516
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10980 3602 11008 5170
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 11072 3466 11100 3878
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 11348 2446 11376 5510
rect 11612 4480 11664 4486
rect 11612 4422 11664 4428
rect 11624 4282 11652 4422
rect 11612 4276 11664 4282
rect 11612 4218 11664 4224
rect 11900 4214 11928 6310
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12268 5574 12296 6190
rect 12256 5568 12308 5574
rect 12256 5510 12308 5516
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 12084 4826 12112 5102
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 12360 4622 12388 7482
rect 12530 7440 12586 7449
rect 12636 7410 12664 8894
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12530 7375 12586 7384
rect 12624 7404 12676 7410
rect 12544 7342 12572 7375
rect 12624 7346 12676 7352
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 12544 6798 12572 7278
rect 12728 7002 12756 8026
rect 14016 7886 14044 16594
rect 14096 16584 14148 16590
rect 14096 16526 14148 16532
rect 14108 16182 14136 16526
rect 14188 16448 14240 16454
rect 14188 16390 14240 16396
rect 14096 16176 14148 16182
rect 14096 16118 14148 16124
rect 14200 15910 14228 16390
rect 14384 16046 14412 16594
rect 14476 16590 14504 16646
rect 14464 16584 14516 16590
rect 14464 16526 14516 16532
rect 14556 16584 14608 16590
rect 14556 16526 14608 16532
rect 14568 16182 14596 16526
rect 14464 16176 14516 16182
rect 14464 16118 14516 16124
rect 14556 16176 14608 16182
rect 14556 16118 14608 16124
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14476 15994 14504 16118
rect 14476 15966 14596 15994
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 14108 12646 14136 13670
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14384 12850 14412 13262
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 14384 11150 14412 12786
rect 14476 11898 14504 13874
rect 14568 12850 14596 15966
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14752 14618 14780 14758
rect 14740 14612 14792 14618
rect 14740 14554 14792 14560
rect 14752 13394 14780 14554
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14568 12306 14596 12786
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14844 12102 14872 14826
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14384 9994 14412 11086
rect 14740 10736 14792 10742
rect 14740 10678 14792 10684
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14372 9988 14424 9994
rect 14372 9930 14424 9936
rect 14384 9586 14412 9930
rect 14476 9722 14504 10610
rect 14752 10470 14780 10678
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14936 10266 14964 17190
rect 15198 17096 15254 17105
rect 15198 17031 15254 17040
rect 15016 16652 15068 16658
rect 15016 16594 15068 16600
rect 15028 10554 15056 16594
rect 15212 16130 15240 17031
rect 15120 16114 15240 16130
rect 15108 16108 15240 16114
rect 15160 16102 15240 16108
rect 15108 16050 15160 16056
rect 15120 15026 15148 16050
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 15212 13326 15240 13738
rect 15304 13326 15332 14282
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15304 12850 15332 13262
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15200 12708 15252 12714
rect 15200 12650 15252 12656
rect 15212 12238 15240 12650
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 15108 12164 15160 12170
rect 15108 12106 15160 12112
rect 15120 11354 15148 12106
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 15212 11830 15240 12038
rect 15200 11824 15252 11830
rect 15200 11766 15252 11772
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15212 10606 15240 11154
rect 15396 10674 15424 12922
rect 15488 11762 15516 18090
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15580 13802 15608 14350
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15672 13190 15700 14554
rect 15764 14550 15792 18022
rect 15856 15978 15884 18822
rect 15948 18766 15976 19110
rect 15936 18760 15988 18766
rect 15936 18702 15988 18708
rect 16040 18426 16068 25774
rect 16120 24608 16172 24614
rect 16120 24550 16172 24556
rect 16132 23730 16160 24550
rect 16120 23724 16172 23730
rect 16120 23666 16172 23672
rect 16120 20800 16172 20806
rect 16120 20742 16172 20748
rect 16028 18420 16080 18426
rect 16028 18362 16080 18368
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 15844 15972 15896 15978
rect 15844 15914 15896 15920
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 15856 14618 15884 14962
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 15948 14550 15976 18226
rect 16132 16114 16160 20742
rect 16224 19496 16252 26182
rect 16316 25294 16344 26318
rect 16868 26314 16896 26415
rect 16960 26353 16988 26930
rect 17144 26874 17172 29582
rect 17236 27033 17264 31214
rect 17408 30932 17460 30938
rect 17408 30874 17460 30880
rect 17420 27962 17448 30874
rect 17512 28150 17540 31282
rect 17868 31272 17920 31278
rect 17868 31214 17920 31220
rect 17880 30938 17908 31214
rect 17868 30932 17920 30938
rect 17868 30874 17920 30880
rect 17684 30660 17736 30666
rect 17684 30602 17736 30608
rect 17696 30190 17724 30602
rect 17776 30592 17828 30598
rect 17776 30534 17828 30540
rect 17684 30184 17736 30190
rect 17684 30126 17736 30132
rect 17592 29164 17644 29170
rect 17592 29106 17644 29112
rect 17604 28694 17632 29106
rect 17592 28688 17644 28694
rect 17592 28630 17644 28636
rect 17696 28540 17724 30126
rect 17788 29209 17816 30534
rect 17774 29200 17830 29209
rect 17774 29135 17830 29144
rect 17868 29164 17920 29170
rect 17604 28512 17724 28540
rect 17500 28144 17552 28150
rect 17500 28086 17552 28092
rect 17420 27934 17540 27962
rect 17316 27872 17368 27878
rect 17316 27814 17368 27820
rect 17408 27872 17460 27878
rect 17408 27814 17460 27820
rect 17222 27024 17278 27033
rect 17328 26994 17356 27814
rect 17420 27470 17448 27814
rect 17408 27464 17460 27470
rect 17408 27406 17460 27412
rect 17222 26959 17224 26968
rect 17276 26959 17278 26968
rect 17316 26988 17368 26994
rect 17224 26930 17276 26936
rect 17316 26930 17368 26936
rect 17052 26846 17172 26874
rect 16946 26344 17002 26353
rect 16856 26308 16908 26314
rect 16946 26279 17002 26288
rect 16856 26250 16908 26256
rect 16764 26240 16816 26246
rect 16764 26182 16816 26188
rect 16776 26042 16804 26182
rect 16764 26036 16816 26042
rect 16764 25978 16816 25984
rect 16856 25696 16908 25702
rect 16856 25638 16908 25644
rect 16304 25288 16356 25294
rect 16304 25230 16356 25236
rect 16396 25288 16448 25294
rect 16396 25230 16448 25236
rect 16304 25152 16356 25158
rect 16304 25094 16356 25100
rect 16316 24818 16344 25094
rect 16304 24812 16356 24818
rect 16304 24754 16356 24760
rect 16316 24274 16344 24754
rect 16304 24268 16356 24274
rect 16304 24210 16356 24216
rect 16408 24206 16436 25230
rect 16396 24200 16448 24206
rect 16396 24142 16448 24148
rect 16764 23724 16816 23730
rect 16764 23666 16816 23672
rect 16580 23588 16632 23594
rect 16580 23530 16632 23536
rect 16592 23322 16620 23530
rect 16580 23316 16632 23322
rect 16580 23258 16632 23264
rect 16672 23316 16724 23322
rect 16672 23258 16724 23264
rect 16488 22432 16540 22438
rect 16488 22374 16540 22380
rect 16302 20496 16358 20505
rect 16302 20431 16304 20440
rect 16356 20431 16358 20440
rect 16396 20460 16448 20466
rect 16304 20402 16356 20408
rect 16396 20402 16448 20408
rect 16224 19468 16344 19496
rect 16212 19372 16264 19378
rect 16212 19314 16264 19320
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16120 15972 16172 15978
rect 16120 15914 16172 15920
rect 16028 14612 16080 14618
rect 16028 14554 16080 14560
rect 15752 14544 15804 14550
rect 15752 14486 15804 14492
rect 15936 14544 15988 14550
rect 15936 14486 15988 14492
rect 15948 14414 15976 14486
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 16040 13530 16068 14554
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 15660 13184 15712 13190
rect 15660 13126 15712 13132
rect 16132 11762 16160 15914
rect 16224 14006 16252 19314
rect 16316 19258 16344 19468
rect 16408 19378 16436 20402
rect 16396 19372 16448 19378
rect 16396 19314 16448 19320
rect 16316 19230 16436 19258
rect 16304 18352 16356 18358
rect 16304 18294 16356 18300
rect 16212 14000 16264 14006
rect 16212 13942 16264 13948
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15200 10600 15252 10606
rect 15028 10526 15148 10554
rect 15200 10542 15252 10548
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 14372 9580 14424 9586
rect 14372 9522 14424 9528
rect 14476 9382 14504 9658
rect 14568 9518 14596 10202
rect 15028 10062 15056 10406
rect 15016 10056 15068 10062
rect 15016 9998 15068 10004
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14372 8560 14424 8566
rect 14372 8502 14424 8508
rect 14094 7984 14150 7993
rect 14094 7919 14150 7928
rect 14108 7886 14136 7919
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 13004 7002 13032 7278
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12992 6996 13044 7002
rect 12992 6938 13044 6944
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 11888 4208 11940 4214
rect 11888 4150 11940 4156
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11624 3058 11652 3674
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 11808 2514 11836 2926
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 11336 2440 11388 2446
rect 11336 2382 11388 2388
rect 11900 2378 11928 3878
rect 12268 3738 12296 4558
rect 12728 4282 12756 6938
rect 13832 6866 13860 7686
rect 14016 7342 14044 7822
rect 14108 7528 14136 7822
rect 14280 7540 14332 7546
rect 14108 7500 14280 7528
rect 14280 7482 14332 7488
rect 14384 7478 14412 8502
rect 14568 8412 14596 9454
rect 14660 8974 14688 9862
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 14740 8560 14792 8566
rect 14844 8548 14872 9862
rect 15028 9722 15056 9998
rect 15016 9716 15068 9722
rect 15016 9658 15068 9664
rect 15028 9450 15056 9658
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 14792 8520 14872 8548
rect 14740 8502 14792 8508
rect 14740 8424 14792 8430
rect 14568 8384 14740 8412
rect 15120 8378 15148 10526
rect 15384 9988 15436 9994
rect 15384 9930 15436 9936
rect 15396 9722 15424 9930
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15396 8838 15424 9522
rect 15488 9042 15516 11698
rect 16132 11218 16160 11698
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 16316 9674 16344 18294
rect 16408 16794 16436 19230
rect 16396 16788 16448 16794
rect 16396 16730 16448 16736
rect 16500 16182 16528 22374
rect 16580 22024 16632 22030
rect 16580 21966 16632 21972
rect 16592 21486 16620 21966
rect 16580 21480 16632 21486
rect 16580 21422 16632 21428
rect 16592 20398 16620 21422
rect 16580 20392 16632 20398
rect 16580 20334 16632 20340
rect 16580 18148 16632 18154
rect 16580 18090 16632 18096
rect 16592 17882 16620 18090
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16684 17218 16712 23258
rect 16776 19310 16804 23666
rect 16868 20806 16896 25638
rect 17052 24138 17080 26846
rect 17132 26308 17184 26314
rect 17132 26250 17184 26256
rect 17144 25265 17172 26250
rect 17316 26240 17368 26246
rect 17314 26208 17316 26217
rect 17368 26208 17370 26217
rect 17314 26143 17370 26152
rect 17408 25424 17460 25430
rect 17408 25366 17460 25372
rect 17130 25256 17186 25265
rect 17130 25191 17186 25200
rect 17316 25220 17368 25226
rect 17316 25162 17368 25168
rect 17132 25152 17184 25158
rect 17132 25094 17184 25100
rect 17144 24954 17172 25094
rect 17132 24948 17184 24954
rect 17132 24890 17184 24896
rect 17144 24818 17172 24890
rect 17328 24818 17356 25162
rect 17420 24818 17448 25366
rect 17132 24812 17184 24818
rect 17132 24754 17184 24760
rect 17316 24812 17368 24818
rect 17316 24754 17368 24760
rect 17408 24812 17460 24818
rect 17408 24754 17460 24760
rect 17328 24410 17356 24754
rect 17316 24404 17368 24410
rect 17316 24346 17368 24352
rect 17040 24132 17092 24138
rect 17040 24074 17092 24080
rect 17052 23662 17080 24074
rect 17040 23656 17092 23662
rect 17040 23598 17092 23604
rect 17408 23656 17460 23662
rect 17408 23598 17460 23604
rect 16948 23112 17000 23118
rect 16948 23054 17000 23060
rect 16960 22506 16988 23054
rect 16948 22500 17000 22506
rect 16948 22442 17000 22448
rect 16960 22030 16988 22442
rect 16948 22024 17000 22030
rect 16948 21966 17000 21972
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17144 21690 17172 21966
rect 17420 21962 17448 23598
rect 17408 21956 17460 21962
rect 17408 21898 17460 21904
rect 17224 21888 17276 21894
rect 17224 21830 17276 21836
rect 17132 21684 17184 21690
rect 17132 21626 17184 21632
rect 17040 21480 17092 21486
rect 17040 21422 17092 21428
rect 17052 20942 17080 21422
rect 17132 21072 17184 21078
rect 17132 21014 17184 21020
rect 17040 20936 17092 20942
rect 17040 20878 17092 20884
rect 16856 20800 16908 20806
rect 16856 20742 16908 20748
rect 17144 20534 17172 21014
rect 17132 20528 17184 20534
rect 17132 20470 17184 20476
rect 17040 19984 17092 19990
rect 17040 19926 17092 19932
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16776 18426 16804 19246
rect 16856 19236 16908 19242
rect 16856 19178 16908 19184
rect 16764 18420 16816 18426
rect 16764 18362 16816 18368
rect 16592 17190 16712 17218
rect 16868 17202 16896 19178
rect 17052 17882 17080 19926
rect 17144 19514 17172 20470
rect 17132 19508 17184 19514
rect 17132 19450 17184 19456
rect 17040 17876 17092 17882
rect 17040 17818 17092 17824
rect 16946 17776 17002 17785
rect 16946 17711 17002 17720
rect 17052 17728 17080 17818
rect 16960 17678 16988 17711
rect 17052 17700 17172 17728
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 16856 17196 16908 17202
rect 16488 16176 16540 16182
rect 16488 16118 16540 16124
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16408 15706 16436 16050
rect 16396 15700 16448 15706
rect 16396 15642 16448 15648
rect 16500 15026 16528 16118
rect 16488 15020 16540 15026
rect 16488 14962 16540 14968
rect 16500 14822 16528 14962
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16592 11150 16620 17190
rect 16856 17138 16908 17144
rect 16960 17082 16988 17614
rect 17040 17604 17092 17610
rect 17040 17546 17092 17552
rect 17052 17202 17080 17546
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 16776 17054 16988 17082
rect 16672 16448 16724 16454
rect 16672 16390 16724 16396
rect 16684 15586 16712 16390
rect 16776 15706 16804 17054
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16764 15700 16816 15706
rect 16764 15642 16816 15648
rect 16684 15558 16804 15586
rect 16776 15502 16804 15558
rect 16960 15502 16988 16934
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16764 15496 16816 15502
rect 16764 15438 16816 15444
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16684 14074 16712 15438
rect 16764 15088 16816 15094
rect 17052 15042 17080 15642
rect 16764 15030 16816 15036
rect 16776 14414 16804 15030
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16960 15014 17080 15042
rect 16868 14482 16896 14962
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16764 14408 16816 14414
rect 16816 14356 16896 14362
rect 16764 14350 16896 14356
rect 16776 14334 16896 14350
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16776 14074 16804 14214
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 16684 13530 16712 14010
rect 16868 13682 16896 14334
rect 16776 13654 16896 13682
rect 16672 13524 16724 13530
rect 16672 13466 16724 13472
rect 16776 13326 16804 13654
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16684 12918 16712 13262
rect 16672 12912 16724 12918
rect 16672 12854 16724 12860
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16224 9646 16344 9674
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15856 9382 15884 9522
rect 15948 9450 15976 9522
rect 15936 9444 15988 9450
rect 15936 9386 15988 9392
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15488 8786 15516 8978
rect 15488 8758 15792 8786
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 14740 8366 14792 8372
rect 15028 8350 15148 8378
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14568 7546 14596 7686
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 14372 7472 14424 7478
rect 14372 7414 14424 7420
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14200 6934 14228 7142
rect 14384 6934 14412 7414
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14188 6928 14240 6934
rect 14188 6870 14240 6876
rect 14372 6928 14424 6934
rect 14372 6870 14424 6876
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 12912 3534 12940 6802
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13648 6458 13676 6734
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 12992 6180 13044 6186
rect 12992 6122 13044 6128
rect 13004 4690 13032 6122
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13360 5296 13412 5302
rect 13360 5238 13412 5244
rect 12992 4684 13044 4690
rect 12992 4626 13044 4632
rect 13004 4078 13032 4626
rect 12992 4072 13044 4078
rect 13044 4032 13124 4060
rect 12992 4014 13044 4020
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13004 3602 13032 3878
rect 13096 3602 13124 4032
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12544 3126 12572 3334
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 13372 3058 13400 5238
rect 13832 4622 13860 5306
rect 13912 4752 13964 4758
rect 13912 4694 13964 4700
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13924 4185 13952 4694
rect 14200 4554 14228 6870
rect 14568 6798 14596 7142
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14292 4826 14320 5102
rect 14280 4820 14332 4826
rect 14280 4762 14332 4768
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14188 4548 14240 4554
rect 14188 4490 14240 4496
rect 13910 4176 13966 4185
rect 13910 4111 13966 4120
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 12348 2848 12400 2854
rect 12348 2790 12400 2796
rect 11888 2372 11940 2378
rect 11888 2314 11940 2320
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 11624 800 11652 2246
rect 12360 1442 12388 2790
rect 12820 2378 12848 2926
rect 13832 2922 13860 4014
rect 13924 3534 13952 4111
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 13820 2916 13872 2922
rect 13820 2858 13872 2864
rect 12900 2576 12952 2582
rect 12900 2518 12952 2524
rect 13544 2576 13596 2582
rect 13544 2518 13596 2524
rect 12808 2372 12860 2378
rect 12808 2314 12860 2320
rect 12268 1414 12388 1442
rect 12268 800 12296 1414
rect 12912 800 12940 2518
rect 13556 800 13584 2518
rect 13832 2378 13860 2858
rect 14016 2446 14044 4014
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 14108 3126 14136 3334
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 14292 2446 14320 4558
rect 14660 3534 14688 7278
rect 14752 7206 14780 7822
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 15028 6662 15056 8350
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 15120 8022 15148 8230
rect 15212 8090 15240 8434
rect 15304 8090 15332 8434
rect 15384 8424 15436 8430
rect 15488 8412 15516 8758
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15436 8384 15516 8412
rect 15384 8366 15436 8372
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 15108 8016 15160 8022
rect 15396 7970 15424 8366
rect 15580 8129 15608 8570
rect 15658 8528 15714 8537
rect 15658 8463 15660 8472
rect 15712 8463 15714 8472
rect 15660 8434 15712 8440
rect 15566 8120 15622 8129
rect 15566 8055 15622 8064
rect 15580 8022 15608 8055
rect 15108 7958 15160 7964
rect 15212 7942 15424 7970
rect 15568 8016 15620 8022
rect 15568 7958 15620 7964
rect 15108 6860 15160 6866
rect 15108 6802 15160 6808
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 15120 6458 15148 6802
rect 15108 6452 15160 6458
rect 15108 6394 15160 6400
rect 15212 6390 15240 7942
rect 15292 7880 15344 7886
rect 15672 7834 15700 8434
rect 15764 7954 15792 8758
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15856 7886 15884 8230
rect 15344 7828 15700 7834
rect 15292 7822 15700 7828
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15936 7880 15988 7886
rect 15936 7822 15988 7828
rect 15304 7806 15700 7822
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15304 7410 15332 7686
rect 15948 7546 15976 7822
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15304 6798 15332 7346
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15384 6928 15436 6934
rect 15384 6870 15436 6876
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15396 6390 15424 6870
rect 15580 6866 15608 7142
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15948 6730 15976 7278
rect 15936 6724 15988 6730
rect 15936 6666 15988 6672
rect 15200 6384 15252 6390
rect 15200 6326 15252 6332
rect 15384 6384 15436 6390
rect 15384 6326 15436 6332
rect 14924 5092 14976 5098
rect 14924 5034 14976 5040
rect 14936 4758 14964 5034
rect 15212 5030 15240 6326
rect 15396 5302 15424 6326
rect 15948 6186 15976 6666
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 16224 6118 16252 9646
rect 16486 9616 16542 9625
rect 16486 9551 16542 9560
rect 16500 8974 16528 9551
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16316 7410 16344 7890
rect 16500 7478 16528 8910
rect 16684 8090 16712 12582
rect 16868 11898 16896 13466
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16960 11778 16988 15014
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 17052 13530 17080 14894
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 17144 13258 17172 17700
rect 17236 16590 17264 21830
rect 17420 21418 17448 21898
rect 17408 21412 17460 21418
rect 17408 21354 17460 21360
rect 17316 21344 17368 21350
rect 17316 21286 17368 21292
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17328 14414 17356 21286
rect 17420 20806 17448 21354
rect 17408 20800 17460 20806
rect 17512 20777 17540 27934
rect 17408 20742 17460 20748
rect 17498 20768 17554 20777
rect 17498 20703 17554 20712
rect 17604 20398 17632 28512
rect 17684 28076 17736 28082
rect 17684 28018 17736 28024
rect 17696 27674 17724 28018
rect 17684 27668 17736 27674
rect 17684 27610 17736 27616
rect 17788 27554 17816 29135
rect 17868 29106 17920 29112
rect 17880 28626 17908 29106
rect 17868 28620 17920 28626
rect 17868 28562 17920 28568
rect 17868 27872 17920 27878
rect 17868 27814 17920 27820
rect 17880 27674 17908 27814
rect 17868 27668 17920 27674
rect 17868 27610 17920 27616
rect 17788 27526 17908 27554
rect 17776 27396 17828 27402
rect 17776 27338 17828 27344
rect 17788 26994 17816 27338
rect 17776 26988 17828 26994
rect 17776 26930 17828 26936
rect 17684 25832 17736 25838
rect 17684 25774 17736 25780
rect 17696 24886 17724 25774
rect 17684 24880 17736 24886
rect 17684 24822 17736 24828
rect 17788 24188 17816 26930
rect 17880 26314 17908 27526
rect 17868 26308 17920 26314
rect 17868 26250 17920 26256
rect 17880 25498 17908 26250
rect 17972 26234 18000 31690
rect 18064 31482 18092 31826
rect 18524 31686 18552 33390
rect 18616 32842 18644 33594
rect 18604 32836 18656 32842
rect 18604 32778 18656 32784
rect 18512 31680 18564 31686
rect 18512 31622 18564 31628
rect 19064 31680 19116 31686
rect 19064 31622 19116 31628
rect 18052 31476 18104 31482
rect 18052 31418 18104 31424
rect 18236 31340 18288 31346
rect 18236 31282 18288 31288
rect 18420 31340 18472 31346
rect 18420 31282 18472 31288
rect 18248 30394 18276 31282
rect 18432 30938 18460 31282
rect 19076 31278 19104 31622
rect 19168 31414 19196 34564
rect 19248 34546 19300 34552
rect 19248 34468 19300 34474
rect 19248 34410 19300 34416
rect 19260 33590 19288 34410
rect 19248 33584 19300 33590
rect 19248 33526 19300 33532
rect 19432 32360 19484 32366
rect 19432 32302 19484 32308
rect 19248 31748 19300 31754
rect 19248 31690 19300 31696
rect 19260 31414 19288 31690
rect 19156 31408 19208 31414
rect 19156 31350 19208 31356
rect 19248 31408 19300 31414
rect 19248 31350 19300 31356
rect 19064 31272 19116 31278
rect 19064 31214 19116 31220
rect 18420 30932 18472 30938
rect 18420 30874 18472 30880
rect 18696 30932 18748 30938
rect 18696 30874 18748 30880
rect 18328 30728 18380 30734
rect 18328 30670 18380 30676
rect 18236 30388 18288 30394
rect 18236 30330 18288 30336
rect 18340 30138 18368 30670
rect 18432 30258 18460 30874
rect 18604 30660 18656 30666
rect 18604 30602 18656 30608
rect 18420 30252 18472 30258
rect 18420 30194 18472 30200
rect 18616 30190 18644 30602
rect 18604 30184 18656 30190
rect 18340 30110 18460 30138
rect 18604 30126 18656 30132
rect 18326 30016 18382 30025
rect 18326 29951 18382 29960
rect 18340 29850 18368 29951
rect 18328 29844 18380 29850
rect 18328 29786 18380 29792
rect 18144 28008 18196 28014
rect 18144 27950 18196 27956
rect 18052 27328 18104 27334
rect 18052 27270 18104 27276
rect 18064 26926 18092 27270
rect 18052 26920 18104 26926
rect 18052 26862 18104 26868
rect 18064 26382 18092 26862
rect 18156 26382 18184 27950
rect 18236 27396 18288 27402
rect 18236 27338 18288 27344
rect 18248 27282 18276 27338
rect 18248 27254 18368 27282
rect 18340 26994 18368 27254
rect 18328 26988 18380 26994
rect 18328 26930 18380 26936
rect 18340 26586 18368 26930
rect 18328 26580 18380 26586
rect 18328 26522 18380 26528
rect 18052 26376 18104 26382
rect 18052 26318 18104 26324
rect 18144 26376 18196 26382
rect 18144 26318 18196 26324
rect 18236 26376 18288 26382
rect 18236 26318 18288 26324
rect 17972 26206 18092 26234
rect 17868 25492 17920 25498
rect 17868 25434 17920 25440
rect 17960 24200 18012 24206
rect 17788 24160 17960 24188
rect 17960 24142 18012 24148
rect 17972 23730 18000 24142
rect 18064 23798 18092 26206
rect 18248 25906 18276 26318
rect 18236 25900 18288 25906
rect 18236 25842 18288 25848
rect 18328 25900 18380 25906
rect 18328 25842 18380 25848
rect 18144 25764 18196 25770
rect 18144 25706 18196 25712
rect 18156 25158 18184 25706
rect 18248 25412 18276 25842
rect 18340 25537 18368 25842
rect 18326 25528 18382 25537
rect 18326 25463 18382 25472
rect 18248 25384 18368 25412
rect 18144 25152 18196 25158
rect 18144 25094 18196 25100
rect 18052 23792 18104 23798
rect 18052 23734 18104 23740
rect 17960 23724 18012 23730
rect 17960 23666 18012 23672
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 18064 23322 18092 23598
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 18050 23080 18106 23089
rect 18050 23015 18106 23024
rect 18064 22982 18092 23015
rect 17684 22976 17736 22982
rect 17684 22918 17736 22924
rect 17960 22976 18012 22982
rect 17960 22918 18012 22924
rect 18052 22976 18104 22982
rect 18052 22918 18104 22924
rect 17696 22098 17724 22918
rect 17684 22092 17736 22098
rect 17684 22034 17736 22040
rect 17684 21888 17736 21894
rect 17684 21830 17736 21836
rect 17868 21888 17920 21894
rect 17868 21830 17920 21836
rect 17592 20392 17644 20398
rect 17592 20334 17644 20340
rect 17592 19780 17644 19786
rect 17592 19722 17644 19728
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 17420 19514 17448 19654
rect 17408 19508 17460 19514
rect 17460 19468 17540 19496
rect 17408 19450 17460 19456
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 17420 16726 17448 17274
rect 17408 16720 17460 16726
rect 17408 16662 17460 16668
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 17420 15706 17448 15982
rect 17408 15700 17460 15706
rect 17408 15642 17460 15648
rect 17512 15094 17540 19468
rect 17604 19378 17632 19722
rect 17592 19372 17644 19378
rect 17592 19314 17644 19320
rect 17592 15564 17644 15570
rect 17592 15506 17644 15512
rect 17500 15088 17552 15094
rect 17500 15030 17552 15036
rect 17604 14482 17632 15506
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17224 14000 17276 14006
rect 17224 13942 17276 13948
rect 17236 13530 17264 13942
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 17420 13326 17448 14214
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17408 13320 17460 13326
rect 17604 13308 17632 14418
rect 17696 13818 17724 21830
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 17788 19378 17816 21626
rect 17880 21554 17908 21830
rect 17972 21593 18000 22918
rect 18052 22772 18104 22778
rect 18052 22714 18104 22720
rect 17958 21584 18014 21593
rect 17868 21548 17920 21554
rect 17958 21519 18014 21528
rect 17868 21490 17920 21496
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17788 17270 17816 19314
rect 17776 17264 17828 17270
rect 17776 17206 17828 17212
rect 17776 15428 17828 15434
rect 17776 15370 17828 15376
rect 17788 14822 17816 15370
rect 17880 15094 17908 21490
rect 17972 19258 18000 21519
rect 18064 19446 18092 22714
rect 18052 19440 18104 19446
rect 18052 19382 18104 19388
rect 17972 19230 18092 19258
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17972 15502 18000 18566
rect 18064 17882 18092 19230
rect 18156 18222 18184 25094
rect 18236 23112 18288 23118
rect 18236 23054 18288 23060
rect 18248 22778 18276 23054
rect 18236 22772 18288 22778
rect 18236 22714 18288 22720
rect 18236 22228 18288 22234
rect 18236 22170 18288 22176
rect 18248 22030 18276 22170
rect 18340 22098 18368 25384
rect 18432 24750 18460 30110
rect 18512 29844 18564 29850
rect 18512 29786 18564 29792
rect 18524 29646 18552 29786
rect 18512 29640 18564 29646
rect 18616 29617 18644 30126
rect 18708 30122 18736 30874
rect 18696 30116 18748 30122
rect 18696 30058 18748 30064
rect 18788 29640 18840 29646
rect 18512 29582 18564 29588
rect 18602 29608 18658 29617
rect 18788 29582 18840 29588
rect 18880 29640 18932 29646
rect 18880 29582 18932 29588
rect 18972 29640 19024 29646
rect 18972 29582 19024 29588
rect 18602 29543 18658 29552
rect 18800 29238 18828 29582
rect 18788 29232 18840 29238
rect 18788 29174 18840 29180
rect 18604 29028 18656 29034
rect 18604 28970 18656 28976
rect 18510 27568 18566 27577
rect 18510 27503 18566 27512
rect 18524 27470 18552 27503
rect 18512 27464 18564 27470
rect 18512 27406 18564 27412
rect 18616 26858 18644 28970
rect 18696 28008 18748 28014
rect 18696 27950 18748 27956
rect 18708 27470 18736 27950
rect 18696 27464 18748 27470
rect 18696 27406 18748 27412
rect 18788 27464 18840 27470
rect 18788 27406 18840 27412
rect 18708 27062 18736 27406
rect 18696 27056 18748 27062
rect 18696 26998 18748 27004
rect 18800 26926 18828 27406
rect 18696 26920 18748 26926
rect 18696 26862 18748 26868
rect 18788 26920 18840 26926
rect 18788 26862 18840 26868
rect 18604 26852 18656 26858
rect 18604 26794 18656 26800
rect 18708 26586 18736 26862
rect 18696 26580 18748 26586
rect 18696 26522 18748 26528
rect 18696 26240 18748 26246
rect 18696 26182 18748 26188
rect 18604 25220 18656 25226
rect 18604 25162 18656 25168
rect 18616 24954 18644 25162
rect 18604 24948 18656 24954
rect 18604 24890 18656 24896
rect 18512 24812 18564 24818
rect 18512 24754 18564 24760
rect 18420 24744 18472 24750
rect 18420 24686 18472 24692
rect 18524 24138 18552 24754
rect 18604 24268 18656 24274
rect 18604 24210 18656 24216
rect 18420 24132 18472 24138
rect 18420 24074 18472 24080
rect 18512 24132 18564 24138
rect 18512 24074 18564 24080
rect 18432 23866 18460 24074
rect 18420 23860 18472 23866
rect 18420 23802 18472 23808
rect 18420 23656 18472 23662
rect 18418 23624 18420 23633
rect 18472 23624 18474 23633
rect 18418 23559 18474 23568
rect 18420 23112 18472 23118
rect 18524 23100 18552 24074
rect 18472 23072 18552 23100
rect 18420 23054 18472 23060
rect 18328 22092 18380 22098
rect 18432 22094 18460 23054
rect 18616 22778 18644 24210
rect 18708 23322 18736 26182
rect 18892 26042 18920 29582
rect 18984 29102 19012 29582
rect 18972 29096 19024 29102
rect 18972 29038 19024 29044
rect 18970 27568 19026 27577
rect 18970 27503 19026 27512
rect 18984 27470 19012 27503
rect 18972 27464 19024 27470
rect 18972 27406 19024 27412
rect 18880 26036 18932 26042
rect 18880 25978 18932 25984
rect 19076 25906 19104 31214
rect 19444 30666 19472 32302
rect 19536 31142 19564 35634
rect 19628 34542 19656 36110
rect 19720 35222 19748 37198
rect 19904 37194 19932 38490
rect 20088 38010 20116 38830
rect 20628 38480 20680 38486
rect 20628 38422 20680 38428
rect 20076 38004 20128 38010
rect 20076 37946 20128 37952
rect 20640 37942 20668 38422
rect 20628 37936 20680 37942
rect 20628 37878 20680 37884
rect 19892 37188 19944 37194
rect 19892 37130 19944 37136
rect 20640 36650 20668 37878
rect 20732 36854 20760 39034
rect 20812 39024 20864 39030
rect 20812 38966 20864 38972
rect 23204 39024 23256 39030
rect 23204 38966 23256 38972
rect 20824 38486 20852 38966
rect 23020 38888 23072 38894
rect 23020 38830 23072 38836
rect 20812 38480 20864 38486
rect 20812 38422 20864 38428
rect 21272 38480 21324 38486
rect 21272 38422 21324 38428
rect 21180 38344 21232 38350
rect 21180 38286 21232 38292
rect 20720 36848 20772 36854
rect 20720 36790 20772 36796
rect 20628 36644 20680 36650
rect 20628 36586 20680 36592
rect 20640 36106 20668 36586
rect 19892 36100 19944 36106
rect 19892 36042 19944 36048
rect 20628 36100 20680 36106
rect 20628 36042 20680 36048
rect 19904 35834 19932 36042
rect 19892 35828 19944 35834
rect 19892 35770 19944 35776
rect 19800 35692 19852 35698
rect 19800 35634 19852 35640
rect 19708 35216 19760 35222
rect 19708 35158 19760 35164
rect 19708 34944 19760 34950
rect 19812 34932 19840 35634
rect 19892 35080 19944 35086
rect 20536 35080 20588 35086
rect 19892 35022 19944 35028
rect 20534 35048 20536 35057
rect 20588 35048 20590 35057
rect 19760 34904 19840 34932
rect 19708 34886 19760 34892
rect 19616 34536 19668 34542
rect 19616 34478 19668 34484
rect 19720 33454 19748 34886
rect 19708 33448 19760 33454
rect 19708 33390 19760 33396
rect 19904 33318 19932 35022
rect 20534 34983 20590 34992
rect 20168 34060 20220 34066
rect 20168 34002 20220 34008
rect 20180 33658 20208 34002
rect 20168 33652 20220 33658
rect 20168 33594 20220 33600
rect 19892 33312 19944 33318
rect 19892 33254 19944 33260
rect 20352 32496 20404 32502
rect 20352 32438 20404 32444
rect 20364 32366 20392 32438
rect 20352 32360 20404 32366
rect 20352 32302 20404 32308
rect 20352 32224 20404 32230
rect 20352 32166 20404 32172
rect 19616 31748 19668 31754
rect 19616 31690 19668 31696
rect 19628 31482 19656 31690
rect 19616 31476 19668 31482
rect 19616 31418 19668 31424
rect 20364 31278 20392 32166
rect 20640 31890 20668 36042
rect 20812 35284 20864 35290
rect 20812 35226 20864 35232
rect 20824 35068 20852 35226
rect 20996 35080 21048 35086
rect 20824 35040 20996 35068
rect 21048 35040 21128 35068
rect 20996 35022 21048 35028
rect 20904 34944 20956 34950
rect 20904 34886 20956 34892
rect 20916 34066 20944 34886
rect 21100 34542 21128 35040
rect 21192 34950 21220 38286
rect 21284 37262 21312 38422
rect 23032 38350 23060 38830
rect 23216 38554 23244 38966
rect 23204 38548 23256 38554
rect 23204 38490 23256 38496
rect 22100 38344 22152 38350
rect 22100 38286 22152 38292
rect 23020 38344 23072 38350
rect 23020 38286 23072 38292
rect 21456 38208 21508 38214
rect 21456 38150 21508 38156
rect 21640 38208 21692 38214
rect 21640 38150 21692 38156
rect 21468 37670 21496 38150
rect 21548 37868 21600 37874
rect 21548 37810 21600 37816
rect 21456 37664 21508 37670
rect 21456 37606 21508 37612
rect 21468 37262 21496 37606
rect 21560 37398 21588 37810
rect 21548 37392 21600 37398
rect 21548 37334 21600 37340
rect 21652 37330 21680 38150
rect 22112 37874 22140 38286
rect 22376 38004 22428 38010
rect 22376 37946 22428 37952
rect 22100 37868 22152 37874
rect 22100 37810 22152 37816
rect 21824 37800 21876 37806
rect 21824 37742 21876 37748
rect 21836 37466 21864 37742
rect 21916 37664 21968 37670
rect 21916 37606 21968 37612
rect 21824 37460 21876 37466
rect 21824 37402 21876 37408
rect 21640 37324 21692 37330
rect 21640 37266 21692 37272
rect 21272 37256 21324 37262
rect 21272 37198 21324 37204
rect 21456 37256 21508 37262
rect 21456 37198 21508 37204
rect 21928 36174 21956 37606
rect 22112 37398 22140 37810
rect 22388 37806 22416 37946
rect 22376 37800 22428 37806
rect 22376 37742 22428 37748
rect 22652 37800 22704 37806
rect 22652 37742 22704 37748
rect 22664 37466 22692 37742
rect 23032 37670 23060 38286
rect 23860 37806 23888 43101
rect 24504 39030 24532 43101
rect 24492 39024 24544 39030
rect 24492 38966 24544 38972
rect 24504 38282 24532 38966
rect 24492 38276 24544 38282
rect 24492 38218 24544 38224
rect 24952 38276 25004 38282
rect 24952 38218 25004 38224
rect 24964 38010 24992 38218
rect 24952 38004 25004 38010
rect 24952 37946 25004 37952
rect 23848 37800 23900 37806
rect 23848 37742 23900 37748
rect 23020 37664 23072 37670
rect 23020 37606 23072 37612
rect 22652 37460 22704 37466
rect 22652 37402 22704 37408
rect 22100 37392 22152 37398
rect 22100 37334 22152 37340
rect 22560 37188 22612 37194
rect 22560 37130 22612 37136
rect 21916 36168 21968 36174
rect 21916 36110 21968 36116
rect 22284 36168 22336 36174
rect 22284 36110 22336 36116
rect 22468 36168 22520 36174
rect 22468 36110 22520 36116
rect 21364 36032 21416 36038
rect 21364 35974 21416 35980
rect 21376 35766 21404 35974
rect 21928 35766 21956 36110
rect 21364 35760 21416 35766
rect 21364 35702 21416 35708
rect 21916 35760 21968 35766
rect 21916 35702 21968 35708
rect 22006 35728 22062 35737
rect 21272 35624 21324 35630
rect 21272 35566 21324 35572
rect 21284 35154 21312 35566
rect 21376 35465 21404 35702
rect 22006 35663 22008 35672
rect 22060 35663 22062 35672
rect 22008 35634 22060 35640
rect 21640 35556 21692 35562
rect 21640 35498 21692 35504
rect 21456 35488 21508 35494
rect 21362 35456 21418 35465
rect 21456 35430 21508 35436
rect 21362 35391 21418 35400
rect 21272 35148 21324 35154
rect 21272 35090 21324 35096
rect 21468 35057 21496 35430
rect 21652 35222 21680 35498
rect 21640 35216 21692 35222
rect 21640 35158 21692 35164
rect 21454 35048 21510 35057
rect 21454 34983 21510 34992
rect 21180 34944 21232 34950
rect 21180 34886 21232 34892
rect 21180 34672 21232 34678
rect 21180 34614 21232 34620
rect 21088 34536 21140 34542
rect 21088 34478 21140 34484
rect 21192 34388 21220 34614
rect 21468 34610 21496 34983
rect 21548 34740 21600 34746
rect 21548 34682 21600 34688
rect 21456 34604 21508 34610
rect 21456 34546 21508 34552
rect 21100 34360 21220 34388
rect 20904 34060 20956 34066
rect 20904 34002 20956 34008
rect 20904 32428 20956 32434
rect 20904 32370 20956 32376
rect 20628 31884 20680 31890
rect 20628 31826 20680 31832
rect 20352 31272 20404 31278
rect 20352 31214 20404 31220
rect 20444 31272 20496 31278
rect 20444 31214 20496 31220
rect 19524 31136 19576 31142
rect 19524 31078 19576 31084
rect 20456 30802 20484 31214
rect 20916 31142 20944 32370
rect 21100 32026 21128 34360
rect 21560 34134 21588 34682
rect 21652 34678 21680 35158
rect 21732 35148 21784 35154
rect 21732 35090 21784 35096
rect 21640 34672 21692 34678
rect 21640 34614 21692 34620
rect 21744 34490 21772 35090
rect 21824 34536 21876 34542
rect 21744 34484 21824 34490
rect 21744 34478 21876 34484
rect 21744 34462 21864 34478
rect 21548 34128 21600 34134
rect 21548 34070 21600 34076
rect 21744 33930 21772 34462
rect 21824 34400 21876 34406
rect 21824 34342 21876 34348
rect 21836 33998 21864 34342
rect 21824 33992 21876 33998
rect 21824 33934 21876 33940
rect 21732 33924 21784 33930
rect 21732 33866 21784 33872
rect 21456 32496 21508 32502
rect 21456 32438 21508 32444
rect 21088 32020 21140 32026
rect 21088 31962 21140 31968
rect 20996 31340 21048 31346
rect 20996 31282 21048 31288
rect 20812 31136 20864 31142
rect 20812 31078 20864 31084
rect 20904 31136 20956 31142
rect 20904 31078 20956 31084
rect 20824 30802 20852 31078
rect 20444 30796 20496 30802
rect 20444 30738 20496 30744
rect 20812 30796 20864 30802
rect 20812 30738 20864 30744
rect 19432 30660 19484 30666
rect 19432 30602 19484 30608
rect 19156 29776 19208 29782
rect 19156 29718 19208 29724
rect 19168 28966 19196 29718
rect 19984 29708 20036 29714
rect 19984 29650 20036 29656
rect 19432 29572 19484 29578
rect 19432 29514 19484 29520
rect 19156 28960 19208 28966
rect 19156 28902 19208 28908
rect 19444 28150 19472 29514
rect 19524 29504 19576 29510
rect 19524 29446 19576 29452
rect 19536 29306 19564 29446
rect 19524 29300 19576 29306
rect 19524 29242 19576 29248
rect 19432 28144 19484 28150
rect 19432 28086 19484 28092
rect 19156 28008 19208 28014
rect 19156 27950 19208 27956
rect 19248 28008 19300 28014
rect 19248 27950 19300 27956
rect 19168 27878 19196 27950
rect 19156 27872 19208 27878
rect 19156 27814 19208 27820
rect 19168 26994 19196 27814
rect 19156 26988 19208 26994
rect 19156 26930 19208 26936
rect 19168 26586 19196 26930
rect 19260 26926 19288 27950
rect 19444 27402 19472 28086
rect 19708 28076 19760 28082
rect 19708 28018 19760 28024
rect 19616 28008 19668 28014
rect 19616 27950 19668 27956
rect 19524 27940 19576 27946
rect 19524 27882 19576 27888
rect 19432 27396 19484 27402
rect 19432 27338 19484 27344
rect 19444 27010 19472 27338
rect 19536 27282 19564 27882
rect 19628 27470 19656 27950
rect 19720 27470 19748 28018
rect 19892 27600 19944 27606
rect 19892 27542 19944 27548
rect 19616 27464 19668 27470
rect 19616 27406 19668 27412
rect 19708 27464 19760 27470
rect 19708 27406 19760 27412
rect 19904 27402 19932 27542
rect 19892 27396 19944 27402
rect 19892 27338 19944 27344
rect 19708 27328 19760 27334
rect 19536 27276 19708 27282
rect 19904 27282 19932 27338
rect 19536 27270 19760 27276
rect 19536 27254 19748 27270
rect 19720 27130 19748 27254
rect 19812 27254 19932 27282
rect 19708 27124 19760 27130
rect 19708 27066 19760 27072
rect 19444 26982 19748 27010
rect 19248 26920 19300 26926
rect 19248 26862 19300 26868
rect 19430 26888 19486 26897
rect 19430 26823 19486 26832
rect 19156 26580 19208 26586
rect 19156 26522 19208 26528
rect 19340 26376 19392 26382
rect 19340 26318 19392 26324
rect 19352 25974 19380 26318
rect 19340 25968 19392 25974
rect 19340 25910 19392 25916
rect 19064 25900 19116 25906
rect 19064 25842 19116 25848
rect 19076 25362 19104 25842
rect 19064 25356 19116 25362
rect 19064 25298 19116 25304
rect 19064 24812 19116 24818
rect 19064 24754 19116 24760
rect 18880 24744 18932 24750
rect 18880 24686 18932 24692
rect 18696 23316 18748 23322
rect 18696 23258 18748 23264
rect 18694 23216 18750 23225
rect 18694 23151 18696 23160
rect 18748 23151 18750 23160
rect 18696 23122 18748 23128
rect 18788 23112 18840 23118
rect 18788 23054 18840 23060
rect 18696 22976 18748 22982
rect 18696 22918 18748 22924
rect 18604 22772 18656 22778
rect 18604 22714 18656 22720
rect 18432 22066 18552 22094
rect 18328 22034 18380 22040
rect 18236 22024 18288 22030
rect 18236 21966 18288 21972
rect 18248 21486 18276 21966
rect 18236 21480 18288 21486
rect 18236 21422 18288 21428
rect 18420 21072 18472 21078
rect 18420 21014 18472 21020
rect 18236 20936 18288 20942
rect 18236 20878 18288 20884
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 18248 17678 18276 20878
rect 18328 20528 18380 20534
rect 18328 20470 18380 20476
rect 18340 19378 18368 20470
rect 18432 20262 18460 21014
rect 18524 20942 18552 22066
rect 18604 22092 18656 22098
rect 18604 22034 18656 22040
rect 18512 20936 18564 20942
rect 18512 20878 18564 20884
rect 18616 20874 18644 22034
rect 18604 20868 18656 20874
rect 18604 20810 18656 20816
rect 18420 20256 18472 20262
rect 18420 20198 18472 20204
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18236 17672 18288 17678
rect 18236 17614 18288 17620
rect 18052 17536 18104 17542
rect 18052 17478 18104 17484
rect 18064 16726 18092 17478
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18052 16720 18104 16726
rect 18052 16662 18104 16668
rect 18064 15502 18092 16662
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17868 15088 17920 15094
rect 17868 15030 17920 15036
rect 17972 14958 18000 15302
rect 18156 15094 18184 16526
rect 18248 15502 18276 17138
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 18144 15088 18196 15094
rect 18144 15030 18196 15036
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 17776 14816 17828 14822
rect 17776 14758 17828 14764
rect 17972 14618 18000 14894
rect 18248 14618 18276 15438
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17880 14006 17908 14214
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 17696 13790 18000 13818
rect 17972 13530 18000 13790
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 17960 13524 18012 13530
rect 18012 13484 18092 13512
rect 17960 13466 18012 13472
rect 17868 13320 17920 13326
rect 17604 13280 17868 13308
rect 17408 13262 17460 13268
rect 17868 13262 17920 13268
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 17132 13252 17184 13258
rect 17132 13194 17184 13200
rect 17144 12889 17172 13194
rect 17130 12880 17186 12889
rect 17130 12815 17186 12824
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 17052 12374 17080 12718
rect 17236 12646 17264 13262
rect 17316 12776 17368 12782
rect 17316 12718 17368 12724
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17328 12434 17356 12718
rect 17420 12714 17448 13262
rect 17500 13252 17552 13258
rect 17500 13194 17552 13200
rect 17512 12986 17540 13194
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17604 12986 17632 13126
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17592 12980 17644 12986
rect 17592 12922 17644 12928
rect 17590 12880 17646 12889
rect 17590 12815 17646 12824
rect 17684 12844 17736 12850
rect 17408 12708 17460 12714
rect 17408 12650 17460 12656
rect 17144 12406 17356 12434
rect 17040 12368 17092 12374
rect 17040 12310 17092 12316
rect 16960 11762 17080 11778
rect 16960 11756 17092 11762
rect 16960 11750 17040 11756
rect 17040 11698 17092 11704
rect 16764 11620 16816 11626
rect 16764 11562 16816 11568
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 16592 6866 16620 7278
rect 16684 7274 16712 8026
rect 16776 7818 16804 11562
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16960 10810 16988 11086
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 17052 10470 17080 11698
rect 17040 10464 17092 10470
rect 17040 10406 17092 10412
rect 16854 10296 16910 10305
rect 16854 10231 16856 10240
rect 16908 10231 16910 10240
rect 16856 10202 16908 10208
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 17052 9586 17080 9862
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 16764 7812 16816 7818
rect 16764 7754 16816 7760
rect 16776 7528 16804 7754
rect 16776 7500 16896 7528
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16776 7154 16804 7346
rect 16684 7126 16804 7154
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16684 6662 16712 7126
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16764 6656 16816 6662
rect 16764 6598 16816 6604
rect 16394 6488 16450 6497
rect 16394 6423 16396 6432
rect 16448 6423 16450 6432
rect 16396 6394 16448 6400
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 15384 5296 15436 5302
rect 15384 5238 15436 5244
rect 15396 5114 15424 5238
rect 15396 5086 15516 5114
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 14924 4752 14976 4758
rect 14924 4694 14976 4700
rect 15212 4690 15240 4966
rect 15016 4684 15068 4690
rect 15016 4626 15068 4632
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 15028 4010 15056 4626
rect 15200 4548 15252 4554
rect 15200 4490 15252 4496
rect 15016 4004 15068 4010
rect 15016 3946 15068 3952
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14844 3602 14872 3878
rect 15028 3602 15056 3946
rect 14832 3596 14884 3602
rect 14832 3538 14884 3544
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 15212 3058 15240 4490
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15396 2514 15424 4966
rect 15488 4554 15516 5086
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 15476 4548 15528 4554
rect 15476 4490 15528 4496
rect 16028 4548 16080 4554
rect 16028 4490 16080 4496
rect 16040 4282 16068 4490
rect 16028 4276 16080 4282
rect 16028 4218 16080 4224
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15580 3194 15608 3470
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 14280 2440 14332 2446
rect 14280 2382 14332 2388
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 14200 800 14228 2246
rect 14844 800 14872 2246
rect 15488 800 15516 2994
rect 15672 2922 15700 4014
rect 15752 3460 15804 3466
rect 15752 3402 15804 3408
rect 15764 3126 15792 3402
rect 15752 3120 15804 3126
rect 15752 3062 15804 3068
rect 16592 2922 16620 4626
rect 16684 4146 16712 6598
rect 16776 6254 16804 6598
rect 16868 6390 16896 7500
rect 17144 7002 17172 12406
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17328 11354 17356 12174
rect 17408 11824 17460 11830
rect 17408 11766 17460 11772
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17222 10160 17278 10169
rect 17222 10095 17278 10104
rect 17236 10062 17264 10095
rect 17224 10056 17276 10062
rect 17224 9998 17276 10004
rect 17328 9994 17356 11290
rect 17420 11014 17448 11766
rect 17604 11218 17632 12815
rect 17684 12786 17736 12792
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17696 11762 17724 12786
rect 17788 11830 17816 12786
rect 17776 11824 17828 11830
rect 17776 11766 17828 11772
rect 17684 11756 17736 11762
rect 17684 11698 17736 11704
rect 17776 11620 17828 11626
rect 17776 11562 17828 11568
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17788 11150 17816 11562
rect 17880 11354 17908 13262
rect 17972 12850 18000 13262
rect 18064 12850 18092 13484
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 17960 12708 18012 12714
rect 17960 12650 18012 12656
rect 17972 12442 18000 12650
rect 17960 12436 18012 12442
rect 18248 12434 18276 13670
rect 18340 12646 18368 19110
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18432 17338 18460 17478
rect 18524 17338 18552 19314
rect 18616 18086 18644 20810
rect 18708 20806 18736 22918
rect 18800 22681 18828 23054
rect 18786 22672 18842 22681
rect 18786 22607 18842 22616
rect 18788 22160 18840 22166
rect 18788 22102 18840 22108
rect 18800 21554 18828 22102
rect 18788 21548 18840 21554
rect 18788 21490 18840 21496
rect 18788 20868 18840 20874
rect 18788 20810 18840 20816
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18708 19446 18736 19790
rect 18696 19440 18748 19446
rect 18696 19382 18748 19388
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18512 17332 18564 17338
rect 18512 17274 18564 17280
rect 18616 17270 18644 17546
rect 18604 17264 18656 17270
rect 18604 17206 18656 17212
rect 18696 17264 18748 17270
rect 18696 17206 18748 17212
rect 18420 15904 18472 15910
rect 18420 15846 18472 15852
rect 18432 15502 18460 15846
rect 18512 15564 18564 15570
rect 18512 15506 18564 15512
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18524 13326 18552 15506
rect 18708 14890 18736 17206
rect 18696 14884 18748 14890
rect 18696 14826 18748 14832
rect 18708 14482 18736 14826
rect 18696 14476 18748 14482
rect 18696 14418 18748 14424
rect 18604 13796 18656 13802
rect 18604 13738 18656 13744
rect 18616 13326 18644 13738
rect 18512 13320 18564 13326
rect 18512 13262 18564 13268
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18524 12850 18552 13126
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 18248 12406 18368 12434
rect 17960 12378 18012 12384
rect 18236 12368 18288 12374
rect 18236 12310 18288 12316
rect 18248 11694 18276 12310
rect 18236 11688 18288 11694
rect 18236 11630 18288 11636
rect 18248 11354 18276 11630
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 18236 11348 18288 11354
rect 18236 11290 18288 11296
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17408 11008 17460 11014
rect 17408 10950 17460 10956
rect 17420 9994 17448 10950
rect 18340 10062 18368 12406
rect 18524 12238 18552 12786
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18616 12102 18644 12922
rect 18696 12776 18748 12782
rect 18694 12744 18696 12753
rect 18748 12744 18750 12753
rect 18694 12679 18750 12688
rect 18696 12368 18748 12374
rect 18696 12310 18748 12316
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18510 11248 18566 11257
rect 18510 11183 18566 11192
rect 18524 11150 18552 11183
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18708 10690 18736 12310
rect 18616 10662 18736 10690
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 17316 9988 17368 9994
rect 17316 9930 17368 9936
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17420 9042 17448 9930
rect 17500 9512 17552 9518
rect 17500 9454 17552 9460
rect 17408 9036 17460 9042
rect 17408 8978 17460 8984
rect 17316 8424 17368 8430
rect 17316 8366 17368 8372
rect 17328 8090 17356 8366
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17224 7404 17276 7410
rect 17328 7392 17356 8026
rect 17276 7364 17356 7392
rect 17224 7346 17276 7352
rect 17328 7206 17356 7364
rect 17316 7200 17368 7206
rect 17316 7142 17368 7148
rect 17132 6996 17184 7002
rect 17132 6938 17184 6944
rect 17132 6656 17184 6662
rect 17132 6598 17184 6604
rect 17144 6458 17172 6598
rect 17132 6452 17184 6458
rect 17132 6394 17184 6400
rect 16856 6384 16908 6390
rect 16856 6326 16908 6332
rect 16764 6248 16816 6254
rect 16764 6190 16816 6196
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 17052 5302 17080 5510
rect 17040 5296 17092 5302
rect 17040 5238 17092 5244
rect 17040 5160 17092 5166
rect 17236 5148 17264 6190
rect 17512 5166 17540 9454
rect 17604 9382 17632 9998
rect 17776 9920 17828 9926
rect 17776 9862 17828 9868
rect 17788 9586 17816 9862
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17788 8906 17816 9522
rect 18236 9036 18288 9042
rect 18236 8978 18288 8984
rect 17776 8900 17828 8906
rect 17776 8842 17828 8848
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17604 7546 17632 8434
rect 17684 8424 17736 8430
rect 17684 8366 17736 8372
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 17696 7274 17724 8366
rect 17776 7812 17828 7818
rect 17776 7754 17828 7760
rect 17788 7478 17816 7754
rect 17776 7472 17828 7478
rect 17776 7414 17828 7420
rect 17684 7268 17736 7274
rect 17684 7210 17736 7216
rect 17684 6384 17736 6390
rect 17684 6326 17736 6332
rect 17696 5302 17724 6326
rect 17684 5296 17736 5302
rect 17684 5238 17736 5244
rect 17092 5120 17264 5148
rect 17040 5102 17092 5108
rect 17236 4622 17264 5120
rect 17500 5160 17552 5166
rect 17500 5102 17552 5108
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16868 4078 16896 4422
rect 16948 4208 17000 4214
rect 16948 4150 17000 4156
rect 16856 4072 16908 4078
rect 16856 4014 16908 4020
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 16684 3058 16712 3130
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 15660 2916 15712 2922
rect 15660 2858 15712 2864
rect 16580 2916 16632 2922
rect 16580 2858 16632 2864
rect 15672 2774 15700 2858
rect 15580 2746 15700 2774
rect 15580 2446 15608 2746
rect 16684 2514 16712 2994
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 16868 2446 16896 4014
rect 16960 3534 16988 4150
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 16948 3528 17000 3534
rect 16948 3470 17000 3476
rect 17052 3194 17080 3878
rect 17144 3194 17172 3878
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 17236 3058 17264 4558
rect 17696 4554 17724 5238
rect 17684 4548 17736 4554
rect 17684 4490 17736 4496
rect 17696 4214 17724 4490
rect 17684 4208 17736 4214
rect 17684 4150 17736 4156
rect 17880 3670 17908 8570
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 17972 7546 18000 8366
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 18156 7206 18184 7822
rect 18248 7410 18276 8978
rect 18340 8974 18368 9998
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 18340 8362 18368 8910
rect 18328 8356 18380 8362
rect 18328 8298 18380 8304
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18432 7206 18460 8230
rect 18144 7200 18196 7206
rect 18144 7142 18196 7148
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18616 6730 18644 10662
rect 18696 10532 18748 10538
rect 18696 10474 18748 10480
rect 18708 10266 18736 10474
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18696 9512 18748 9518
rect 18696 9454 18748 9460
rect 18708 8498 18736 9454
rect 18800 8634 18828 20810
rect 18892 19718 18920 24686
rect 18972 24336 19024 24342
rect 18972 24278 19024 24284
rect 18984 23798 19012 24278
rect 18972 23792 19024 23798
rect 18972 23734 19024 23740
rect 18984 21010 19012 23734
rect 19076 23662 19104 24754
rect 19340 24744 19392 24750
rect 19260 24692 19340 24698
rect 19260 24686 19392 24692
rect 19260 24670 19380 24686
rect 19156 24200 19208 24206
rect 19156 24142 19208 24148
rect 19168 23866 19196 24142
rect 19156 23860 19208 23866
rect 19156 23802 19208 23808
rect 19064 23656 19116 23662
rect 19156 23656 19208 23662
rect 19064 23598 19116 23604
rect 19154 23624 19156 23633
rect 19208 23624 19210 23633
rect 19076 23254 19104 23598
rect 19154 23559 19210 23568
rect 19064 23248 19116 23254
rect 19064 23190 19116 23196
rect 19156 23248 19208 23254
rect 19156 23190 19208 23196
rect 18972 21004 19024 21010
rect 18972 20946 19024 20952
rect 18972 20800 19024 20806
rect 18972 20742 19024 20748
rect 18880 19712 18932 19718
rect 18880 19654 18932 19660
rect 18984 17814 19012 20742
rect 18972 17808 19024 17814
rect 18972 17750 19024 17756
rect 19168 17542 19196 23190
rect 19260 22982 19288 24670
rect 19338 23760 19394 23769
rect 19338 23695 19394 23704
rect 19352 23662 19380 23695
rect 19340 23656 19392 23662
rect 19340 23598 19392 23604
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 19352 23118 19380 23462
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 19340 22636 19392 22642
rect 19340 22578 19392 22584
rect 19352 22234 19380 22578
rect 19340 22228 19392 22234
rect 19340 22170 19392 22176
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 19352 19786 19380 21830
rect 19444 21486 19472 26823
rect 19524 24268 19576 24274
rect 19524 24210 19576 24216
rect 19536 23905 19564 24210
rect 19522 23896 19578 23905
rect 19522 23831 19578 23840
rect 19524 23724 19576 23730
rect 19524 23666 19576 23672
rect 19536 23322 19564 23666
rect 19524 23316 19576 23322
rect 19524 23258 19576 23264
rect 19536 23050 19564 23258
rect 19524 23044 19576 23050
rect 19524 22986 19576 22992
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19536 19854 19564 22986
rect 19720 22250 19748 26982
rect 19628 22222 19748 22250
rect 19628 22098 19656 22222
rect 19616 22092 19668 22098
rect 19812 22094 19840 27254
rect 19892 27124 19944 27130
rect 19892 27066 19944 27072
rect 19904 26994 19932 27066
rect 19892 26988 19944 26994
rect 19892 26930 19944 26936
rect 19892 24880 19944 24886
rect 19892 24822 19944 24828
rect 19904 24342 19932 24822
rect 19892 24336 19944 24342
rect 19892 24278 19944 24284
rect 19996 24154 20024 29650
rect 20352 27940 20404 27946
rect 20352 27882 20404 27888
rect 20364 27470 20392 27882
rect 20352 27464 20404 27470
rect 20352 27406 20404 27412
rect 20260 27328 20312 27334
rect 20260 27270 20312 27276
rect 20272 26994 20300 27270
rect 20076 26988 20128 26994
rect 20076 26930 20128 26936
rect 20260 26988 20312 26994
rect 20260 26930 20312 26936
rect 20088 26586 20116 26930
rect 20076 26580 20128 26586
rect 20456 26568 20484 30738
rect 20916 30682 20944 31078
rect 21008 30938 21036 31282
rect 20996 30932 21048 30938
rect 20996 30874 21048 30880
rect 21100 30802 21128 31962
rect 21364 31748 21416 31754
rect 21364 31690 21416 31696
rect 21180 31680 21232 31686
rect 21180 31622 21232 31628
rect 21192 31482 21220 31622
rect 21376 31482 21404 31690
rect 21180 31476 21232 31482
rect 21180 31418 21232 31424
rect 21364 31476 21416 31482
rect 21364 31418 21416 31424
rect 21088 30796 21140 30802
rect 21088 30738 21140 30744
rect 20824 30654 20944 30682
rect 21376 30666 21404 31418
rect 21364 30660 21416 30666
rect 20720 29504 20772 29510
rect 20720 29446 20772 29452
rect 20732 29170 20760 29446
rect 20720 29164 20772 29170
rect 20720 29106 20772 29112
rect 20824 29102 20852 30654
rect 21364 30602 21416 30608
rect 20996 30592 21048 30598
rect 20996 30534 21048 30540
rect 20904 29164 20956 29170
rect 20904 29106 20956 29112
rect 20812 29096 20864 29102
rect 20718 29064 20774 29073
rect 20812 29038 20864 29044
rect 20718 28999 20720 29008
rect 20772 28999 20774 29008
rect 20720 28970 20772 28976
rect 20824 28014 20852 29038
rect 20916 28762 20944 29106
rect 20904 28756 20956 28762
rect 20904 28698 20956 28704
rect 20904 28416 20956 28422
rect 20904 28358 20956 28364
rect 20812 28008 20864 28014
rect 20812 27950 20864 27956
rect 20536 27872 20588 27878
rect 20536 27814 20588 27820
rect 20076 26522 20128 26528
rect 20364 26540 20484 26568
rect 20364 26382 20392 26540
rect 20444 26444 20496 26450
rect 20444 26386 20496 26392
rect 20352 26376 20404 26382
rect 20352 26318 20404 26324
rect 20260 25288 20312 25294
rect 20260 25230 20312 25236
rect 20166 24984 20222 24993
rect 20272 24954 20300 25230
rect 20166 24919 20222 24928
rect 20260 24948 20312 24954
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 20088 24274 20116 24754
rect 20076 24268 20128 24274
rect 20076 24210 20128 24216
rect 19996 24126 20116 24154
rect 20088 24070 20116 24126
rect 19984 24064 20036 24070
rect 19890 24032 19946 24041
rect 19984 24006 20036 24012
rect 20076 24064 20128 24070
rect 20076 24006 20128 24012
rect 19890 23967 19946 23976
rect 19904 23866 19932 23967
rect 19892 23860 19944 23866
rect 19892 23802 19944 23808
rect 19892 23724 19944 23730
rect 19892 23666 19944 23672
rect 19904 22642 19932 23666
rect 19996 22982 20024 24006
rect 20076 23520 20128 23526
rect 20180 23508 20208 24919
rect 20260 24890 20312 24896
rect 20364 23798 20392 26318
rect 20456 24041 20484 26386
rect 20442 24032 20498 24041
rect 20442 23967 20498 23976
rect 20456 23866 20484 23967
rect 20444 23860 20496 23866
rect 20444 23802 20496 23808
rect 20352 23792 20404 23798
rect 20352 23734 20404 23740
rect 20128 23480 20208 23508
rect 20076 23462 20128 23468
rect 20076 23112 20128 23118
rect 20076 23054 20128 23060
rect 19984 22976 20036 22982
rect 19984 22918 20036 22924
rect 19892 22636 19944 22642
rect 19892 22578 19944 22584
rect 19984 22500 20036 22506
rect 19984 22442 20036 22448
rect 19890 22264 19946 22273
rect 19890 22199 19946 22208
rect 19616 22034 19668 22040
rect 19720 22066 19840 22094
rect 19628 20942 19656 22034
rect 19616 20936 19668 20942
rect 19616 20878 19668 20884
rect 19720 19922 19748 22066
rect 19904 22030 19932 22199
rect 19996 22166 20024 22442
rect 19984 22160 20036 22166
rect 19984 22102 20036 22108
rect 19892 22024 19944 22030
rect 19892 21966 19944 21972
rect 19800 21888 19852 21894
rect 19800 21830 19852 21836
rect 19892 21888 19944 21894
rect 19892 21830 19944 21836
rect 19812 21729 19840 21830
rect 19798 21720 19854 21729
rect 19798 21655 19854 21664
rect 19800 21004 19852 21010
rect 19800 20946 19852 20952
rect 19812 20602 19840 20946
rect 19800 20596 19852 20602
rect 19800 20538 19852 20544
rect 19708 19916 19760 19922
rect 19708 19858 19760 19864
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19340 19780 19392 19786
rect 19340 19722 19392 19728
rect 19616 19780 19668 19786
rect 19616 19722 19668 19728
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 19260 17610 19288 19314
rect 19340 17740 19392 17746
rect 19340 17682 19392 17688
rect 19248 17604 19300 17610
rect 19248 17546 19300 17552
rect 19156 17536 19208 17542
rect 19156 17478 19208 17484
rect 19260 17270 19288 17546
rect 19248 17264 19300 17270
rect 19248 17206 19300 17212
rect 19156 16992 19208 16998
rect 19156 16934 19208 16940
rect 19064 16788 19116 16794
rect 19064 16730 19116 16736
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 18892 14482 18920 14554
rect 18880 14476 18932 14482
rect 18880 14418 18932 14424
rect 18892 13190 18920 14418
rect 18972 14340 19024 14346
rect 18972 14282 19024 14288
rect 18984 14006 19012 14282
rect 18972 14000 19024 14006
rect 18972 13942 19024 13948
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18984 12986 19012 13194
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 18880 12912 18932 12918
rect 18880 12854 18932 12860
rect 18892 12238 18920 12854
rect 18972 12844 19024 12850
rect 18972 12786 19024 12792
rect 18984 12442 19012 12786
rect 18972 12436 19024 12442
rect 18972 12378 19024 12384
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18972 12232 19024 12238
rect 18972 12174 19024 12180
rect 18984 11898 19012 12174
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 19076 10146 19104 16730
rect 19168 12186 19196 16934
rect 19352 15638 19380 17682
rect 19628 17270 19656 19722
rect 19708 18692 19760 18698
rect 19708 18634 19760 18640
rect 19616 17264 19668 17270
rect 19616 17206 19668 17212
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19444 16658 19472 17138
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 19628 16454 19656 17206
rect 19616 16448 19668 16454
rect 19616 16390 19668 16396
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 19340 15632 19392 15638
rect 19340 15574 19392 15580
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19248 13932 19300 13938
rect 19248 13874 19300 13880
rect 19260 12442 19288 13874
rect 19352 13326 19380 14962
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19352 12442 19380 13262
rect 19248 12436 19300 12442
rect 19248 12378 19300 12384
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19168 12158 19288 12186
rect 19352 12170 19380 12378
rect 19444 12306 19472 15642
rect 19628 15026 19656 16390
rect 19616 15020 19668 15026
rect 19616 14962 19668 14968
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19536 14618 19564 14758
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 19536 12442 19564 13670
rect 19524 12436 19576 12442
rect 19524 12378 19576 12384
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19156 12096 19208 12102
rect 19156 12038 19208 12044
rect 19168 11898 19196 12038
rect 19156 11892 19208 11898
rect 19156 11834 19208 11840
rect 19260 11354 19288 12158
rect 19340 12164 19392 12170
rect 19340 12106 19392 12112
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19340 11076 19392 11082
rect 19340 11018 19392 11024
rect 19076 10118 19196 10146
rect 19352 10130 19380 11018
rect 19444 10146 19472 12242
rect 19524 11756 19576 11762
rect 19524 11698 19576 11704
rect 19536 11665 19564 11698
rect 19522 11656 19578 11665
rect 19522 11591 19578 11600
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19536 10266 19564 10406
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 19064 10056 19116 10062
rect 19064 9998 19116 10004
rect 19076 9654 19104 9998
rect 19064 9648 19116 9654
rect 19064 9590 19116 9596
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 19168 8498 19196 10118
rect 19340 10124 19392 10130
rect 19444 10118 19564 10146
rect 19628 10130 19656 14350
rect 19720 13161 19748 18634
rect 19800 17808 19852 17814
rect 19800 17750 19852 17756
rect 19812 17202 19840 17750
rect 19800 17196 19852 17202
rect 19800 17138 19852 17144
rect 19800 16652 19852 16658
rect 19800 16594 19852 16600
rect 19812 15026 19840 16594
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19798 14648 19854 14657
rect 19798 14583 19800 14592
rect 19852 14583 19854 14592
rect 19800 14554 19852 14560
rect 19800 14476 19852 14482
rect 19800 14418 19852 14424
rect 19812 13258 19840 14418
rect 19904 13938 19932 21830
rect 20088 19854 20116 23054
rect 20364 22778 20392 23734
rect 20352 22772 20404 22778
rect 20352 22714 20404 22720
rect 20352 22636 20404 22642
rect 20352 22578 20404 22584
rect 20168 22568 20220 22574
rect 20168 22510 20220 22516
rect 20180 22234 20208 22510
rect 20168 22228 20220 22234
rect 20168 22170 20220 22176
rect 20180 20058 20208 22170
rect 20260 22024 20312 22030
rect 20260 21966 20312 21972
rect 20272 21690 20300 21966
rect 20364 21690 20392 22578
rect 20444 22500 20496 22506
rect 20444 22442 20496 22448
rect 20456 22409 20484 22442
rect 20442 22400 20498 22409
rect 20442 22335 20498 22344
rect 20548 22216 20576 27814
rect 20916 27606 20944 28358
rect 20904 27600 20956 27606
rect 20904 27542 20956 27548
rect 20812 27532 20864 27538
rect 20812 27474 20864 27480
rect 20628 27464 20680 27470
rect 20628 27406 20680 27412
rect 20640 26994 20668 27406
rect 20824 27130 20852 27474
rect 20812 27124 20864 27130
rect 20812 27066 20864 27072
rect 20628 26988 20680 26994
rect 20628 26930 20680 26936
rect 20640 25498 20668 26930
rect 20720 26784 20772 26790
rect 20718 26752 20720 26761
rect 20772 26752 20774 26761
rect 20718 26687 20774 26696
rect 20812 26240 20864 26246
rect 20812 26182 20864 26188
rect 20628 25492 20680 25498
rect 20628 25434 20680 25440
rect 20824 25362 20852 26182
rect 20812 25356 20864 25362
rect 20812 25298 20864 25304
rect 20628 24880 20680 24886
rect 20628 24822 20680 24828
rect 20640 24206 20668 24822
rect 20720 24812 20772 24818
rect 20720 24754 20772 24760
rect 20628 24200 20680 24206
rect 20628 24142 20680 24148
rect 20628 23792 20680 23798
rect 20628 23734 20680 23740
rect 20640 22778 20668 23734
rect 20628 22772 20680 22778
rect 20628 22714 20680 22720
rect 20732 22216 20760 24754
rect 20824 23662 20852 25298
rect 20904 24336 20956 24342
rect 20904 24278 20956 24284
rect 20916 24138 20944 24278
rect 20904 24132 20956 24138
rect 20904 24074 20956 24080
rect 20812 23656 20864 23662
rect 20812 23598 20864 23604
rect 20824 22642 20852 23598
rect 20916 23118 20944 24074
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 21008 22522 21036 30534
rect 21180 30320 21232 30326
rect 21180 30262 21232 30268
rect 21192 29238 21220 30262
rect 21468 29850 21496 32438
rect 21824 32224 21876 32230
rect 21824 32166 21876 32172
rect 21836 32065 21864 32166
rect 21822 32056 21878 32065
rect 21822 31991 21878 32000
rect 21824 31476 21876 31482
rect 21824 31418 21876 31424
rect 21640 31136 21692 31142
rect 21640 31078 21692 31084
rect 21456 29844 21508 29850
rect 21456 29786 21508 29792
rect 21180 29232 21232 29238
rect 21180 29174 21232 29180
rect 21468 29170 21496 29786
rect 21088 29164 21140 29170
rect 21088 29106 21140 29112
rect 21456 29164 21508 29170
rect 21456 29106 21508 29112
rect 21548 29164 21600 29170
rect 21548 29106 21600 29112
rect 21100 28422 21128 29106
rect 21272 29096 21324 29102
rect 21560 29073 21588 29106
rect 21272 29038 21324 29044
rect 21546 29064 21602 29073
rect 21180 28552 21232 28558
rect 21178 28520 21180 28529
rect 21232 28520 21234 28529
rect 21178 28455 21234 28464
rect 21088 28416 21140 28422
rect 21088 28358 21140 28364
rect 21178 28248 21234 28257
rect 21178 28183 21234 28192
rect 21088 27940 21140 27946
rect 21088 27882 21140 27888
rect 21100 25294 21128 27882
rect 21088 25288 21140 25294
rect 21088 25230 21140 25236
rect 21086 24848 21142 24857
rect 21086 24783 21142 24792
rect 21100 24682 21128 24783
rect 21088 24676 21140 24682
rect 21088 24618 21140 24624
rect 20456 22188 20576 22216
rect 20640 22188 20760 22216
rect 20824 22494 21036 22522
rect 20260 21684 20312 21690
rect 20260 21626 20312 21632
rect 20352 21684 20404 21690
rect 20352 21626 20404 21632
rect 20272 21418 20300 21626
rect 20260 21412 20312 21418
rect 20260 21354 20312 21360
rect 20456 20942 20484 22188
rect 20534 22128 20590 22137
rect 20534 22063 20590 22072
rect 20444 20936 20496 20942
rect 20444 20878 20496 20884
rect 20444 20256 20496 20262
rect 20442 20224 20444 20233
rect 20496 20224 20498 20233
rect 20442 20159 20498 20168
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 20548 19938 20576 22063
rect 20640 22012 20668 22188
rect 20640 21984 20760 22012
rect 20628 21616 20680 21622
rect 20628 21558 20680 21564
rect 20640 21350 20668 21558
rect 20628 21344 20680 21350
rect 20628 21286 20680 21292
rect 20628 20936 20680 20942
rect 20628 20878 20680 20884
rect 20640 20398 20668 20878
rect 20628 20392 20680 20398
rect 20626 20360 20628 20369
rect 20680 20360 20682 20369
rect 20626 20295 20682 20304
rect 20456 19910 20576 19938
rect 20076 19848 20128 19854
rect 20074 19816 20076 19825
rect 20128 19816 20130 19825
rect 20074 19751 20130 19760
rect 20456 19334 20484 19910
rect 20536 19848 20588 19854
rect 20536 19790 20588 19796
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20548 19689 20576 19790
rect 20534 19680 20590 19689
rect 20534 19615 20590 19624
rect 20364 19306 20484 19334
rect 20260 18896 20312 18902
rect 20260 18838 20312 18844
rect 20272 18426 20300 18838
rect 20364 18766 20392 19306
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 20260 18420 20312 18426
rect 20260 18362 20312 18368
rect 20168 17128 20220 17134
rect 20168 17070 20220 17076
rect 19984 16992 20036 16998
rect 19984 16934 20036 16940
rect 19996 16454 20024 16934
rect 19984 16448 20036 16454
rect 19984 16390 20036 16396
rect 20180 15094 20208 17070
rect 20168 15088 20220 15094
rect 20168 15030 20220 15036
rect 19984 15020 20036 15026
rect 20036 14980 20116 15008
rect 19984 14962 20036 14968
rect 20088 14074 20116 14980
rect 20168 14544 20220 14550
rect 20166 14512 20168 14521
rect 20220 14512 20222 14521
rect 20166 14447 20222 14456
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 19892 13932 19944 13938
rect 19892 13874 19944 13880
rect 19892 13796 19944 13802
rect 19892 13738 19944 13744
rect 19800 13252 19852 13258
rect 19800 13194 19852 13200
rect 19706 13152 19762 13161
rect 19706 13087 19762 13096
rect 19708 12980 19760 12986
rect 19708 12922 19760 12928
rect 19720 12442 19748 12922
rect 19812 12646 19840 13194
rect 19800 12640 19852 12646
rect 19800 12582 19852 12588
rect 19904 12442 19932 13738
rect 20088 13326 20116 14010
rect 20180 13870 20208 14350
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 19708 12436 19760 12442
rect 19708 12378 19760 12384
rect 19892 12436 19944 12442
rect 19892 12378 19944 12384
rect 19800 12232 19852 12238
rect 19720 12180 19800 12186
rect 19720 12174 19852 12180
rect 19720 12158 19840 12174
rect 19720 11082 19748 12158
rect 19800 11620 19852 11626
rect 19996 11608 20024 13262
rect 20088 12850 20116 13262
rect 20180 12986 20208 13806
rect 20272 13802 20300 18362
rect 20364 14346 20392 18702
rect 20442 16688 20498 16697
rect 20442 16623 20444 16632
rect 20496 16623 20498 16632
rect 20444 16594 20496 16600
rect 20548 15502 20576 19615
rect 20640 18970 20668 19790
rect 20732 19334 20760 21984
rect 20824 21554 20852 22494
rect 20904 22432 20956 22438
rect 20904 22374 20956 22380
rect 21088 22432 21140 22438
rect 21088 22374 21140 22380
rect 20916 22030 20944 22374
rect 21100 22234 21128 22374
rect 21088 22228 21140 22234
rect 21088 22170 21140 22176
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 20996 21956 21048 21962
rect 20996 21898 21048 21904
rect 20812 21548 20864 21554
rect 20812 21490 20864 21496
rect 20824 21078 20852 21490
rect 20812 21072 20864 21078
rect 20812 21014 20864 21020
rect 20810 20904 20866 20913
rect 20810 20839 20812 20848
rect 20864 20839 20866 20848
rect 20812 20810 20864 20816
rect 20904 20800 20956 20806
rect 20810 20768 20866 20777
rect 20866 20748 20904 20754
rect 20866 20742 20956 20748
rect 20866 20726 20944 20742
rect 20810 20703 20866 20712
rect 20824 19854 20852 20703
rect 20812 19848 20864 19854
rect 20812 19790 20864 19796
rect 20824 19514 20852 19790
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20732 19306 20852 19334
rect 20628 18964 20680 18970
rect 20628 18906 20680 18912
rect 20640 18748 20668 18906
rect 20720 18760 20772 18766
rect 20640 18720 20720 18748
rect 20720 18702 20772 18708
rect 20824 17762 20852 19306
rect 20732 17734 20852 17762
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 20640 17066 20668 17274
rect 20628 17060 20680 17066
rect 20628 17002 20680 17008
rect 20628 16652 20680 16658
rect 20628 16594 20680 16600
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20444 14952 20496 14958
rect 20444 14894 20496 14900
rect 20352 14340 20404 14346
rect 20352 14282 20404 14288
rect 20352 14000 20404 14006
rect 20352 13942 20404 13948
rect 20260 13796 20312 13802
rect 20260 13738 20312 13744
rect 20364 13326 20392 13942
rect 20352 13320 20404 13326
rect 20352 13262 20404 13268
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20076 12844 20128 12850
rect 20076 12786 20128 12792
rect 20364 12442 20392 13262
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 20168 12300 20220 12306
rect 20088 12260 20168 12288
rect 20088 11762 20116 12260
rect 20168 12242 20220 12248
rect 20076 11756 20128 11762
rect 20076 11698 20128 11704
rect 20260 11756 20312 11762
rect 20364 11744 20392 12378
rect 20312 11716 20392 11744
rect 20260 11698 20312 11704
rect 19852 11580 20024 11608
rect 20168 11620 20220 11626
rect 19800 11562 19852 11568
rect 20168 11562 20220 11568
rect 19708 11076 19760 11082
rect 19708 11018 19760 11024
rect 19340 10066 19392 10072
rect 19248 9988 19300 9994
rect 19248 9930 19300 9936
rect 19260 9586 19288 9930
rect 19352 9586 19380 10066
rect 19536 10062 19564 10118
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19524 10056 19576 10062
rect 19812 10033 19840 11562
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 19984 10192 20036 10198
rect 19984 10134 20036 10140
rect 19996 10062 20024 10134
rect 19984 10056 20036 10062
rect 19524 9998 19576 10004
rect 19798 10024 19854 10033
rect 19432 9988 19484 9994
rect 19432 9930 19484 9936
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 18800 8090 18828 8434
rect 18880 8356 18932 8362
rect 18880 8298 18932 8304
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 18604 6724 18656 6730
rect 18604 6666 18656 6672
rect 17960 6112 18012 6118
rect 17960 6054 18012 6060
rect 17972 4282 18000 6054
rect 18616 5778 18644 6666
rect 18800 5914 18828 7346
rect 18892 6866 18920 8298
rect 19168 7970 19196 8434
rect 19260 8430 19288 9522
rect 19352 9450 19380 9522
rect 19340 9444 19392 9450
rect 19340 9386 19392 9392
rect 19444 8566 19472 9930
rect 19536 9674 19564 9998
rect 19984 9998 20036 10004
rect 19798 9959 19800 9968
rect 19852 9959 19854 9968
rect 19800 9930 19852 9936
rect 19536 9646 19932 9674
rect 19616 8900 19668 8906
rect 19616 8842 19668 8848
rect 19432 8560 19484 8566
rect 19432 8502 19484 8508
rect 19628 8498 19656 8842
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 19430 8392 19486 8401
rect 19076 7942 19196 7970
rect 18972 7812 19024 7818
rect 18972 7754 19024 7760
rect 18984 7478 19012 7754
rect 18972 7472 19024 7478
rect 18972 7414 19024 7420
rect 18880 6860 18932 6866
rect 18880 6802 18932 6808
rect 19076 6458 19104 7942
rect 19156 7880 19208 7886
rect 19260 7868 19288 8366
rect 19430 8327 19486 8336
rect 19444 8090 19472 8327
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19340 7948 19392 7954
rect 19628 7936 19656 8434
rect 19392 7908 19656 7936
rect 19340 7890 19392 7896
rect 19208 7840 19288 7868
rect 19156 7822 19208 7828
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 18788 5908 18840 5914
rect 18788 5850 18840 5856
rect 18604 5772 18656 5778
rect 18604 5714 18656 5720
rect 18696 5772 18748 5778
rect 18696 5714 18748 5720
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 18144 5636 18196 5642
rect 18144 5578 18196 5584
rect 18156 5030 18184 5578
rect 18524 5370 18552 5646
rect 18512 5364 18564 5370
rect 18512 5306 18564 5312
rect 18616 5234 18644 5714
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 17960 4276 18012 4282
rect 17960 4218 18012 4224
rect 17868 3664 17920 3670
rect 17868 3606 17920 3612
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 17420 2514 17448 3334
rect 17880 2990 17908 3606
rect 17868 2984 17920 2990
rect 17868 2926 17920 2932
rect 17408 2508 17460 2514
rect 17408 2450 17460 2456
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 17972 2378 18000 4218
rect 18156 2774 18184 4966
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18340 4078 18368 4422
rect 18616 4078 18644 5170
rect 18708 4146 18736 5714
rect 18800 5710 18828 5850
rect 18788 5704 18840 5710
rect 19076 5692 19104 6394
rect 19352 6390 19380 7142
rect 19628 6934 19656 7908
rect 19904 7732 19932 9646
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19996 8498 20024 8774
rect 20088 8634 20116 11494
rect 20180 8906 20208 11562
rect 20364 11218 20392 11716
rect 20456 11558 20484 14894
rect 20548 14414 20576 15302
rect 20640 15162 20668 16594
rect 20732 16522 20760 17734
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20824 16561 20852 17614
rect 20810 16552 20866 16561
rect 20720 16516 20772 16522
rect 20810 16487 20812 16496
rect 20720 16458 20772 16464
rect 20864 16487 20866 16496
rect 20904 16516 20956 16522
rect 20812 16458 20864 16464
rect 20904 16458 20956 16464
rect 20732 15978 20760 16458
rect 20720 15972 20772 15978
rect 20720 15914 20772 15920
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20640 14618 20668 15098
rect 20916 14906 20944 16458
rect 20732 14878 20944 14906
rect 20732 14822 20760 14878
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 20536 14408 20588 14414
rect 20588 14368 20668 14396
rect 20536 14350 20588 14356
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20548 12238 20576 14214
rect 20640 13258 20668 14368
rect 20732 13938 20760 14758
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20718 13424 20774 13433
rect 20718 13359 20720 13368
rect 20772 13359 20774 13368
rect 20720 13330 20772 13336
rect 20628 13252 20680 13258
rect 20628 13194 20680 13200
rect 20824 13138 20852 14758
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 20640 13110 20852 13138
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 20548 11286 20576 12174
rect 20536 11280 20588 11286
rect 20536 11222 20588 11228
rect 20352 11212 20404 11218
rect 20352 11154 20404 11160
rect 20260 11076 20312 11082
rect 20260 11018 20312 11024
rect 20272 8906 20300 11018
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20364 10266 20392 10406
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20640 9704 20668 13110
rect 20812 12980 20864 12986
rect 20812 12922 20864 12928
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 20732 11694 20760 12038
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20824 11218 20852 12922
rect 20916 11762 20944 13262
rect 21008 12986 21036 21898
rect 21192 20754 21220 28183
rect 21284 24954 21312 29038
rect 21546 28999 21602 29008
rect 21364 28552 21416 28558
rect 21364 28494 21416 28500
rect 21376 26897 21404 28494
rect 21454 28384 21510 28393
rect 21454 28319 21510 28328
rect 21468 28150 21496 28319
rect 21652 28200 21680 31078
rect 21732 30728 21784 30734
rect 21732 30670 21784 30676
rect 21744 30190 21772 30670
rect 21836 30666 21864 31418
rect 21824 30660 21876 30666
rect 21824 30602 21876 30608
rect 21732 30184 21784 30190
rect 21732 30126 21784 30132
rect 21916 29844 21968 29850
rect 21916 29786 21968 29792
rect 21928 29510 21956 29786
rect 21916 29504 21968 29510
rect 21916 29446 21968 29452
rect 21732 29028 21784 29034
rect 21732 28970 21784 28976
rect 21560 28172 21680 28200
rect 21456 28144 21508 28150
rect 21456 28086 21508 28092
rect 21456 28008 21508 28014
rect 21456 27950 21508 27956
rect 21468 26926 21496 27950
rect 21456 26920 21508 26926
rect 21362 26888 21418 26897
rect 21456 26862 21508 26868
rect 21362 26823 21418 26832
rect 21364 26784 21416 26790
rect 21364 26726 21416 26732
rect 21376 26382 21404 26726
rect 21364 26376 21416 26382
rect 21364 26318 21416 26324
rect 21272 24948 21324 24954
rect 21272 24890 21324 24896
rect 21284 23798 21312 24890
rect 21376 24750 21404 26318
rect 21468 25362 21496 26862
rect 21456 25356 21508 25362
rect 21456 25298 21508 25304
rect 21364 24744 21416 24750
rect 21364 24686 21416 24692
rect 21456 24744 21508 24750
rect 21456 24686 21508 24692
rect 21468 24614 21496 24686
rect 21456 24608 21508 24614
rect 21456 24550 21508 24556
rect 21272 23792 21324 23798
rect 21324 23752 21404 23780
rect 21272 23734 21324 23740
rect 21272 23520 21324 23526
rect 21272 23462 21324 23468
rect 21284 22438 21312 23462
rect 21376 23118 21404 23752
rect 21364 23112 21416 23118
rect 21364 23054 21416 23060
rect 21456 23044 21508 23050
rect 21456 22986 21508 22992
rect 21364 22976 21416 22982
rect 21364 22918 21416 22924
rect 21272 22432 21324 22438
rect 21272 22374 21324 22380
rect 21100 20726 21220 20754
rect 21100 13138 21128 20726
rect 21284 20074 21312 22374
rect 21376 22094 21404 22918
rect 21468 22710 21496 22986
rect 21456 22704 21508 22710
rect 21456 22646 21508 22652
rect 21560 22098 21588 28172
rect 21640 28076 21692 28082
rect 21640 28018 21692 28024
rect 21376 22066 21496 22094
rect 21364 22024 21416 22030
rect 21364 21966 21416 21972
rect 21376 21865 21404 21966
rect 21362 21856 21418 21865
rect 21362 21791 21418 21800
rect 21362 21720 21418 21729
rect 21362 21655 21364 21664
rect 21416 21655 21418 21664
rect 21364 21626 21416 21632
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 21192 20046 21312 20074
rect 21192 19990 21220 20046
rect 21376 19990 21404 20402
rect 21180 19984 21232 19990
rect 21180 19926 21232 19932
rect 21272 19984 21324 19990
rect 21272 19926 21324 19932
rect 21364 19984 21416 19990
rect 21364 19926 21416 19932
rect 21284 19854 21312 19926
rect 21272 19848 21324 19854
rect 21272 19790 21324 19796
rect 21284 19689 21312 19790
rect 21270 19680 21326 19689
rect 21270 19615 21326 19624
rect 21364 19508 21416 19514
rect 21364 19450 21416 19456
rect 21270 19408 21326 19417
rect 21270 19343 21272 19352
rect 21324 19343 21326 19352
rect 21272 19314 21324 19320
rect 21272 18828 21324 18834
rect 21272 18770 21324 18776
rect 21178 18728 21234 18737
rect 21178 18663 21234 18672
rect 21192 16590 21220 18663
rect 21180 16584 21232 16590
rect 21180 16526 21232 16532
rect 21192 14890 21220 16526
rect 21284 15094 21312 18770
rect 21272 15088 21324 15094
rect 21272 15030 21324 15036
rect 21272 14952 21324 14958
rect 21272 14894 21324 14900
rect 21180 14884 21232 14890
rect 21180 14826 21232 14832
rect 21192 14482 21220 14826
rect 21180 14476 21232 14482
rect 21180 14418 21232 14424
rect 21284 14346 21312 14894
rect 21272 14340 21324 14346
rect 21272 14282 21324 14288
rect 21376 14226 21404 19450
rect 21284 14198 21404 14226
rect 21284 13802 21312 14198
rect 21272 13796 21324 13802
rect 21272 13738 21324 13744
rect 21180 13320 21232 13326
rect 21232 13280 21312 13308
rect 21180 13262 21232 13268
rect 21100 13110 21220 13138
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 20996 12164 21048 12170
rect 20996 12106 21048 12112
rect 21008 11830 21036 12106
rect 20996 11824 21048 11830
rect 20996 11766 21048 11772
rect 20904 11756 20956 11762
rect 20904 11698 20956 11704
rect 21100 11354 21128 12922
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 20812 11212 20864 11218
rect 20812 11154 20864 11160
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20456 9676 20668 9704
rect 20352 9376 20404 9382
rect 20352 9318 20404 9324
rect 20364 9178 20392 9318
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 20168 8900 20220 8906
rect 20168 8842 20220 8848
rect 20260 8900 20312 8906
rect 20260 8842 20312 8848
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 20272 8566 20300 8842
rect 20260 8560 20312 8566
rect 20260 8502 20312 8508
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 20088 8401 20116 8434
rect 20074 8392 20130 8401
rect 20074 8327 20130 8336
rect 20088 7886 20116 8327
rect 20364 8022 20392 9114
rect 20456 8294 20484 9676
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20548 8820 20576 9522
rect 20732 8906 20760 10950
rect 20810 10704 20866 10713
rect 21008 10674 21036 11290
rect 21088 10736 21140 10742
rect 21192 10724 21220 13110
rect 21284 12442 21312 13280
rect 21364 12844 21416 12850
rect 21364 12786 21416 12792
rect 21272 12436 21324 12442
rect 21272 12378 21324 12384
rect 21284 11694 21312 12378
rect 21272 11688 21324 11694
rect 21272 11630 21324 11636
rect 21376 11558 21404 12786
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21140 10696 21220 10724
rect 21088 10678 21140 10684
rect 20810 10639 20812 10648
rect 20864 10639 20866 10648
rect 20996 10668 21048 10674
rect 20812 10610 20864 10616
rect 20996 10610 21048 10616
rect 21008 10470 21036 10610
rect 20996 10464 21048 10470
rect 20996 10406 21048 10412
rect 20810 9616 20866 9625
rect 20810 9551 20812 9560
rect 20864 9551 20866 9560
rect 20812 9522 20864 9528
rect 20902 9480 20958 9489
rect 20902 9415 20958 9424
rect 20916 9382 20944 9415
rect 20904 9376 20956 9382
rect 20904 9318 20956 9324
rect 20996 9172 21048 9178
rect 20996 9114 21048 9120
rect 20812 9104 20864 9110
rect 20812 9046 20864 9052
rect 20902 9072 20958 9081
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 20628 8832 20680 8838
rect 20548 8792 20628 8820
rect 20628 8774 20680 8780
rect 20732 8566 20760 8842
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 20824 8498 20852 9046
rect 20902 9007 20958 9016
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20812 8492 20864 8498
rect 20812 8434 20864 8440
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 20352 8016 20404 8022
rect 20352 7958 20404 7964
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 20352 7880 20404 7886
rect 20456 7868 20484 8230
rect 20640 8022 20668 8434
rect 20916 8378 20944 9007
rect 21008 8634 21036 9114
rect 20996 8628 21048 8634
rect 20996 8570 21048 8576
rect 20824 8350 20944 8378
rect 20628 8016 20680 8022
rect 20628 7958 20680 7964
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 20404 7840 20484 7868
rect 20536 7880 20588 7886
rect 20352 7822 20404 7828
rect 20536 7822 20588 7828
rect 20076 7744 20128 7750
rect 19904 7704 20076 7732
rect 20076 7686 20128 7692
rect 20442 7712 20498 7721
rect 20442 7647 20498 7656
rect 20456 7546 20484 7647
rect 20444 7540 20496 7546
rect 20444 7482 20496 7488
rect 20548 7002 20576 7822
rect 20628 7812 20680 7818
rect 20628 7754 20680 7760
rect 20640 7002 20668 7754
rect 20732 7410 20760 7890
rect 20824 7478 20852 8350
rect 20904 8288 20956 8294
rect 20904 8230 20956 8236
rect 20916 7954 20944 8230
rect 20904 7948 20956 7954
rect 20904 7890 20956 7896
rect 21100 7528 21128 10678
rect 21284 10674 21312 11290
rect 21468 11082 21496 22066
rect 21548 22092 21600 22098
rect 21548 22034 21600 22040
rect 21548 21956 21600 21962
rect 21548 21898 21600 21904
rect 21560 21350 21588 21898
rect 21548 21344 21600 21350
rect 21548 21286 21600 21292
rect 21548 20800 21600 20806
rect 21548 20742 21600 20748
rect 21560 15706 21588 20742
rect 21652 19514 21680 28018
rect 21744 21894 21772 28970
rect 21824 28076 21876 28082
rect 21824 28018 21876 28024
rect 21836 27713 21864 28018
rect 21822 27704 21878 27713
rect 21822 27639 21878 27648
rect 21824 26988 21876 26994
rect 21824 26930 21876 26936
rect 21836 26353 21864 26930
rect 21822 26344 21878 26353
rect 21822 26279 21878 26288
rect 21824 24880 21876 24886
rect 21824 24822 21876 24828
rect 21836 24698 21864 24822
rect 21928 24818 21956 29446
rect 21916 24812 21968 24818
rect 21916 24754 21968 24760
rect 21836 24670 21956 24698
rect 21824 24608 21876 24614
rect 21824 24550 21876 24556
rect 21836 23361 21864 24550
rect 21822 23352 21878 23361
rect 21822 23287 21878 23296
rect 21822 22400 21878 22409
rect 21822 22335 21878 22344
rect 21836 22166 21864 22335
rect 21928 22273 21956 24670
rect 21914 22264 21970 22273
rect 21914 22199 21970 22208
rect 21824 22160 21876 22166
rect 21824 22102 21876 22108
rect 22020 22001 22048 35634
rect 22296 35290 22324 36110
rect 22480 35834 22508 36110
rect 22572 36038 22600 37130
rect 23032 36718 23060 37606
rect 23860 37398 23888 37742
rect 23848 37392 23900 37398
rect 23848 37334 23900 37340
rect 25044 37120 25096 37126
rect 25044 37062 25096 37068
rect 24952 36916 25004 36922
rect 24952 36858 25004 36864
rect 23756 36780 23808 36786
rect 23756 36722 23808 36728
rect 23020 36712 23072 36718
rect 23020 36654 23072 36660
rect 23032 36174 23060 36654
rect 23020 36168 23072 36174
rect 23020 36110 23072 36116
rect 22560 36032 22612 36038
rect 22560 35974 22612 35980
rect 22468 35828 22520 35834
rect 22468 35770 22520 35776
rect 23032 35698 23060 36110
rect 23480 36032 23532 36038
rect 23480 35974 23532 35980
rect 23492 35834 23520 35974
rect 23480 35828 23532 35834
rect 23480 35770 23532 35776
rect 23768 35737 23796 36722
rect 24768 36712 24820 36718
rect 24768 36654 24820 36660
rect 24780 36242 24808 36654
rect 24768 36236 24820 36242
rect 24768 36178 24820 36184
rect 24964 35766 24992 36858
rect 25056 36854 25084 37062
rect 25044 36848 25096 36854
rect 25044 36790 25096 36796
rect 25148 36106 25176 43101
rect 25792 41414 25820 43101
rect 25700 41386 25820 41414
rect 25228 38956 25280 38962
rect 25228 38898 25280 38904
rect 25240 38654 25268 38898
rect 25504 38888 25556 38894
rect 25504 38830 25556 38836
rect 25240 38626 25360 38654
rect 25332 38282 25360 38626
rect 25516 38418 25544 38830
rect 25504 38412 25556 38418
rect 25504 38354 25556 38360
rect 25320 38276 25372 38282
rect 25320 38218 25372 38224
rect 25228 37868 25280 37874
rect 25332 37856 25360 38218
rect 25280 37828 25360 37856
rect 25228 37810 25280 37816
rect 25332 36922 25360 37828
rect 25516 37806 25544 38354
rect 25504 37800 25556 37806
rect 25504 37742 25556 37748
rect 25516 37330 25544 37742
rect 25504 37324 25556 37330
rect 25504 37266 25556 37272
rect 25320 36916 25372 36922
rect 25320 36858 25372 36864
rect 25136 36100 25188 36106
rect 25136 36042 25188 36048
rect 25412 36100 25464 36106
rect 25412 36042 25464 36048
rect 25148 35766 25176 36042
rect 25424 35834 25452 36042
rect 25412 35828 25464 35834
rect 25412 35770 25464 35776
rect 24952 35760 25004 35766
rect 23754 35728 23810 35737
rect 23020 35692 23072 35698
rect 24952 35702 25004 35708
rect 25136 35760 25188 35766
rect 25136 35702 25188 35708
rect 23754 35663 23810 35672
rect 23020 35634 23072 35640
rect 22466 35456 22522 35465
rect 22466 35391 22522 35400
rect 22284 35284 22336 35290
rect 22204 35244 22284 35272
rect 22204 34610 22232 35244
rect 22284 35226 22336 35232
rect 22480 35086 22508 35391
rect 22468 35080 22520 35086
rect 22468 35022 22520 35028
rect 22560 35012 22612 35018
rect 22560 34954 22612 34960
rect 22928 35012 22980 35018
rect 22928 34954 22980 34960
rect 22572 34610 22600 34954
rect 22836 34944 22888 34950
rect 22836 34886 22888 34892
rect 22848 34610 22876 34886
rect 22192 34604 22244 34610
rect 22192 34546 22244 34552
rect 22560 34604 22612 34610
rect 22560 34546 22612 34552
rect 22836 34604 22888 34610
rect 22836 34546 22888 34552
rect 22560 33040 22612 33046
rect 22560 32982 22612 32988
rect 22190 32464 22246 32473
rect 22246 32408 22324 32416
rect 22190 32399 22192 32408
rect 22244 32388 22324 32408
rect 22192 32370 22244 32376
rect 22100 31884 22152 31890
rect 22100 31826 22152 31832
rect 22112 31414 22140 31826
rect 22192 31816 22244 31822
rect 22190 31784 22192 31793
rect 22244 31784 22246 31793
rect 22190 31719 22246 31728
rect 22192 31680 22244 31686
rect 22192 31622 22244 31628
rect 22100 31408 22152 31414
rect 22100 31350 22152 31356
rect 22204 31210 22232 31622
rect 22192 31204 22244 31210
rect 22192 31146 22244 31152
rect 22100 30592 22152 30598
rect 22100 30534 22152 30540
rect 22112 30258 22140 30534
rect 22100 30252 22152 30258
rect 22100 30194 22152 30200
rect 22112 28558 22140 30194
rect 22296 29889 22324 32388
rect 22572 32026 22600 32982
rect 22744 32428 22796 32434
rect 22744 32370 22796 32376
rect 22652 32360 22704 32366
rect 22756 32337 22784 32370
rect 22652 32302 22704 32308
rect 22742 32328 22798 32337
rect 22560 32020 22612 32026
rect 22560 31962 22612 31968
rect 22572 31278 22600 31962
rect 22664 31890 22692 32302
rect 22742 32263 22798 32272
rect 22744 32224 22796 32230
rect 22744 32166 22796 32172
rect 22652 31884 22704 31890
rect 22652 31826 22704 31832
rect 22376 31272 22428 31278
rect 22374 31240 22376 31249
rect 22560 31272 22612 31278
rect 22428 31240 22430 31249
rect 22560 31214 22612 31220
rect 22374 31175 22430 31184
rect 22376 31136 22428 31142
rect 22376 31078 22428 31084
rect 22388 30433 22416 31078
rect 22374 30424 22430 30433
rect 22374 30359 22430 30368
rect 22376 30320 22428 30326
rect 22376 30262 22428 30268
rect 22282 29880 22338 29889
rect 22282 29815 22338 29824
rect 22296 29646 22324 29815
rect 22284 29640 22336 29646
rect 22284 29582 22336 29588
rect 22388 29102 22416 30262
rect 22756 29730 22784 32166
rect 22836 31680 22888 31686
rect 22836 31622 22888 31628
rect 22848 30938 22876 31622
rect 22940 31482 22968 34954
rect 23768 34746 23796 35663
rect 23756 34740 23808 34746
rect 23756 34682 23808 34688
rect 24964 34610 24992 35702
rect 25700 34678 25728 41386
rect 26436 38418 26464 43101
rect 27080 39030 27108 43101
rect 27068 39024 27120 39030
rect 27068 38966 27120 38972
rect 27080 38418 27108 38966
rect 27436 38752 27488 38758
rect 27436 38694 27488 38700
rect 27448 38418 27476 38694
rect 26424 38412 26476 38418
rect 26424 38354 26476 38360
rect 27068 38412 27120 38418
rect 27068 38354 27120 38360
rect 27436 38412 27488 38418
rect 27436 38354 27488 38360
rect 26436 38010 26464 38354
rect 26424 38004 26476 38010
rect 26424 37946 26476 37952
rect 25964 37324 26016 37330
rect 25964 37266 26016 37272
rect 25976 36242 26004 37266
rect 27724 37262 27752 43101
rect 27712 37256 27764 37262
rect 27712 37198 27764 37204
rect 27724 36854 27752 37198
rect 27712 36848 27764 36854
rect 27712 36790 27764 36796
rect 28368 36242 28396 43101
rect 30944 41138 30972 43101
rect 35594 41372 35902 41381
rect 35594 41370 35600 41372
rect 35656 41370 35680 41372
rect 35736 41370 35760 41372
rect 35816 41370 35840 41372
rect 35896 41370 35902 41372
rect 35656 41318 35658 41370
rect 35838 41318 35840 41370
rect 35594 41316 35600 41318
rect 35656 41316 35680 41318
rect 35736 41316 35760 41318
rect 35816 41316 35840 41318
rect 35896 41316 35902 41318
rect 35594 41307 35902 41316
rect 30932 41132 30984 41138
rect 30932 41074 30984 41080
rect 31208 41064 31260 41070
rect 31208 41006 31260 41012
rect 28908 38344 28960 38350
rect 28908 38286 28960 38292
rect 25780 36236 25832 36242
rect 25780 36178 25832 36184
rect 25964 36236 26016 36242
rect 25964 36178 26016 36184
rect 27160 36236 27212 36242
rect 27160 36178 27212 36184
rect 28356 36236 28408 36242
rect 28356 36178 28408 36184
rect 25792 35612 25820 36178
rect 27172 35834 27200 36178
rect 27160 35828 27212 35834
rect 27160 35770 27212 35776
rect 25872 35624 25924 35630
rect 25792 35584 25872 35612
rect 25872 35566 25924 35572
rect 25688 34672 25740 34678
rect 25688 34614 25740 34620
rect 24952 34604 25004 34610
rect 24952 34546 25004 34552
rect 23848 34536 23900 34542
rect 23848 34478 23900 34484
rect 23860 34202 23888 34478
rect 23848 34196 23900 34202
rect 23848 34138 23900 34144
rect 25136 34060 25188 34066
rect 25136 34002 25188 34008
rect 24400 33312 24452 33318
rect 24400 33254 24452 33260
rect 24124 32904 24176 32910
rect 23846 32872 23902 32881
rect 23664 32836 23716 32842
rect 24124 32846 24176 32852
rect 23846 32807 23902 32816
rect 23664 32778 23716 32784
rect 23020 32428 23072 32434
rect 23020 32370 23072 32376
rect 23296 32428 23348 32434
rect 23296 32370 23348 32376
rect 23388 32428 23440 32434
rect 23388 32370 23440 32376
rect 23032 32026 23060 32370
rect 23020 32020 23072 32026
rect 23020 31962 23072 31968
rect 23020 31816 23072 31822
rect 23020 31758 23072 31764
rect 22928 31476 22980 31482
rect 22928 31418 22980 31424
rect 23032 31385 23060 31758
rect 23308 31686 23336 32370
rect 23204 31680 23256 31686
rect 23204 31622 23256 31628
rect 23296 31680 23348 31686
rect 23296 31622 23348 31628
rect 23018 31376 23074 31385
rect 22928 31340 22980 31346
rect 23018 31311 23074 31320
rect 23112 31340 23164 31346
rect 22928 31282 22980 31288
rect 23112 31282 23164 31288
rect 22836 30932 22888 30938
rect 22836 30874 22888 30880
rect 22940 30870 22968 31282
rect 23020 31136 23072 31142
rect 23020 31078 23072 31084
rect 22928 30864 22980 30870
rect 22928 30806 22980 30812
rect 22834 29880 22890 29889
rect 22834 29815 22890 29824
rect 22664 29702 22784 29730
rect 22664 29646 22692 29702
rect 22652 29640 22704 29646
rect 22744 29640 22796 29646
rect 22652 29582 22704 29588
rect 22742 29608 22744 29617
rect 22796 29608 22798 29617
rect 22560 29572 22612 29578
rect 22560 29514 22612 29520
rect 22468 29504 22520 29510
rect 22468 29446 22520 29452
rect 22376 29096 22428 29102
rect 22376 29038 22428 29044
rect 22284 29028 22336 29034
rect 22284 28970 22336 28976
rect 22100 28552 22152 28558
rect 22100 28494 22152 28500
rect 22100 28076 22152 28082
rect 22100 28018 22152 28024
rect 22112 26976 22140 28018
rect 22192 26988 22244 26994
rect 22112 26948 22192 26976
rect 22192 26930 22244 26936
rect 22204 26897 22232 26930
rect 22190 26888 22246 26897
rect 22190 26823 22246 26832
rect 22190 26616 22246 26625
rect 22190 26551 22246 26560
rect 22204 26382 22232 26551
rect 22192 26376 22244 26382
rect 22190 26344 22192 26353
rect 22244 26344 22246 26353
rect 22190 26279 22246 26288
rect 22296 25498 22324 28970
rect 22480 28558 22508 29446
rect 22572 29102 22600 29514
rect 22664 29238 22692 29582
rect 22742 29543 22798 29552
rect 22652 29232 22704 29238
rect 22652 29174 22704 29180
rect 22560 29096 22612 29102
rect 22560 29038 22612 29044
rect 22468 28552 22520 28558
rect 22468 28494 22520 28500
rect 22480 28082 22508 28494
rect 22468 28076 22520 28082
rect 22468 28018 22520 28024
rect 22466 26616 22522 26625
rect 22466 26551 22468 26560
rect 22520 26551 22522 26560
rect 22468 26522 22520 26528
rect 22376 26376 22428 26382
rect 22374 26344 22376 26353
rect 22428 26344 22430 26353
rect 22374 26279 22430 26288
rect 22284 25492 22336 25498
rect 22284 25434 22336 25440
rect 22192 24948 22244 24954
rect 22192 24890 22244 24896
rect 22100 24676 22152 24682
rect 22100 24618 22152 24624
rect 22112 24041 22140 24618
rect 22098 24032 22154 24041
rect 22098 23967 22154 23976
rect 22100 23588 22152 23594
rect 22100 23530 22152 23536
rect 22006 21992 22062 22001
rect 22006 21927 22062 21936
rect 21732 21888 21784 21894
rect 21732 21830 21784 21836
rect 21824 21548 21876 21554
rect 21824 21490 21876 21496
rect 21732 20868 21784 20874
rect 21732 20810 21784 20816
rect 21744 19961 21772 20810
rect 21836 20806 21864 21490
rect 21916 21072 21968 21078
rect 21916 21014 21968 21020
rect 21824 20800 21876 20806
rect 21824 20742 21876 20748
rect 21822 20632 21878 20641
rect 21928 20618 21956 21014
rect 22020 20806 22048 21927
rect 22112 21418 22140 23530
rect 22204 22778 22232 24890
rect 22296 24818 22324 25434
rect 22572 24954 22600 29038
rect 22664 28422 22692 29174
rect 22652 28416 22704 28422
rect 22652 28358 22704 28364
rect 22744 28076 22796 28082
rect 22848 28064 22876 29815
rect 22796 28036 22876 28064
rect 22744 28018 22796 28024
rect 22756 27946 22784 28018
rect 22744 27940 22796 27946
rect 22744 27882 22796 27888
rect 22756 26994 22784 27882
rect 22836 27532 22888 27538
rect 22836 27474 22888 27480
rect 22652 26988 22704 26994
rect 22652 26930 22704 26936
rect 22744 26988 22796 26994
rect 22744 26930 22796 26936
rect 22664 26761 22692 26930
rect 22744 26784 22796 26790
rect 22650 26752 22706 26761
rect 22744 26726 22796 26732
rect 22650 26687 22706 26696
rect 22664 26586 22692 26687
rect 22652 26580 22704 26586
rect 22652 26522 22704 26528
rect 22756 25158 22784 26726
rect 22848 26450 22876 27474
rect 22940 27112 22968 30806
rect 23032 29714 23060 31078
rect 23124 30258 23152 31282
rect 23216 31210 23244 31622
rect 23308 31346 23336 31622
rect 23296 31340 23348 31346
rect 23296 31282 23348 31288
rect 23204 31204 23256 31210
rect 23204 31146 23256 31152
rect 23216 30938 23244 31146
rect 23204 30932 23256 30938
rect 23204 30874 23256 30880
rect 23204 30728 23256 30734
rect 23204 30670 23256 30676
rect 23112 30252 23164 30258
rect 23112 30194 23164 30200
rect 23020 29708 23072 29714
rect 23020 29650 23072 29656
rect 23216 29594 23244 30670
rect 23308 30394 23336 31282
rect 23400 30598 23428 32370
rect 23572 31340 23624 31346
rect 23572 31282 23624 31288
rect 23584 30734 23612 31282
rect 23676 30938 23704 32778
rect 23756 32768 23808 32774
rect 23756 32710 23808 32716
rect 23768 32434 23796 32710
rect 23756 32428 23808 32434
rect 23756 32370 23808 32376
rect 23860 32366 23888 32807
rect 23848 32360 23900 32366
rect 23848 32302 23900 32308
rect 23756 31884 23808 31890
rect 23756 31826 23808 31832
rect 23768 31668 23796 31826
rect 23848 31816 23900 31822
rect 23900 31776 24072 31804
rect 23848 31758 23900 31764
rect 23768 31640 23980 31668
rect 23848 31476 23900 31482
rect 23848 31418 23900 31424
rect 23860 31278 23888 31418
rect 23848 31272 23900 31278
rect 23848 31214 23900 31220
rect 23860 30938 23888 31214
rect 23664 30932 23716 30938
rect 23664 30874 23716 30880
rect 23848 30932 23900 30938
rect 23848 30874 23900 30880
rect 23572 30728 23624 30734
rect 23492 30688 23572 30716
rect 23388 30592 23440 30598
rect 23388 30534 23440 30540
rect 23296 30388 23348 30394
rect 23296 30330 23348 30336
rect 23400 30258 23428 30534
rect 23388 30252 23440 30258
rect 23124 29566 23244 29594
rect 23308 30212 23388 30240
rect 23018 29472 23074 29481
rect 23018 29407 23074 29416
rect 23032 29170 23060 29407
rect 23020 29164 23072 29170
rect 23020 29106 23072 29112
rect 23020 28960 23072 28966
rect 23020 28902 23072 28908
rect 23032 28082 23060 28902
rect 23124 28422 23152 29566
rect 23308 28994 23336 30212
rect 23388 30194 23440 30200
rect 23388 30048 23440 30054
rect 23388 29990 23440 29996
rect 23400 29646 23428 29990
rect 23492 29782 23520 30688
rect 23572 30670 23624 30676
rect 23676 30258 23704 30874
rect 23756 30728 23808 30734
rect 23756 30670 23808 30676
rect 23664 30252 23716 30258
rect 23664 30194 23716 30200
rect 23570 29880 23626 29889
rect 23570 29815 23626 29824
rect 23480 29776 23532 29782
rect 23480 29718 23532 29724
rect 23388 29640 23440 29646
rect 23388 29582 23440 29588
rect 23492 29170 23520 29718
rect 23584 29646 23612 29815
rect 23572 29640 23624 29646
rect 23572 29582 23624 29588
rect 23572 29504 23624 29510
rect 23572 29446 23624 29452
rect 23584 29170 23612 29446
rect 23662 29336 23718 29345
rect 23662 29271 23718 29280
rect 23676 29238 23704 29271
rect 23664 29232 23716 29238
rect 23664 29174 23716 29180
rect 23480 29164 23532 29170
rect 23480 29106 23532 29112
rect 23572 29164 23624 29170
rect 23572 29106 23624 29112
rect 23216 28966 23336 28994
rect 23216 28937 23244 28966
rect 23480 28960 23532 28966
rect 23202 28928 23258 28937
rect 23480 28902 23532 28908
rect 23202 28863 23258 28872
rect 23112 28416 23164 28422
rect 23112 28358 23164 28364
rect 23020 28076 23072 28082
rect 23020 28018 23072 28024
rect 23216 27538 23244 28863
rect 23492 28558 23520 28902
rect 23584 28626 23612 29106
rect 23664 28960 23716 28966
rect 23664 28902 23716 28908
rect 23572 28620 23624 28626
rect 23572 28562 23624 28568
rect 23388 28552 23440 28558
rect 23388 28494 23440 28500
rect 23480 28552 23532 28558
rect 23480 28494 23532 28500
rect 23296 27872 23348 27878
rect 23296 27814 23348 27820
rect 23204 27532 23256 27538
rect 23204 27474 23256 27480
rect 22940 27084 23060 27112
rect 22928 26580 22980 26586
rect 22928 26522 22980 26528
rect 22836 26444 22888 26450
rect 22836 26386 22888 26392
rect 22836 26240 22888 26246
rect 22836 26182 22888 26188
rect 22744 25152 22796 25158
rect 22744 25094 22796 25100
rect 22560 24948 22612 24954
rect 22560 24890 22612 24896
rect 22284 24812 22336 24818
rect 22284 24754 22336 24760
rect 22376 24608 22428 24614
rect 22376 24550 22428 24556
rect 22284 23112 22336 23118
rect 22284 23054 22336 23060
rect 22192 22772 22244 22778
rect 22192 22714 22244 22720
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 22204 21418 22232 21626
rect 22100 21412 22152 21418
rect 22100 21354 22152 21360
rect 22192 21412 22244 21418
rect 22192 21354 22244 21360
rect 22008 20800 22060 20806
rect 22006 20768 22008 20777
rect 22060 20768 22062 20777
rect 22006 20703 22062 20712
rect 21928 20590 22048 20618
rect 21822 20567 21878 20576
rect 21730 19952 21786 19961
rect 21730 19887 21786 19896
rect 21836 19854 21864 20567
rect 22020 20534 22048 20590
rect 22008 20528 22060 20534
rect 22008 20470 22060 20476
rect 21732 19848 21784 19854
rect 21732 19790 21784 19796
rect 21824 19848 21876 19854
rect 21824 19790 21876 19796
rect 21640 19508 21692 19514
rect 21640 19450 21692 19456
rect 21640 19304 21692 19310
rect 21744 19281 21772 19790
rect 21824 19508 21876 19514
rect 21824 19450 21876 19456
rect 21916 19508 21968 19514
rect 21916 19450 21968 19456
rect 21640 19246 21692 19252
rect 21730 19272 21786 19281
rect 21652 18970 21680 19246
rect 21836 19242 21864 19450
rect 21928 19417 21956 19450
rect 21914 19408 21970 19417
rect 21914 19343 21970 19352
rect 21730 19207 21786 19216
rect 21824 19236 21876 19242
rect 21824 19178 21876 19184
rect 21640 18964 21692 18970
rect 21640 18906 21692 18912
rect 21652 18766 21680 18906
rect 22020 18850 22048 20470
rect 22296 20466 22324 23054
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 22100 19984 22152 19990
rect 22100 19926 22152 19932
rect 21928 18822 22048 18850
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 21824 18760 21876 18766
rect 21824 18702 21876 18708
rect 21640 18624 21692 18630
rect 21836 18601 21864 18702
rect 21640 18566 21692 18572
rect 21822 18592 21878 18601
rect 21548 15700 21600 15706
rect 21548 15642 21600 15648
rect 21548 15088 21600 15094
rect 21548 15030 21600 15036
rect 21560 13326 21588 15030
rect 21652 13376 21680 18566
rect 21822 18527 21878 18536
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21836 17678 21864 18226
rect 21824 17672 21876 17678
rect 21824 17614 21876 17620
rect 21836 16590 21864 17614
rect 21824 16584 21876 16590
rect 21824 16526 21876 16532
rect 21732 15360 21784 15366
rect 21732 15302 21784 15308
rect 21744 14550 21772 15302
rect 21732 14544 21784 14550
rect 21732 14486 21784 14492
rect 21732 14408 21784 14414
rect 21732 14350 21784 14356
rect 21744 14074 21772 14350
rect 21732 14068 21784 14074
rect 21732 14010 21784 14016
rect 21744 13530 21772 14010
rect 21732 13524 21784 13530
rect 21732 13466 21784 13472
rect 21732 13388 21784 13394
rect 21652 13348 21732 13376
rect 21732 13330 21784 13336
rect 21548 13320 21600 13326
rect 21600 13280 21680 13308
rect 21548 13262 21600 13268
rect 21548 13184 21600 13190
rect 21548 13126 21600 13132
rect 21560 12646 21588 13126
rect 21652 12986 21680 13280
rect 21640 12980 21692 12986
rect 21640 12922 21692 12928
rect 21836 12866 21864 16526
rect 21652 12838 21864 12866
rect 21548 12640 21600 12646
rect 21548 12582 21600 12588
rect 21548 11756 21600 11762
rect 21548 11698 21600 11704
rect 21456 11076 21508 11082
rect 21456 11018 21508 11024
rect 21362 10704 21418 10713
rect 21272 10668 21324 10674
rect 21560 10674 21588 11698
rect 21362 10639 21418 10648
rect 21548 10668 21600 10674
rect 21272 10610 21324 10616
rect 21180 9512 21232 9518
rect 21180 9454 21232 9460
rect 21192 9217 21220 9454
rect 21178 9208 21234 9217
rect 21178 9143 21234 9152
rect 21180 8492 21232 8498
rect 21180 8434 21232 8440
rect 20916 7500 21128 7528
rect 20812 7472 20864 7478
rect 20812 7414 20864 7420
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20916 7342 20944 7500
rect 21086 7440 21142 7449
rect 21086 7375 21088 7384
rect 21140 7375 21142 7384
rect 21088 7346 21140 7352
rect 20904 7336 20956 7342
rect 20904 7278 20956 7284
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20536 6996 20588 7002
rect 20536 6938 20588 6944
rect 20628 6996 20680 7002
rect 20628 6938 20680 6944
rect 19616 6928 19668 6934
rect 19616 6870 19668 6876
rect 20548 6798 20576 6938
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 19340 6384 19392 6390
rect 20260 6384 20312 6390
rect 19340 6326 19392 6332
rect 20180 6344 20260 6372
rect 19524 6112 19576 6118
rect 19524 6054 19576 6060
rect 19340 5840 19392 5846
rect 19340 5782 19392 5788
rect 19156 5704 19208 5710
rect 18840 5664 18920 5692
rect 19076 5664 19156 5692
rect 18788 5646 18840 5652
rect 18892 4146 18920 5664
rect 19156 5646 19208 5652
rect 19248 5568 19300 5574
rect 19248 5510 19300 5516
rect 18972 5160 19024 5166
rect 18972 5102 19024 5108
rect 19260 5114 19288 5510
rect 19352 5234 19380 5782
rect 19536 5710 19564 6054
rect 19982 5944 20038 5953
rect 19982 5879 19984 5888
rect 20036 5879 20038 5888
rect 19984 5850 20036 5856
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19892 5704 19944 5710
rect 19892 5646 19944 5652
rect 20076 5704 20128 5710
rect 20076 5646 20128 5652
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 18984 4826 19012 5102
rect 19260 5098 19380 5114
rect 19260 5092 19392 5098
rect 19260 5086 19340 5092
rect 19340 5034 19392 5040
rect 18972 4820 19024 4826
rect 18972 4762 19024 4768
rect 19352 4214 19380 5034
rect 19340 4208 19392 4214
rect 19340 4150 19392 4156
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18880 4140 18932 4146
rect 18880 4082 18932 4088
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 18604 4072 18656 4078
rect 18604 4014 18656 4020
rect 19444 4010 19472 5646
rect 19524 5024 19576 5030
rect 19524 4966 19576 4972
rect 19536 4690 19564 4966
rect 19708 4820 19760 4826
rect 19708 4762 19760 4768
rect 19524 4684 19576 4690
rect 19524 4626 19576 4632
rect 19720 4146 19748 4762
rect 19904 4146 19932 5646
rect 20088 5302 20116 5646
rect 20076 5296 20128 5302
rect 20076 5238 20128 5244
rect 20088 5098 20116 5238
rect 20076 5092 20128 5098
rect 20076 5034 20128 5040
rect 20088 4690 20116 5034
rect 20076 4684 20128 4690
rect 20076 4626 20128 4632
rect 20180 4554 20208 6344
rect 20260 6326 20312 6332
rect 20444 6248 20496 6254
rect 20444 6190 20496 6196
rect 20456 5914 20484 6190
rect 20444 5908 20496 5914
rect 20444 5850 20496 5856
rect 20732 5846 20760 7142
rect 20720 5840 20772 5846
rect 20720 5782 20772 5788
rect 20536 5704 20588 5710
rect 20536 5646 20588 5652
rect 20548 4826 20576 5646
rect 20628 5228 20680 5234
rect 20628 5170 20680 5176
rect 20640 5030 20668 5170
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 20536 4820 20588 4826
rect 20536 4762 20588 4768
rect 20640 4758 20668 4966
rect 20628 4752 20680 4758
rect 20628 4694 20680 4700
rect 20168 4548 20220 4554
rect 20168 4490 20220 4496
rect 20180 4214 20208 4490
rect 20168 4208 20220 4214
rect 20168 4150 20220 4156
rect 20732 4146 20760 5782
rect 20916 5114 20944 7278
rect 20824 5086 20944 5114
rect 19708 4140 19760 4146
rect 19708 4082 19760 4088
rect 19892 4140 19944 4146
rect 19892 4082 19944 4088
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 19432 4004 19484 4010
rect 19432 3946 19484 3952
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18800 3534 18828 3878
rect 20088 3738 20116 4082
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 18788 3528 18840 3534
rect 18788 3470 18840 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 18800 3126 18828 3470
rect 18788 3120 18840 3126
rect 18788 3062 18840 3068
rect 18064 2746 18184 2774
rect 17960 2372 18012 2378
rect 17960 2314 18012 2320
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 16132 800 16160 2246
rect 16776 800 16804 2246
rect 18064 800 18092 2746
rect 19260 2650 19288 3470
rect 20824 2990 20852 5086
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20916 4282 20944 4966
rect 20904 4276 20956 4282
rect 20904 4218 20956 4224
rect 21192 4078 21220 8434
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21284 7342 21312 7482
rect 21272 7336 21324 7342
rect 21272 7278 21324 7284
rect 21284 6458 21312 7278
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 21284 6118 21312 6394
rect 21272 6112 21324 6118
rect 21272 6054 21324 6060
rect 21284 5710 21312 6054
rect 21376 5846 21404 10639
rect 21548 10610 21600 10616
rect 21652 8294 21680 12838
rect 21928 12764 21956 18822
rect 22008 18760 22060 18766
rect 22112 18748 22140 19926
rect 22296 19854 22324 20402
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 22388 19802 22416 24550
rect 22558 23896 22614 23905
rect 22558 23831 22614 23840
rect 22572 23730 22600 23831
rect 22742 23760 22798 23769
rect 22560 23724 22612 23730
rect 22742 23695 22744 23704
rect 22560 23666 22612 23672
rect 22796 23695 22798 23704
rect 22744 23666 22796 23672
rect 22848 23202 22876 26182
rect 22940 24052 22968 26522
rect 23032 26353 23060 27084
rect 23308 26994 23336 27814
rect 23296 26988 23348 26994
rect 23296 26930 23348 26936
rect 23400 26874 23428 28494
rect 23676 28014 23704 28902
rect 23768 28558 23796 30670
rect 23848 30592 23900 30598
rect 23848 30534 23900 30540
rect 23860 29782 23888 30534
rect 23848 29776 23900 29782
rect 23848 29718 23900 29724
rect 23848 29640 23900 29646
rect 23848 29582 23900 29588
rect 23860 29170 23888 29582
rect 23848 29164 23900 29170
rect 23848 29106 23900 29112
rect 23848 29028 23900 29034
rect 23848 28970 23900 28976
rect 23860 28937 23888 28970
rect 23846 28928 23902 28937
rect 23846 28863 23902 28872
rect 23756 28552 23808 28558
rect 23756 28494 23808 28500
rect 23756 28416 23808 28422
rect 23756 28358 23808 28364
rect 23768 28014 23796 28358
rect 23664 28008 23716 28014
rect 23664 27950 23716 27956
rect 23756 28008 23808 28014
rect 23756 27950 23808 27956
rect 23204 26852 23256 26858
rect 23204 26794 23256 26800
rect 23308 26846 23428 26874
rect 23480 26920 23532 26926
rect 23480 26862 23532 26868
rect 23018 26344 23074 26353
rect 23018 26279 23074 26288
rect 23112 26240 23164 26246
rect 23112 26182 23164 26188
rect 23020 25356 23072 25362
rect 23020 25298 23072 25304
rect 23032 24206 23060 25298
rect 23124 25226 23152 26182
rect 23216 25838 23244 26794
rect 23204 25832 23256 25838
rect 23204 25774 23256 25780
rect 23308 25673 23336 26846
rect 23492 26364 23520 26862
rect 23572 26376 23624 26382
rect 23492 26336 23572 26364
rect 23388 26308 23440 26314
rect 23388 26250 23440 26256
rect 23294 25664 23350 25673
rect 23294 25599 23350 25608
rect 23112 25220 23164 25226
rect 23112 25162 23164 25168
rect 23020 24200 23072 24206
rect 23020 24142 23072 24148
rect 22940 24024 23244 24052
rect 23018 23896 23074 23905
rect 23018 23831 23074 23840
rect 22756 23174 22876 23202
rect 22468 22024 22520 22030
rect 22466 21992 22468 22001
rect 22520 21992 22522 22001
rect 22466 21927 22522 21936
rect 22756 19854 22784 23174
rect 22836 23112 22888 23118
rect 22836 23054 22888 23060
rect 22848 20466 22876 23054
rect 22928 22772 22980 22778
rect 22928 22714 22980 22720
rect 22940 22030 22968 22714
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 22836 20460 22888 20466
rect 22836 20402 22888 20408
rect 22848 20058 22876 20402
rect 22836 20052 22888 20058
rect 22836 19994 22888 20000
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 22744 19848 22796 19854
rect 22192 19780 22244 19786
rect 22388 19774 22600 19802
rect 22744 19790 22796 19796
rect 22192 19722 22244 19728
rect 22204 19378 22232 19722
rect 22376 19712 22428 19718
rect 22376 19654 22428 19660
rect 22388 19514 22416 19654
rect 22376 19508 22428 19514
rect 22376 19450 22428 19456
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22060 18720 22140 18748
rect 22008 18702 22060 18708
rect 22192 18624 22244 18630
rect 22192 18566 22244 18572
rect 22204 18290 22232 18566
rect 22284 18352 22336 18358
rect 22284 18294 22336 18300
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 22192 17808 22244 17814
rect 22192 17750 22244 17756
rect 22204 16658 22232 17750
rect 22296 16674 22324 18294
rect 22388 18290 22416 19450
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22376 18080 22428 18086
rect 22376 18022 22428 18028
rect 22388 17678 22416 18022
rect 22376 17672 22428 17678
rect 22376 17614 22428 17620
rect 22192 16652 22244 16658
rect 22296 16646 22416 16674
rect 22192 16594 22244 16600
rect 22284 16516 22336 16522
rect 22284 16458 22336 16464
rect 22296 16182 22324 16458
rect 22284 16176 22336 16182
rect 22284 16118 22336 16124
rect 22006 15872 22062 15881
rect 22006 15807 22062 15816
rect 22020 15706 22048 15807
rect 22008 15700 22060 15706
rect 22008 15642 22060 15648
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22098 15600 22154 15609
rect 22008 15564 22060 15570
rect 22098 15535 22100 15544
rect 22008 15506 22060 15512
rect 22152 15535 22154 15544
rect 22100 15506 22152 15512
rect 22020 14006 22048 15506
rect 22204 15502 22232 15642
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 22204 14770 22232 15438
rect 22296 15026 22324 16118
rect 22388 15348 22416 16646
rect 22572 16454 22600 19774
rect 22848 19378 22876 19858
rect 22928 19440 22980 19446
rect 22928 19382 22980 19388
rect 22836 19372 22888 19378
rect 22836 19314 22888 19320
rect 22940 18873 22968 19382
rect 22926 18864 22982 18873
rect 22926 18799 22982 18808
rect 22652 17672 22704 17678
rect 22652 17614 22704 17620
rect 22664 16833 22692 17614
rect 22926 17368 22982 17377
rect 22926 17303 22982 17312
rect 22940 17134 22968 17303
rect 22928 17128 22980 17134
rect 22928 17070 22980 17076
rect 22836 16992 22888 16998
rect 22836 16934 22888 16940
rect 22650 16824 22706 16833
rect 22650 16759 22706 16768
rect 22664 16726 22692 16759
rect 22652 16720 22704 16726
rect 22652 16662 22704 16668
rect 22652 16584 22704 16590
rect 22848 16538 22876 16934
rect 22926 16824 22982 16833
rect 22926 16759 22928 16768
rect 22980 16759 22982 16768
rect 22928 16730 22980 16736
rect 22928 16652 22980 16658
rect 22928 16594 22980 16600
rect 22704 16532 22876 16538
rect 22652 16526 22876 16532
rect 22664 16510 22876 16526
rect 22560 16448 22612 16454
rect 22560 16390 22612 16396
rect 22468 15496 22520 15502
rect 22520 15456 22692 15484
rect 22468 15438 22520 15444
rect 22664 15366 22692 15456
rect 22652 15360 22704 15366
rect 22388 15320 22600 15348
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22204 14742 22324 14770
rect 22190 14648 22246 14657
rect 22190 14583 22192 14592
rect 22244 14583 22246 14592
rect 22192 14554 22244 14560
rect 22100 14408 22152 14414
rect 22100 14350 22152 14356
rect 22008 14000 22060 14006
rect 22008 13942 22060 13948
rect 22112 13870 22140 14350
rect 22296 14074 22324 14742
rect 22468 14340 22520 14346
rect 22468 14282 22520 14288
rect 22374 14240 22430 14249
rect 22374 14175 22430 14184
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 22388 13462 22416 14175
rect 22376 13456 22428 13462
rect 22376 13398 22428 13404
rect 22100 13388 22152 13394
rect 22100 13330 22152 13336
rect 22112 13297 22140 13330
rect 22376 13320 22428 13326
rect 22098 13288 22154 13297
rect 22376 13262 22428 13268
rect 22098 13223 22154 13232
rect 22006 13152 22062 13161
rect 22006 13087 22062 13096
rect 21836 12736 21956 12764
rect 21732 12640 21784 12646
rect 21732 12582 21784 12588
rect 21744 12442 21772 12582
rect 21732 12436 21784 12442
rect 21732 12378 21784 12384
rect 21836 10810 21864 12736
rect 22020 12050 22048 13087
rect 22112 12850 22140 13223
rect 22388 12850 22416 13262
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 22192 12776 22244 12782
rect 22192 12718 22244 12724
rect 22204 12102 22232 12718
rect 22376 12232 22428 12238
rect 22376 12174 22428 12180
rect 22192 12096 22244 12102
rect 22020 12022 22140 12050
rect 22192 12038 22244 12044
rect 22006 11928 22062 11937
rect 22006 11863 22062 11872
rect 22020 11830 22048 11863
rect 22008 11824 22060 11830
rect 22008 11766 22060 11772
rect 22112 11694 22140 12022
rect 22282 11792 22338 11801
rect 22282 11727 22338 11736
rect 22100 11688 22152 11694
rect 22100 11630 22152 11636
rect 22192 11348 22244 11354
rect 22192 11290 22244 11296
rect 21916 11008 21968 11014
rect 21916 10950 21968 10956
rect 21824 10804 21876 10810
rect 21824 10746 21876 10752
rect 21822 10704 21878 10713
rect 21822 10639 21824 10648
rect 21876 10639 21878 10648
rect 21824 10610 21876 10616
rect 21928 10606 21956 10950
rect 22100 10736 22152 10742
rect 22020 10684 22100 10690
rect 22020 10678 22152 10684
rect 22020 10662 22140 10678
rect 21732 10600 21784 10606
rect 21732 10542 21784 10548
rect 21916 10600 21968 10606
rect 21916 10542 21968 10548
rect 21744 8430 21772 10542
rect 22020 10470 22048 10662
rect 21824 10464 21876 10470
rect 21824 10406 21876 10412
rect 22008 10464 22060 10470
rect 22008 10406 22060 10412
rect 21732 8424 21784 8430
rect 21732 8366 21784 8372
rect 21836 8294 21864 10406
rect 22204 9518 22232 11290
rect 22296 11218 22324 11727
rect 22284 11212 22336 11218
rect 22284 11154 22336 11160
rect 22388 10656 22416 12174
rect 22480 11354 22508 14282
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 22468 11144 22520 11150
rect 22468 11086 22520 11092
rect 22480 10810 22508 11086
rect 22468 10804 22520 10810
rect 22468 10746 22520 10752
rect 22468 10668 22520 10674
rect 22388 10628 22468 10656
rect 22468 10610 22520 10616
rect 22376 10464 22428 10470
rect 22376 10406 22428 10412
rect 22388 9722 22416 10406
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 22284 9580 22336 9586
rect 22284 9522 22336 9528
rect 22008 9512 22060 9518
rect 22008 9454 22060 9460
rect 22192 9512 22244 9518
rect 22192 9454 22244 9460
rect 21640 8288 21692 8294
rect 21640 8230 21692 8236
rect 21824 8288 21876 8294
rect 21824 8230 21876 8236
rect 21836 7954 21864 8230
rect 21824 7948 21876 7954
rect 21824 7890 21876 7896
rect 22020 7546 22048 9454
rect 22204 9178 22232 9454
rect 22192 9172 22244 9178
rect 22192 9114 22244 9120
rect 22296 9058 22324 9522
rect 22204 9030 22324 9058
rect 22204 8401 22232 9030
rect 22284 8560 22336 8566
rect 22284 8502 22336 8508
rect 22190 8392 22246 8401
rect 22190 8327 22192 8336
rect 22244 8327 22246 8336
rect 22192 8298 22244 8304
rect 22296 7886 22324 8502
rect 22376 8016 22428 8022
rect 22376 7958 22428 7964
rect 22100 7880 22152 7886
rect 22100 7822 22152 7828
rect 22284 7880 22336 7886
rect 22284 7822 22336 7828
rect 22008 7540 22060 7546
rect 22112 7528 22140 7822
rect 22192 7540 22244 7546
rect 22112 7500 22192 7528
rect 22008 7482 22060 7488
rect 22192 7482 22244 7488
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21468 6934 21496 7142
rect 22296 6934 22324 7822
rect 22388 7478 22416 7958
rect 22480 7886 22508 10610
rect 22572 9654 22600 15320
rect 22652 15302 22704 15308
rect 22664 15162 22692 15302
rect 22652 15156 22704 15162
rect 22652 15098 22704 15104
rect 22652 14952 22704 14958
rect 22652 14894 22704 14900
rect 22664 14618 22692 14894
rect 22652 14612 22704 14618
rect 22652 14554 22704 14560
rect 22756 14498 22784 16510
rect 22836 15564 22888 15570
rect 22836 15506 22888 15512
rect 22848 15026 22876 15506
rect 22836 15020 22888 15026
rect 22836 14962 22888 14968
rect 22940 14822 22968 16594
rect 22928 14816 22980 14822
rect 22928 14758 22980 14764
rect 22664 14470 22784 14498
rect 22836 14544 22888 14550
rect 22836 14486 22888 14492
rect 22560 9648 22612 9654
rect 22560 9590 22612 9596
rect 22664 9466 22692 14470
rect 22744 14408 22796 14414
rect 22744 14350 22796 14356
rect 22756 13462 22784 14350
rect 22848 13802 22876 14486
rect 23032 14396 23060 23831
rect 23112 23724 23164 23730
rect 23112 23666 23164 23672
rect 23124 23118 23152 23666
rect 23112 23112 23164 23118
rect 23112 23054 23164 23060
rect 23216 21078 23244 24024
rect 23400 23497 23428 26250
rect 23492 24290 23520 26336
rect 23572 26318 23624 26324
rect 23572 25696 23624 25702
rect 23572 25638 23624 25644
rect 23584 25294 23612 25638
rect 23664 25356 23716 25362
rect 23664 25298 23716 25304
rect 23572 25288 23624 25294
rect 23572 25230 23624 25236
rect 23676 24857 23704 25298
rect 23952 24954 23980 31640
rect 24044 29646 24072 31776
rect 24136 31754 24164 32846
rect 24216 32224 24268 32230
rect 24216 32166 24268 32172
rect 24124 31748 24176 31754
rect 24124 31690 24176 31696
rect 24228 31686 24256 32166
rect 24216 31680 24268 31686
rect 24216 31622 24268 31628
rect 24228 30326 24256 31622
rect 24308 31136 24360 31142
rect 24308 31078 24360 31084
rect 24320 30841 24348 31078
rect 24306 30832 24362 30841
rect 24306 30767 24362 30776
rect 24216 30320 24268 30326
rect 24216 30262 24268 30268
rect 24216 30048 24268 30054
rect 24216 29990 24268 29996
rect 24124 29776 24176 29782
rect 24124 29718 24176 29724
rect 24032 29640 24084 29646
rect 24032 29582 24084 29588
rect 24044 29481 24072 29582
rect 24030 29472 24086 29481
rect 24030 29407 24086 29416
rect 24044 29170 24072 29407
rect 24032 29164 24084 29170
rect 24032 29106 24084 29112
rect 24032 28756 24084 28762
rect 24032 28698 24084 28704
rect 24044 26586 24072 28698
rect 24136 27130 24164 29718
rect 24228 29714 24256 29990
rect 24216 29708 24268 29714
rect 24216 29650 24268 29656
rect 24216 29504 24268 29510
rect 24216 29446 24268 29452
rect 24306 29472 24362 29481
rect 24228 28529 24256 29446
rect 24306 29407 24362 29416
rect 24320 28642 24348 29407
rect 24412 28762 24440 33254
rect 24676 32904 24728 32910
rect 24676 32846 24728 32852
rect 24688 32502 24716 32846
rect 25044 32768 25096 32774
rect 25044 32710 25096 32716
rect 24676 32496 24728 32502
rect 24676 32438 24728 32444
rect 25056 32434 25084 32710
rect 25148 32502 25176 34002
rect 25700 33998 25728 34614
rect 25884 34066 25912 35566
rect 28920 34610 28948 38286
rect 30472 36100 30524 36106
rect 30472 36042 30524 36048
rect 28264 34604 28316 34610
rect 28264 34546 28316 34552
rect 28908 34604 28960 34610
rect 28908 34546 28960 34552
rect 25872 34060 25924 34066
rect 25872 34002 25924 34008
rect 25688 33992 25740 33998
rect 25688 33934 25740 33940
rect 28276 33912 28304 34546
rect 28356 34536 28408 34542
rect 28356 34478 28408 34484
rect 28368 34202 28396 34478
rect 28356 34196 28408 34202
rect 28408 34156 28672 34184
rect 28356 34138 28408 34144
rect 28356 33924 28408 33930
rect 28276 33884 28356 33912
rect 28356 33866 28408 33872
rect 28368 33590 28396 33866
rect 28356 33584 28408 33590
rect 28356 33526 28408 33532
rect 28080 33312 28132 33318
rect 28080 33254 28132 33260
rect 26792 32972 26844 32978
rect 26792 32914 26844 32920
rect 25780 32904 25832 32910
rect 25516 32864 25780 32892
rect 25136 32496 25188 32502
rect 25136 32438 25188 32444
rect 24860 32428 24912 32434
rect 24860 32370 24912 32376
rect 24952 32428 25004 32434
rect 24952 32370 25004 32376
rect 25044 32428 25096 32434
rect 25044 32370 25096 32376
rect 25320 32428 25372 32434
rect 25320 32370 25372 32376
rect 25412 32428 25464 32434
rect 25412 32370 25464 32376
rect 24492 32360 24544 32366
rect 24492 32302 24544 32308
rect 24504 32065 24532 32302
rect 24490 32056 24546 32065
rect 24490 31991 24546 32000
rect 24872 31890 24900 32370
rect 24964 32337 24992 32370
rect 24950 32328 25006 32337
rect 24950 32263 25006 32272
rect 24860 31884 24912 31890
rect 24860 31826 24912 31832
rect 24584 31748 24636 31754
rect 24584 31690 24636 31696
rect 24492 30184 24544 30190
rect 24492 30126 24544 30132
rect 24504 29170 24532 30126
rect 24492 29164 24544 29170
rect 24492 29106 24544 29112
rect 24490 29064 24546 29073
rect 24490 28999 24546 29008
rect 24504 28966 24532 28999
rect 24492 28960 24544 28966
rect 24492 28902 24544 28908
rect 24400 28756 24452 28762
rect 24400 28698 24452 28704
rect 24320 28614 24440 28642
rect 24214 28520 24270 28529
rect 24214 28455 24216 28464
rect 24268 28455 24270 28464
rect 24216 28426 24268 28432
rect 24228 27878 24256 28426
rect 24216 27872 24268 27878
rect 24216 27814 24268 27820
rect 24308 27328 24360 27334
rect 24308 27270 24360 27276
rect 24124 27124 24176 27130
rect 24124 27066 24176 27072
rect 24124 26988 24176 26994
rect 24124 26930 24176 26936
rect 24032 26580 24084 26586
rect 24032 26522 24084 26528
rect 24032 26240 24084 26246
rect 24032 26182 24084 26188
rect 23940 24948 23992 24954
rect 23940 24890 23992 24896
rect 23662 24848 23718 24857
rect 23662 24783 23718 24792
rect 23664 24744 23716 24750
rect 24044 24698 24072 26182
rect 23664 24686 23716 24692
rect 23492 24262 23612 24290
rect 23480 24200 23532 24206
rect 23480 24142 23532 24148
rect 23492 24070 23520 24142
rect 23480 24064 23532 24070
rect 23480 24006 23532 24012
rect 23478 23896 23534 23905
rect 23478 23831 23534 23840
rect 23492 23662 23520 23831
rect 23480 23656 23532 23662
rect 23480 23598 23532 23604
rect 23386 23488 23442 23497
rect 23386 23423 23442 23432
rect 23296 23316 23348 23322
rect 23296 23258 23348 23264
rect 23308 22506 23336 23258
rect 23296 22500 23348 22506
rect 23296 22442 23348 22448
rect 23204 21072 23256 21078
rect 23204 21014 23256 21020
rect 23112 20528 23164 20534
rect 23112 20470 23164 20476
rect 23124 20233 23152 20470
rect 23216 20262 23244 21014
rect 23204 20256 23256 20262
rect 23110 20224 23166 20233
rect 23204 20198 23256 20204
rect 23110 20159 23166 20168
rect 23112 20052 23164 20058
rect 23112 19994 23164 20000
rect 23124 19854 23152 19994
rect 23204 19984 23256 19990
rect 23202 19952 23204 19961
rect 23256 19952 23258 19961
rect 23202 19887 23258 19896
rect 23112 19848 23164 19854
rect 23112 19790 23164 19796
rect 23110 19544 23166 19553
rect 23308 19514 23336 22442
rect 23480 22160 23532 22166
rect 23480 22102 23532 22108
rect 23388 21616 23440 21622
rect 23386 21584 23388 21593
rect 23440 21584 23442 21593
rect 23386 21519 23442 21528
rect 23388 20392 23440 20398
rect 23388 20334 23440 20340
rect 23400 19922 23428 20334
rect 23492 20330 23520 22102
rect 23584 20942 23612 24262
rect 23676 24206 23704 24686
rect 23952 24670 24072 24698
rect 23848 24404 23900 24410
rect 23768 24364 23848 24392
rect 23664 24200 23716 24206
rect 23664 24142 23716 24148
rect 23664 24064 23716 24070
rect 23664 24006 23716 24012
rect 23572 20936 23624 20942
rect 23572 20878 23624 20884
rect 23676 20448 23704 24006
rect 23768 23866 23796 24364
rect 23848 24346 23900 24352
rect 23848 24200 23900 24206
rect 23848 24142 23900 24148
rect 23756 23860 23808 23866
rect 23756 23802 23808 23808
rect 23756 23724 23808 23730
rect 23756 23666 23808 23672
rect 23768 22642 23796 23666
rect 23860 23594 23888 24142
rect 23848 23588 23900 23594
rect 23848 23530 23900 23536
rect 23756 22636 23808 22642
rect 23756 22578 23808 22584
rect 23768 22080 23796 22578
rect 23952 22273 23980 24670
rect 24136 24410 24164 26930
rect 24216 26784 24268 26790
rect 24216 26726 24268 26732
rect 24228 26382 24256 26726
rect 24216 26376 24268 26382
rect 24216 26318 24268 26324
rect 24216 26036 24268 26042
rect 24216 25978 24268 25984
rect 24228 25226 24256 25978
rect 24216 25220 24268 25226
rect 24216 25162 24268 25168
rect 24124 24404 24176 24410
rect 24124 24346 24176 24352
rect 24320 24290 24348 27270
rect 24412 26246 24440 28614
rect 24492 27600 24544 27606
rect 24492 27542 24544 27548
rect 24504 26382 24532 27542
rect 24596 27334 24624 31690
rect 24964 31414 24992 32263
rect 24952 31408 25004 31414
rect 24952 31350 25004 31356
rect 24952 31272 25004 31278
rect 24952 31214 25004 31220
rect 24676 30184 24728 30190
rect 24676 30126 24728 30132
rect 24688 29594 24716 30126
rect 24688 29566 24808 29594
rect 24676 29504 24728 29510
rect 24674 29472 24676 29481
rect 24728 29472 24730 29481
rect 24674 29407 24730 29416
rect 24780 29170 24808 29566
rect 24860 29572 24912 29578
rect 24860 29514 24912 29520
rect 24768 29164 24820 29170
rect 24768 29106 24820 29112
rect 24872 29034 24900 29514
rect 24860 29028 24912 29034
rect 24860 28970 24912 28976
rect 24676 28688 24728 28694
rect 24728 28636 24900 28642
rect 24676 28630 24900 28636
rect 24688 28614 24900 28630
rect 24676 28552 24728 28558
rect 24676 28494 24728 28500
rect 24768 28552 24820 28558
rect 24768 28494 24820 28500
rect 24584 27328 24636 27334
rect 24584 27270 24636 27276
rect 24688 26926 24716 28494
rect 24780 28150 24808 28494
rect 24768 28144 24820 28150
rect 24768 28086 24820 28092
rect 24872 27402 24900 28614
rect 24860 27396 24912 27402
rect 24860 27338 24912 27344
rect 24584 26920 24636 26926
rect 24584 26862 24636 26868
rect 24676 26920 24728 26926
rect 24676 26862 24728 26868
rect 24596 26568 24624 26862
rect 24676 26580 24728 26586
rect 24596 26540 24676 26568
rect 24676 26522 24728 26528
rect 24492 26376 24544 26382
rect 24492 26318 24544 26324
rect 24676 26376 24728 26382
rect 24676 26318 24728 26324
rect 24768 26376 24820 26382
rect 24768 26318 24820 26324
rect 24400 26240 24452 26246
rect 24400 26182 24452 26188
rect 24584 26240 24636 26246
rect 24584 26182 24636 26188
rect 24400 25356 24452 25362
rect 24400 25298 24452 25304
rect 24412 24886 24440 25298
rect 24596 25294 24624 26182
rect 24688 25906 24716 26318
rect 24676 25900 24728 25906
rect 24676 25842 24728 25848
rect 24780 25498 24808 26318
rect 24858 25528 24914 25537
rect 24768 25492 24820 25498
rect 24858 25463 24860 25472
rect 24768 25434 24820 25440
rect 24912 25463 24914 25472
rect 24860 25434 24912 25440
rect 24584 25288 24636 25294
rect 24584 25230 24636 25236
rect 24492 25220 24544 25226
rect 24492 25162 24544 25168
rect 24400 24880 24452 24886
rect 24400 24822 24452 24828
rect 24504 24818 24532 25162
rect 24492 24812 24544 24818
rect 24492 24754 24544 24760
rect 24136 24262 24348 24290
rect 24400 24268 24452 24274
rect 24030 24032 24086 24041
rect 24030 23967 24086 23976
rect 24044 23730 24072 23967
rect 24032 23724 24084 23730
rect 24032 23666 24084 23672
rect 24032 23180 24084 23186
rect 24032 23122 24084 23128
rect 24044 22642 24072 23122
rect 24136 22642 24164 24262
rect 24400 24210 24452 24216
rect 24216 24132 24268 24138
rect 24216 24074 24268 24080
rect 24228 24041 24256 24074
rect 24214 24032 24270 24041
rect 24214 23967 24270 23976
rect 24216 23656 24268 23662
rect 24216 23598 24268 23604
rect 24032 22636 24084 22642
rect 24032 22578 24084 22584
rect 24124 22636 24176 22642
rect 24124 22578 24176 22584
rect 24044 22545 24072 22578
rect 24030 22536 24086 22545
rect 24030 22471 24086 22480
rect 23938 22264 23994 22273
rect 23938 22199 23994 22208
rect 23848 22092 23900 22098
rect 23768 22052 23848 22080
rect 23848 22034 23900 22040
rect 23756 21548 23808 21554
rect 23756 21490 23808 21496
rect 23768 20777 23796 21490
rect 23754 20768 23810 20777
rect 23754 20703 23810 20712
rect 23676 20420 23796 20448
rect 23480 20324 23532 20330
rect 23480 20266 23532 20272
rect 23664 20324 23716 20330
rect 23664 20266 23716 20272
rect 23388 19916 23440 19922
rect 23388 19858 23440 19864
rect 23572 19848 23624 19854
rect 23572 19790 23624 19796
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 23110 19479 23166 19488
rect 23296 19508 23348 19514
rect 23124 19334 23152 19479
rect 23296 19450 23348 19456
rect 23492 19446 23520 19654
rect 23584 19553 23612 19790
rect 23570 19544 23626 19553
rect 23570 19479 23626 19488
rect 23480 19440 23532 19446
rect 23480 19382 23532 19388
rect 23388 19372 23440 19378
rect 23124 19306 23244 19334
rect 23388 19314 23440 19320
rect 23572 19372 23624 19378
rect 23572 19314 23624 19320
rect 23112 18896 23164 18902
rect 23112 18838 23164 18844
rect 23124 15162 23152 18838
rect 23216 18766 23244 19306
rect 23400 18970 23428 19314
rect 23388 18964 23440 18970
rect 23388 18906 23440 18912
rect 23204 18760 23256 18766
rect 23204 18702 23256 18708
rect 23112 15156 23164 15162
rect 23112 15098 23164 15104
rect 23112 14408 23164 14414
rect 23032 14368 23112 14396
rect 23112 14350 23164 14356
rect 23020 13932 23072 13938
rect 23020 13874 23072 13880
rect 22836 13796 22888 13802
rect 22836 13738 22888 13744
rect 22744 13456 22796 13462
rect 22742 13424 22744 13433
rect 22796 13424 22798 13433
rect 22742 13359 22798 13368
rect 22848 13326 22876 13738
rect 23032 13530 23060 13874
rect 23112 13864 23164 13870
rect 23112 13806 23164 13812
rect 23020 13524 23072 13530
rect 23020 13466 23072 13472
rect 22928 13388 22980 13394
rect 22928 13330 22980 13336
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22836 13184 22888 13190
rect 22836 13126 22888 13132
rect 22742 12880 22798 12889
rect 22742 12815 22744 12824
rect 22796 12815 22798 12824
rect 22744 12786 22796 12792
rect 22756 11762 22784 12786
rect 22744 11756 22796 11762
rect 22744 11698 22796 11704
rect 22848 9761 22876 13126
rect 22940 12986 22968 13330
rect 23124 13190 23152 13806
rect 23020 13184 23072 13190
rect 23020 13126 23072 13132
rect 23112 13184 23164 13190
rect 23112 13126 23164 13132
rect 22928 12980 22980 12986
rect 22928 12922 22980 12928
rect 22928 12844 22980 12850
rect 22928 12786 22980 12792
rect 22940 12238 22968 12786
rect 22928 12232 22980 12238
rect 22928 12174 22980 12180
rect 23032 11234 23060 13126
rect 23216 12986 23244 18702
rect 23480 17876 23532 17882
rect 23480 17818 23532 17824
rect 23388 17672 23440 17678
rect 23388 17614 23440 17620
rect 23296 17128 23348 17134
rect 23296 17070 23348 17076
rect 23204 12980 23256 12986
rect 23204 12922 23256 12928
rect 23204 11688 23256 11694
rect 23204 11630 23256 11636
rect 23110 11520 23166 11529
rect 23110 11455 23166 11464
rect 22940 11206 23060 11234
rect 22940 10577 22968 11206
rect 23020 11008 23072 11014
rect 23020 10950 23072 10956
rect 23032 10674 23060 10950
rect 23124 10810 23152 11455
rect 23216 11150 23244 11630
rect 23204 11144 23256 11150
rect 23204 11086 23256 11092
rect 23112 10804 23164 10810
rect 23112 10746 23164 10752
rect 23020 10668 23072 10674
rect 23020 10610 23072 10616
rect 22926 10568 22982 10577
rect 23124 10554 23152 10746
rect 22926 10503 22982 10512
rect 23032 10526 23152 10554
rect 22834 9752 22890 9761
rect 22834 9687 22890 9696
rect 22572 9438 22692 9466
rect 22572 9382 22600 9438
rect 22560 9376 22612 9382
rect 22560 9318 22612 9324
rect 22560 9104 22612 9110
rect 22560 9046 22612 9052
rect 22468 7880 22520 7886
rect 22468 7822 22520 7828
rect 22376 7472 22428 7478
rect 22376 7414 22428 7420
rect 21456 6928 21508 6934
rect 21456 6870 21508 6876
rect 22284 6928 22336 6934
rect 22284 6870 22336 6876
rect 21548 6724 21600 6730
rect 21548 6666 21600 6672
rect 21560 5914 21588 6666
rect 22388 6390 22416 7414
rect 22572 7206 22600 9046
rect 22744 8900 22796 8906
rect 22744 8842 22796 8848
rect 22756 8498 22784 8842
rect 22744 8492 22796 8498
rect 22744 8434 22796 8440
rect 22652 8424 22704 8430
rect 22652 8366 22704 8372
rect 22664 7818 22692 8366
rect 22756 7886 22784 8434
rect 22848 8022 22876 9687
rect 22940 8838 22968 10503
rect 23032 8906 23060 10526
rect 23112 9648 23164 9654
rect 23112 9590 23164 9596
rect 23124 8974 23152 9590
rect 23112 8968 23164 8974
rect 23112 8910 23164 8916
rect 23020 8900 23072 8906
rect 23020 8842 23072 8848
rect 22928 8832 22980 8838
rect 22928 8774 22980 8780
rect 22836 8016 22888 8022
rect 22836 7958 22888 7964
rect 22744 7880 22796 7886
rect 22744 7822 22796 7828
rect 22652 7812 22704 7818
rect 22652 7754 22704 7760
rect 22940 7750 22968 8774
rect 23124 8634 23152 8910
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 23020 7948 23072 7954
rect 23124 7936 23152 8570
rect 23072 7908 23152 7936
rect 23020 7890 23072 7896
rect 22928 7744 22980 7750
rect 22928 7686 22980 7692
rect 22560 7200 22612 7206
rect 22560 7142 22612 7148
rect 22376 6384 22428 6390
rect 22376 6326 22428 6332
rect 23020 6248 23072 6254
rect 22374 6216 22430 6225
rect 22284 6180 22336 6186
rect 23020 6190 23072 6196
rect 22374 6151 22430 6160
rect 22284 6122 22336 6128
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 21364 5840 21416 5846
rect 21364 5782 21416 5788
rect 21560 5710 21588 5850
rect 21272 5704 21324 5710
rect 21272 5646 21324 5652
rect 21548 5704 21600 5710
rect 21548 5646 21600 5652
rect 21732 5704 21784 5710
rect 21732 5646 21784 5652
rect 22100 5704 22152 5710
rect 22100 5646 22152 5652
rect 21744 5574 21772 5646
rect 21732 5568 21784 5574
rect 21732 5510 21784 5516
rect 21362 5400 21418 5409
rect 21362 5335 21364 5344
rect 21416 5335 21418 5344
rect 21364 5306 21416 5312
rect 21456 5228 21508 5234
rect 21456 5170 21508 5176
rect 21272 5024 21324 5030
rect 21272 4966 21324 4972
rect 21284 4214 21312 4966
rect 21468 4826 21496 5170
rect 21456 4820 21508 4826
rect 21456 4762 21508 4768
rect 21468 4214 21496 4762
rect 21640 4548 21692 4554
rect 21640 4490 21692 4496
rect 21272 4208 21324 4214
rect 21272 4150 21324 4156
rect 21456 4208 21508 4214
rect 21456 4150 21508 4156
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 21180 4072 21232 4078
rect 21180 4014 21232 4020
rect 21362 4040 21418 4049
rect 21362 3975 21418 3984
rect 21376 3534 21404 3975
rect 21560 3738 21588 4082
rect 21548 3732 21600 3738
rect 21548 3674 21600 3680
rect 21652 3618 21680 4490
rect 21744 4146 21772 5510
rect 22112 5234 22140 5646
rect 22204 5642 22232 6054
rect 22192 5636 22244 5642
rect 22192 5578 22244 5584
rect 22296 5370 22324 6122
rect 22388 6118 22416 6151
rect 22376 6112 22428 6118
rect 22376 6054 22428 6060
rect 22468 5636 22520 5642
rect 22468 5578 22520 5584
rect 22376 5568 22428 5574
rect 22376 5510 22428 5516
rect 22284 5364 22336 5370
rect 22284 5306 22336 5312
rect 22388 5302 22416 5510
rect 22480 5370 22508 5578
rect 22468 5364 22520 5370
rect 22468 5306 22520 5312
rect 22376 5296 22428 5302
rect 22376 5238 22428 5244
rect 23032 5234 23060 6190
rect 23216 5778 23244 11086
rect 23308 10656 23336 17070
rect 23400 16561 23428 17614
rect 23492 17542 23520 17818
rect 23480 17536 23532 17542
rect 23480 17478 23532 17484
rect 23386 16552 23442 16561
rect 23386 16487 23442 16496
rect 23400 16454 23428 16487
rect 23388 16448 23440 16454
rect 23388 16390 23440 16396
rect 23492 14362 23520 17478
rect 23584 14482 23612 19314
rect 23676 17610 23704 20266
rect 23768 19718 23796 20420
rect 23756 19712 23808 19718
rect 23756 19654 23808 19660
rect 23756 19304 23808 19310
rect 23756 19246 23808 19252
rect 23768 18902 23796 19246
rect 23756 18896 23808 18902
rect 23756 18838 23808 18844
rect 23860 18578 23888 22034
rect 23952 20874 23980 22199
rect 24032 22024 24084 22030
rect 24032 21966 24084 21972
rect 23940 20868 23992 20874
rect 23940 20810 23992 20816
rect 24044 20777 24072 21966
rect 24124 21548 24176 21554
rect 24124 21490 24176 21496
rect 24136 21418 24164 21490
rect 24124 21412 24176 21418
rect 24124 21354 24176 21360
rect 24030 20768 24086 20777
rect 24030 20703 24086 20712
rect 23768 18550 23888 18578
rect 23768 17882 23796 18550
rect 23940 18284 23992 18290
rect 23940 18226 23992 18232
rect 23848 18080 23900 18086
rect 23848 18022 23900 18028
rect 23756 17876 23808 17882
rect 23756 17818 23808 17824
rect 23756 17672 23808 17678
rect 23756 17614 23808 17620
rect 23664 17604 23716 17610
rect 23664 17546 23716 17552
rect 23676 15502 23704 17546
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23768 15348 23796 17614
rect 23676 15320 23796 15348
rect 23572 14476 23624 14482
rect 23572 14418 23624 14424
rect 23492 14334 23612 14362
rect 23388 13252 23440 13258
rect 23388 13194 23440 13200
rect 23400 12832 23428 13194
rect 23480 12844 23532 12850
rect 23400 12804 23480 12832
rect 23480 12786 23532 12792
rect 23388 12708 23440 12714
rect 23388 12650 23440 12656
rect 23400 12374 23428 12650
rect 23388 12368 23440 12374
rect 23388 12310 23440 12316
rect 23388 11756 23440 11762
rect 23388 11698 23440 11704
rect 23400 10996 23428 11698
rect 23400 10968 23520 10996
rect 23388 10668 23440 10674
rect 23308 10628 23388 10656
rect 23388 10610 23440 10616
rect 23294 8664 23350 8673
rect 23294 8599 23296 8608
rect 23348 8599 23350 8608
rect 23296 8570 23348 8576
rect 23308 7410 23336 8570
rect 23400 8090 23428 10610
rect 23492 9178 23520 10968
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23492 8294 23520 9114
rect 23480 8288 23532 8294
rect 23480 8230 23532 8236
rect 23388 8084 23440 8090
rect 23388 8026 23440 8032
rect 23296 7404 23348 7410
rect 23296 7346 23348 7352
rect 23584 6118 23612 14334
rect 23676 12628 23704 15320
rect 23756 14272 23808 14278
rect 23756 14214 23808 14220
rect 23768 14074 23796 14214
rect 23756 14068 23808 14074
rect 23756 14010 23808 14016
rect 23756 13524 23808 13530
rect 23756 13466 23808 13472
rect 23768 12730 23796 13466
rect 23860 12850 23888 18022
rect 23952 14521 23980 18226
rect 24124 18216 24176 18222
rect 24124 18158 24176 18164
rect 24136 15434 24164 18158
rect 24228 17678 24256 23598
rect 24308 22636 24360 22642
rect 24308 22578 24360 22584
rect 24320 20262 24348 22578
rect 24412 22522 24440 24210
rect 24492 23316 24544 23322
rect 24492 23258 24544 23264
rect 24504 22642 24532 23258
rect 24492 22636 24544 22642
rect 24492 22578 24544 22584
rect 24412 22494 24532 22522
rect 24400 21888 24452 21894
rect 24400 21830 24452 21836
rect 24412 21690 24440 21830
rect 24400 21684 24452 21690
rect 24400 21626 24452 21632
rect 24400 21548 24452 21554
rect 24400 21490 24452 21496
rect 24308 20256 24360 20262
rect 24308 20198 24360 20204
rect 24308 19712 24360 19718
rect 24308 19654 24360 19660
rect 24320 19417 24348 19654
rect 24306 19408 24362 19417
rect 24306 19343 24362 19352
rect 24320 17746 24348 19343
rect 24412 19334 24440 21490
rect 24504 19854 24532 22494
rect 24596 21554 24624 25230
rect 24766 24848 24822 24857
rect 24964 24818 24992 31214
rect 25056 30054 25084 32370
rect 25332 32230 25360 32370
rect 25424 32337 25452 32370
rect 25410 32328 25466 32337
rect 25410 32263 25466 32272
rect 25320 32224 25372 32230
rect 25320 32166 25372 32172
rect 25332 32026 25360 32166
rect 25320 32020 25372 32026
rect 25320 31962 25372 31968
rect 25228 31816 25280 31822
rect 25228 31758 25280 31764
rect 25044 30048 25096 30054
rect 25044 29990 25096 29996
rect 25056 29714 25084 29990
rect 25044 29708 25096 29714
rect 25044 29650 25096 29656
rect 25136 29640 25188 29646
rect 25042 29608 25098 29617
rect 25136 29582 25188 29588
rect 25042 29543 25098 29552
rect 25056 29084 25084 29543
rect 25148 29238 25176 29582
rect 25136 29232 25188 29238
rect 25136 29174 25188 29180
rect 25136 29096 25188 29102
rect 25056 29056 25136 29084
rect 25136 29038 25188 29044
rect 25044 28552 25096 28558
rect 25044 28494 25096 28500
rect 25136 28552 25188 28558
rect 25136 28494 25188 28500
rect 25056 26586 25084 28494
rect 25148 27878 25176 28494
rect 25136 27872 25188 27878
rect 25136 27814 25188 27820
rect 25240 27062 25268 31758
rect 25332 29646 25360 31962
rect 25424 31414 25452 32263
rect 25516 31804 25544 32864
rect 26148 32904 26200 32910
rect 25780 32846 25832 32852
rect 26146 32872 26148 32881
rect 26200 32872 26202 32881
rect 26146 32807 26202 32816
rect 25596 32768 25648 32774
rect 25596 32710 25648 32716
rect 26424 32768 26476 32774
rect 26424 32710 26476 32716
rect 25608 32473 25636 32710
rect 25688 32564 25740 32570
rect 25688 32506 25740 32512
rect 25780 32564 25832 32570
rect 25780 32506 25832 32512
rect 25594 32464 25650 32473
rect 25594 32399 25596 32408
rect 25648 32399 25650 32408
rect 25596 32370 25648 32376
rect 25700 31822 25728 32506
rect 25792 31958 25820 32506
rect 26436 32502 26464 32710
rect 26424 32496 26476 32502
rect 26424 32438 26476 32444
rect 26056 32428 26108 32434
rect 26056 32370 26108 32376
rect 26332 32428 26384 32434
rect 26332 32370 26384 32376
rect 25780 31952 25832 31958
rect 25780 31894 25832 31900
rect 25596 31816 25648 31822
rect 25516 31776 25596 31804
rect 25596 31758 25648 31764
rect 25688 31816 25740 31822
rect 25688 31758 25740 31764
rect 25412 31408 25464 31414
rect 25412 31350 25464 31356
rect 25410 31104 25466 31113
rect 25410 31039 25466 31048
rect 25424 30054 25452 31039
rect 25608 30190 25636 31758
rect 25792 31482 25820 31894
rect 26068 31482 26096 32370
rect 26148 32224 26200 32230
rect 26148 32166 26200 32172
rect 26160 31822 26188 32166
rect 26148 31816 26200 31822
rect 26148 31758 26200 31764
rect 26148 31680 26200 31686
rect 26148 31622 26200 31628
rect 25780 31476 25832 31482
rect 26056 31476 26108 31482
rect 25780 31418 25832 31424
rect 25884 31436 26056 31464
rect 25884 31362 25912 31436
rect 26056 31418 26108 31424
rect 25700 31346 25912 31362
rect 25688 31340 25912 31346
rect 25740 31334 25912 31340
rect 25964 31340 26016 31346
rect 25688 31282 25740 31288
rect 25964 31282 26016 31288
rect 25976 30841 26004 31282
rect 25962 30832 26018 30841
rect 25962 30767 26018 30776
rect 25872 30660 25924 30666
rect 25872 30602 25924 30608
rect 25884 30326 25912 30602
rect 25872 30320 25924 30326
rect 25872 30262 25924 30268
rect 25596 30184 25648 30190
rect 25596 30126 25648 30132
rect 25780 30116 25832 30122
rect 25780 30058 25832 30064
rect 25412 30048 25464 30054
rect 25412 29990 25464 29996
rect 25320 29640 25372 29646
rect 25318 29608 25320 29617
rect 25372 29608 25374 29617
rect 25318 29543 25374 29552
rect 25424 29170 25452 29990
rect 25792 29889 25820 30058
rect 25778 29880 25834 29889
rect 25778 29815 25834 29824
rect 25688 29572 25740 29578
rect 25740 29532 25820 29560
rect 25688 29514 25740 29520
rect 25516 29260 25728 29288
rect 25516 29170 25544 29260
rect 25412 29164 25464 29170
rect 25412 29106 25464 29112
rect 25504 29164 25556 29170
rect 25504 29106 25556 29112
rect 25596 29164 25648 29170
rect 25596 29106 25648 29112
rect 25320 29028 25372 29034
rect 25320 28970 25372 28976
rect 25228 27056 25280 27062
rect 25228 26998 25280 27004
rect 25332 26994 25360 28970
rect 25424 28218 25452 29106
rect 25608 28626 25636 29106
rect 25596 28620 25648 28626
rect 25596 28562 25648 28568
rect 25504 28552 25556 28558
rect 25608 28529 25636 28562
rect 25504 28494 25556 28500
rect 25594 28520 25650 28529
rect 25516 28218 25544 28494
rect 25594 28455 25650 28464
rect 25412 28212 25464 28218
rect 25412 28154 25464 28160
rect 25504 28212 25556 28218
rect 25504 28154 25556 28160
rect 25700 27520 25728 29260
rect 25792 29238 25820 29532
rect 25780 29232 25832 29238
rect 25780 29174 25832 29180
rect 25792 28558 25820 29174
rect 25884 28626 25912 30262
rect 26056 30184 26108 30190
rect 26056 30126 26108 30132
rect 25964 30116 26016 30122
rect 25964 30058 26016 30064
rect 25872 28620 25924 28626
rect 25872 28562 25924 28568
rect 25780 28552 25832 28558
rect 25780 28494 25832 28500
rect 25780 28008 25832 28014
rect 25780 27950 25832 27956
rect 25516 27492 25728 27520
rect 25320 26988 25372 26994
rect 25320 26930 25372 26936
rect 25516 26874 25544 27492
rect 25792 27402 25820 27950
rect 25872 27940 25924 27946
rect 25872 27882 25924 27888
rect 25596 27396 25648 27402
rect 25780 27396 25832 27402
rect 25596 27338 25648 27344
rect 25700 27356 25780 27384
rect 25332 26846 25544 26874
rect 25044 26580 25096 26586
rect 25044 26522 25096 26528
rect 25136 26512 25188 26518
rect 25136 26454 25188 26460
rect 25228 26512 25280 26518
rect 25228 26454 25280 26460
rect 25044 26308 25096 26314
rect 25044 26250 25096 26256
rect 24766 24783 24768 24792
rect 24820 24783 24822 24792
rect 24952 24812 25004 24818
rect 24768 24754 24820 24760
rect 24952 24754 25004 24760
rect 24676 24676 24728 24682
rect 24676 24618 24728 24624
rect 24688 24206 24716 24618
rect 24780 24274 24808 24754
rect 24768 24268 24820 24274
rect 24768 24210 24820 24216
rect 24676 24200 24728 24206
rect 24676 24142 24728 24148
rect 24952 22636 25004 22642
rect 24952 22578 25004 22584
rect 24676 22432 24728 22438
rect 24676 22374 24728 22380
rect 24584 21548 24636 21554
rect 24584 21490 24636 21496
rect 24492 19848 24544 19854
rect 24492 19790 24544 19796
rect 24504 19446 24532 19790
rect 24584 19712 24636 19718
rect 24584 19654 24636 19660
rect 24492 19440 24544 19446
rect 24492 19382 24544 19388
rect 24412 19306 24532 19334
rect 24398 19000 24454 19009
rect 24398 18935 24454 18944
rect 24412 18766 24440 18935
rect 24400 18760 24452 18766
rect 24400 18702 24452 18708
rect 24308 17740 24360 17746
rect 24308 17682 24360 17688
rect 24216 17672 24268 17678
rect 24216 17614 24268 17620
rect 24400 17604 24452 17610
rect 24400 17546 24452 17552
rect 24216 17536 24268 17542
rect 24216 17478 24268 17484
rect 24228 17202 24256 17478
rect 24412 17338 24440 17546
rect 24400 17332 24452 17338
rect 24400 17274 24452 17280
rect 24216 17196 24268 17202
rect 24216 17138 24268 17144
rect 24504 16590 24532 19306
rect 24596 18834 24624 19654
rect 24584 18828 24636 18834
rect 24584 18770 24636 18776
rect 24596 18630 24624 18770
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 24492 16584 24544 16590
rect 24492 16526 24544 16532
rect 24492 16448 24544 16454
rect 24492 16390 24544 16396
rect 24504 16114 24532 16390
rect 24492 16108 24544 16114
rect 24492 16050 24544 16056
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24032 15428 24084 15434
rect 24032 15370 24084 15376
rect 24124 15428 24176 15434
rect 24124 15370 24176 15376
rect 24044 14550 24072 15370
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 24032 14544 24084 14550
rect 23938 14512 23994 14521
rect 24032 14486 24084 14492
rect 23938 14447 23994 14456
rect 23952 14278 23980 14447
rect 23940 14272 23992 14278
rect 23940 14214 23992 14220
rect 23938 14104 23994 14113
rect 24228 14074 24256 14962
rect 24412 14958 24440 15438
rect 24504 14958 24532 16050
rect 24596 15586 24624 18566
rect 24688 18290 24716 22374
rect 24766 22128 24822 22137
rect 24766 22063 24822 22072
rect 24676 18284 24728 18290
rect 24676 18226 24728 18232
rect 24780 18222 24808 22063
rect 24860 21548 24912 21554
rect 24860 21490 24912 21496
rect 24872 19825 24900 21490
rect 24964 20398 24992 22578
rect 25056 22098 25084 26250
rect 25148 24342 25176 26454
rect 25240 25498 25268 26454
rect 25228 25492 25280 25498
rect 25228 25434 25280 25440
rect 25136 24336 25188 24342
rect 25136 24278 25188 24284
rect 25136 24200 25188 24206
rect 25134 24168 25136 24177
rect 25188 24168 25190 24177
rect 25134 24103 25190 24112
rect 25044 22092 25096 22098
rect 25044 22034 25096 22040
rect 25044 21956 25096 21962
rect 25044 21898 25096 21904
rect 25056 21690 25084 21898
rect 25044 21684 25096 21690
rect 25044 21626 25096 21632
rect 25056 21078 25084 21626
rect 25044 21072 25096 21078
rect 25044 21014 25096 21020
rect 25044 20460 25096 20466
rect 25044 20402 25096 20408
rect 24952 20392 25004 20398
rect 24952 20334 25004 20340
rect 24858 19816 24914 19825
rect 24858 19751 24914 19760
rect 24768 18216 24820 18222
rect 24768 18158 24820 18164
rect 24674 17368 24730 17377
rect 24674 17303 24730 17312
rect 24688 17202 24716 17303
rect 24676 17196 24728 17202
rect 24676 17138 24728 17144
rect 24872 16998 24900 19751
rect 24964 18970 24992 20334
rect 25056 19922 25084 20402
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 25148 20058 25176 20334
rect 25136 20052 25188 20058
rect 25136 19994 25188 20000
rect 25044 19916 25096 19922
rect 25044 19858 25096 19864
rect 24952 18964 25004 18970
rect 24952 18906 25004 18912
rect 24952 18760 25004 18766
rect 24952 18702 25004 18708
rect 24860 16992 24912 16998
rect 24860 16934 24912 16940
rect 24768 16516 24820 16522
rect 24768 16458 24820 16464
rect 24780 16250 24808 16458
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 24676 16108 24728 16114
rect 24676 16050 24728 16056
rect 24688 15706 24716 16050
rect 24676 15700 24728 15706
rect 24676 15642 24728 15648
rect 24596 15558 24808 15586
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24688 15162 24716 15438
rect 24676 15156 24728 15162
rect 24676 15098 24728 15104
rect 24674 15056 24730 15065
rect 24674 14991 24676 15000
rect 24728 14991 24730 15000
rect 24676 14962 24728 14968
rect 24400 14952 24452 14958
rect 24400 14894 24452 14900
rect 24492 14952 24544 14958
rect 24492 14894 24544 14900
rect 24676 14884 24728 14890
rect 24676 14826 24728 14832
rect 24400 14816 24452 14822
rect 24400 14758 24452 14764
rect 24308 14476 24360 14482
rect 24308 14418 24360 14424
rect 24320 14074 24348 14418
rect 23938 14039 23940 14048
rect 23992 14039 23994 14048
rect 24216 14068 24268 14074
rect 23940 14010 23992 14016
rect 24216 14010 24268 14016
rect 24308 14068 24360 14074
rect 24308 14010 24360 14016
rect 24124 14000 24176 14006
rect 24044 13960 24124 13988
rect 23940 13728 23992 13734
rect 23940 13670 23992 13676
rect 23952 12850 23980 13670
rect 23848 12844 23900 12850
rect 23848 12786 23900 12792
rect 23940 12844 23992 12850
rect 23940 12786 23992 12792
rect 23768 12702 23980 12730
rect 23848 12640 23900 12646
rect 23676 12600 23796 12628
rect 23662 12472 23718 12481
rect 23662 12407 23718 12416
rect 23572 6112 23624 6118
rect 23572 6054 23624 6060
rect 23204 5772 23256 5778
rect 23204 5714 23256 5720
rect 23676 5658 23704 12407
rect 23768 8566 23796 12600
rect 23848 12582 23900 12588
rect 23860 12481 23888 12582
rect 23846 12472 23902 12481
rect 23846 12407 23902 12416
rect 23848 12368 23900 12374
rect 23848 12310 23900 12316
rect 23860 10062 23888 12310
rect 23848 10056 23900 10062
rect 23848 9998 23900 10004
rect 23952 9586 23980 12702
rect 24044 10810 24072 13960
rect 24124 13942 24176 13948
rect 24124 13864 24176 13870
rect 24124 13806 24176 13812
rect 24032 10804 24084 10810
rect 24032 10746 24084 10752
rect 24136 10538 24164 13806
rect 24216 13184 24268 13190
rect 24216 13126 24268 13132
rect 24228 11762 24256 13126
rect 24216 11756 24268 11762
rect 24216 11698 24268 11704
rect 24228 10724 24256 11698
rect 24412 11354 24440 14758
rect 24688 14414 24716 14826
rect 24584 14408 24636 14414
rect 24584 14350 24636 14356
rect 24676 14408 24728 14414
rect 24676 14350 24728 14356
rect 24490 14104 24546 14113
rect 24490 14039 24492 14048
rect 24544 14039 24546 14048
rect 24492 14010 24544 14016
rect 24492 13864 24544 13870
rect 24492 13806 24544 13812
rect 24504 13734 24532 13806
rect 24492 13728 24544 13734
rect 24492 13670 24544 13676
rect 24596 12850 24624 14350
rect 24676 14000 24728 14006
rect 24674 13968 24676 13977
rect 24728 13968 24730 13977
rect 24674 13903 24730 13912
rect 24584 12844 24636 12850
rect 24584 12786 24636 12792
rect 24492 12640 24544 12646
rect 24492 12582 24544 12588
rect 24504 11937 24532 12582
rect 24490 11928 24546 11937
rect 24780 11914 24808 15558
rect 24964 14618 24992 18702
rect 25056 17218 25084 19858
rect 25136 19780 25188 19786
rect 25136 19722 25188 19728
rect 25148 19378 25176 19722
rect 25136 19372 25188 19378
rect 25136 19314 25188 19320
rect 25240 18902 25268 25434
rect 25332 23769 25360 26846
rect 25504 26512 25556 26518
rect 25504 26454 25556 26460
rect 25516 26382 25544 26454
rect 25504 26376 25556 26382
rect 25504 26318 25556 26324
rect 25412 25356 25464 25362
rect 25412 25298 25464 25304
rect 25424 24857 25452 25298
rect 25410 24848 25466 24857
rect 25410 24783 25466 24792
rect 25412 24744 25464 24750
rect 25412 24686 25464 24692
rect 25318 23760 25374 23769
rect 25318 23695 25374 23704
rect 25424 22778 25452 24686
rect 25412 22772 25464 22778
rect 25412 22714 25464 22720
rect 25320 22704 25372 22710
rect 25320 22646 25372 22652
rect 25332 22234 25360 22646
rect 25320 22228 25372 22234
rect 25320 22170 25372 22176
rect 25320 20528 25372 20534
rect 25320 20470 25372 20476
rect 25332 20369 25360 20470
rect 25318 20360 25374 20369
rect 25318 20295 25374 20304
rect 25412 20324 25464 20330
rect 25412 20266 25464 20272
rect 25320 20256 25372 20262
rect 25320 20198 25372 20204
rect 25332 20058 25360 20198
rect 25424 20058 25452 20266
rect 25516 20262 25544 26318
rect 25608 26042 25636 27338
rect 25700 26314 25728 27356
rect 25780 27338 25832 27344
rect 25780 26988 25832 26994
rect 25780 26930 25832 26936
rect 25688 26308 25740 26314
rect 25688 26250 25740 26256
rect 25792 26042 25820 26930
rect 25884 26586 25912 27882
rect 25976 27130 26004 30058
rect 26068 28082 26096 30126
rect 26160 29578 26188 31622
rect 26240 30728 26292 30734
rect 26240 30670 26292 30676
rect 26252 30190 26280 30670
rect 26240 30184 26292 30190
rect 26240 30126 26292 30132
rect 26240 30048 26292 30054
rect 26240 29990 26292 29996
rect 26252 29646 26280 29990
rect 26240 29640 26292 29646
rect 26240 29582 26292 29588
rect 26148 29572 26200 29578
rect 26148 29514 26200 29520
rect 26252 29170 26280 29582
rect 26240 29164 26292 29170
rect 26240 29106 26292 29112
rect 26252 28762 26280 29106
rect 26240 28756 26292 28762
rect 26240 28698 26292 28704
rect 26148 28552 26200 28558
rect 26146 28520 26148 28529
rect 26200 28520 26202 28529
rect 26146 28455 26202 28464
rect 26056 28076 26108 28082
rect 26056 28018 26108 28024
rect 25964 27124 26016 27130
rect 25964 27066 26016 27072
rect 25872 26580 25924 26586
rect 25872 26522 25924 26528
rect 26068 26314 26096 28018
rect 26056 26308 26108 26314
rect 26056 26250 26108 26256
rect 25596 26036 25648 26042
rect 25596 25978 25648 25984
rect 25780 26036 25832 26042
rect 25780 25978 25832 25984
rect 26056 25900 26108 25906
rect 26056 25842 26108 25848
rect 26068 25294 26096 25842
rect 26148 25764 26200 25770
rect 26148 25706 26200 25712
rect 25688 25288 25740 25294
rect 25688 25230 25740 25236
rect 25872 25288 25924 25294
rect 25872 25230 25924 25236
rect 26056 25288 26108 25294
rect 26056 25230 26108 25236
rect 26160 25276 26188 25706
rect 26240 25288 26292 25294
rect 26160 25248 26240 25276
rect 25700 24954 25728 25230
rect 25688 24948 25740 24954
rect 25688 24890 25740 24896
rect 25780 24880 25832 24886
rect 25780 24822 25832 24828
rect 25792 24698 25820 24822
rect 25608 24670 25820 24698
rect 25608 24410 25636 24670
rect 25688 24608 25740 24614
rect 25688 24550 25740 24556
rect 25780 24608 25832 24614
rect 25780 24550 25832 24556
rect 25596 24404 25648 24410
rect 25596 24346 25648 24352
rect 25596 23792 25648 23798
rect 25596 23734 25648 23740
rect 25608 21622 25636 23734
rect 25700 22778 25728 24550
rect 25792 24138 25820 24550
rect 25884 24410 25912 25230
rect 25964 24948 26016 24954
rect 25964 24890 26016 24896
rect 25872 24404 25924 24410
rect 25872 24346 25924 24352
rect 25976 24290 26004 24890
rect 25884 24262 26004 24290
rect 25884 24206 25912 24262
rect 25872 24200 25924 24206
rect 25870 24168 25872 24177
rect 25924 24168 25926 24177
rect 25780 24132 25832 24138
rect 25870 24103 25926 24112
rect 25780 24074 25832 24080
rect 25872 24064 25924 24070
rect 25872 24006 25924 24012
rect 25884 23254 25912 24006
rect 25872 23248 25924 23254
rect 25872 23190 25924 23196
rect 25688 22772 25740 22778
rect 25688 22714 25740 22720
rect 25872 22568 25924 22574
rect 25872 22510 25924 22516
rect 25964 22568 26016 22574
rect 25964 22510 26016 22516
rect 25688 22432 25740 22438
rect 25688 22374 25740 22380
rect 25596 21616 25648 21622
rect 25596 21558 25648 21564
rect 25608 20641 25636 21558
rect 25700 21554 25728 22374
rect 25780 22024 25832 22030
rect 25884 21978 25912 22510
rect 25832 21972 25912 21978
rect 25780 21966 25912 21972
rect 25792 21950 25912 21966
rect 25780 21684 25832 21690
rect 25780 21626 25832 21632
rect 25688 21548 25740 21554
rect 25688 21490 25740 21496
rect 25594 20632 25650 20641
rect 25594 20567 25650 20576
rect 25688 20460 25740 20466
rect 25688 20402 25740 20408
rect 25504 20256 25556 20262
rect 25504 20198 25556 20204
rect 25320 20052 25372 20058
rect 25320 19994 25372 20000
rect 25412 20052 25464 20058
rect 25412 19994 25464 20000
rect 25228 18896 25280 18902
rect 25228 18838 25280 18844
rect 25136 18624 25188 18630
rect 25240 18578 25268 18838
rect 25188 18572 25268 18578
rect 25136 18566 25268 18572
rect 25148 18550 25268 18566
rect 25136 17264 25188 17270
rect 25056 17212 25136 17218
rect 25056 17206 25188 17212
rect 25056 17190 25176 17206
rect 25044 17128 25096 17134
rect 25044 17070 25096 17076
rect 24952 14612 25004 14618
rect 24952 14554 25004 14560
rect 25056 14521 25084 17070
rect 25148 15094 25176 17190
rect 25332 17082 25360 19994
rect 25504 19780 25556 19786
rect 25504 19722 25556 19728
rect 25516 19514 25544 19722
rect 25504 19508 25556 19514
rect 25504 19450 25556 19456
rect 25412 19372 25464 19378
rect 25412 19314 25464 19320
rect 25424 18698 25452 19314
rect 25412 18692 25464 18698
rect 25412 18634 25464 18640
rect 25700 18630 25728 20402
rect 25792 20380 25820 21626
rect 25884 20534 25912 21950
rect 25976 21894 26004 22510
rect 25964 21888 26016 21894
rect 25964 21830 26016 21836
rect 25964 20868 26016 20874
rect 25964 20810 26016 20816
rect 25872 20528 25924 20534
rect 25872 20470 25924 20476
rect 25792 20352 25912 20380
rect 25780 19984 25832 19990
rect 25780 19926 25832 19932
rect 25792 18766 25820 19926
rect 25780 18760 25832 18766
rect 25780 18702 25832 18708
rect 25688 18624 25740 18630
rect 25688 18566 25740 18572
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 25228 17060 25280 17066
rect 25332 17054 25452 17082
rect 25228 17002 25280 17008
rect 25240 16946 25268 17002
rect 25240 16918 25360 16946
rect 25228 16108 25280 16114
rect 25228 16050 25280 16056
rect 25136 15088 25188 15094
rect 25136 15030 25188 15036
rect 25042 14512 25098 14521
rect 24952 14476 25004 14482
rect 25042 14447 25098 14456
rect 24952 14418 25004 14424
rect 24860 13252 24912 13258
rect 24860 13194 24912 13200
rect 24872 12850 24900 13194
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24860 12640 24912 12646
rect 24860 12582 24912 12588
rect 24872 12050 24900 12582
rect 24964 12186 24992 14418
rect 25044 14408 25096 14414
rect 25044 14350 25096 14356
rect 25056 13938 25084 14350
rect 25044 13932 25096 13938
rect 25044 13874 25096 13880
rect 25148 12186 25176 15030
rect 25240 12782 25268 16050
rect 25332 14482 25360 16918
rect 25320 14476 25372 14482
rect 25320 14418 25372 14424
rect 25318 14376 25374 14385
rect 25318 14311 25374 14320
rect 25228 12776 25280 12782
rect 25228 12718 25280 12724
rect 25332 12646 25360 14311
rect 25320 12640 25372 12646
rect 25320 12582 25372 12588
rect 25424 12434 25452 17054
rect 25504 16584 25556 16590
rect 25504 16526 25556 16532
rect 25516 14618 25544 16526
rect 25608 16522 25636 17138
rect 25700 16658 25728 18566
rect 25792 18358 25820 18702
rect 25780 18352 25832 18358
rect 25780 18294 25832 18300
rect 25688 16652 25740 16658
rect 25688 16594 25740 16600
rect 25780 16652 25832 16658
rect 25780 16594 25832 16600
rect 25596 16516 25648 16522
rect 25596 16458 25648 16464
rect 25608 15502 25636 16458
rect 25700 16182 25728 16594
rect 25688 16176 25740 16182
rect 25688 16118 25740 16124
rect 25596 15496 25648 15502
rect 25596 15438 25648 15444
rect 25504 14612 25556 14618
rect 25504 14554 25556 14560
rect 25596 13252 25648 13258
rect 25596 13194 25648 13200
rect 25608 12850 25636 13194
rect 25596 12844 25648 12850
rect 25596 12786 25648 12792
rect 25424 12406 25544 12434
rect 24964 12158 25084 12186
rect 25148 12158 25268 12186
rect 24872 12022 24992 12050
rect 24490 11863 24546 11872
rect 24688 11886 24808 11914
rect 24504 11762 24532 11863
rect 24492 11756 24544 11762
rect 24492 11698 24544 11704
rect 24400 11348 24452 11354
rect 24400 11290 24452 11296
rect 24308 10736 24360 10742
rect 24228 10696 24308 10724
rect 24308 10678 24360 10684
rect 24492 10736 24544 10742
rect 24492 10678 24544 10684
rect 24124 10532 24176 10538
rect 24124 10474 24176 10480
rect 24136 9722 24164 10474
rect 24320 10198 24348 10678
rect 24308 10192 24360 10198
rect 24308 10134 24360 10140
rect 24308 10056 24360 10062
rect 24504 10044 24532 10678
rect 24360 10016 24532 10044
rect 24308 9998 24360 10004
rect 24124 9716 24176 9722
rect 24124 9658 24176 9664
rect 23940 9580 23992 9586
rect 23940 9522 23992 9528
rect 23848 8628 23900 8634
rect 23848 8570 23900 8576
rect 23756 8560 23808 8566
rect 23756 8502 23808 8508
rect 23768 6254 23796 8502
rect 23860 8401 23888 8570
rect 23846 8392 23902 8401
rect 23952 8362 23980 9522
rect 24136 9110 24164 9658
rect 24124 9104 24176 9110
rect 24124 9046 24176 9052
rect 24032 8832 24084 8838
rect 24032 8774 24084 8780
rect 24044 8498 24072 8774
rect 24136 8566 24164 9046
rect 24216 8968 24268 8974
rect 24214 8936 24216 8945
rect 24268 8936 24270 8945
rect 24214 8871 24270 8880
rect 24214 8664 24270 8673
rect 24214 8599 24270 8608
rect 24228 8566 24256 8599
rect 24124 8560 24176 8566
rect 24124 8502 24176 8508
rect 24216 8560 24268 8566
rect 24216 8502 24268 8508
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 23846 8327 23902 8336
rect 23940 8356 23992 8362
rect 23940 8298 23992 8304
rect 23848 8288 23900 8294
rect 23848 8230 23900 8236
rect 23860 7721 23888 8230
rect 24124 7880 24176 7886
rect 24122 7848 24124 7857
rect 24176 7848 24178 7857
rect 24122 7783 24178 7792
rect 23846 7712 23902 7721
rect 23846 7647 23902 7656
rect 24320 7410 24348 9998
rect 24400 9920 24452 9926
rect 24400 9862 24452 9868
rect 24412 8906 24440 9862
rect 24688 9194 24716 11886
rect 24860 11824 24912 11830
rect 24860 11766 24912 11772
rect 24768 11552 24820 11558
rect 24768 11494 24820 11500
rect 24780 11354 24808 11494
rect 24768 11348 24820 11354
rect 24768 11290 24820 11296
rect 24768 11144 24820 11150
rect 24872 11121 24900 11766
rect 24964 11762 24992 12022
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 24964 11558 24992 11698
rect 24952 11552 25004 11558
rect 24952 11494 25004 11500
rect 24768 11086 24820 11092
rect 24858 11112 24914 11121
rect 24780 10674 24808 11086
rect 24858 11047 24914 11056
rect 25056 10713 25084 12158
rect 25136 12096 25188 12102
rect 25136 12038 25188 12044
rect 25148 11762 25176 12038
rect 25136 11756 25188 11762
rect 25136 11698 25188 11704
rect 25240 11626 25268 12158
rect 25320 11756 25372 11762
rect 25320 11698 25372 11704
rect 25228 11620 25280 11626
rect 25228 11562 25280 11568
rect 25332 11529 25360 11698
rect 25412 11688 25464 11694
rect 25412 11630 25464 11636
rect 25318 11520 25374 11529
rect 25318 11455 25374 11464
rect 25424 11286 25452 11630
rect 25412 11280 25464 11286
rect 25412 11222 25464 11228
rect 25136 11144 25188 11150
rect 25136 11086 25188 11092
rect 25410 11112 25466 11121
rect 25042 10704 25098 10713
rect 24768 10668 24820 10674
rect 25042 10639 25098 10648
rect 24768 10610 24820 10616
rect 24860 10600 24912 10606
rect 24860 10542 24912 10548
rect 24872 10062 24900 10542
rect 25044 10464 25096 10470
rect 25044 10406 25096 10412
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 24766 9344 24822 9353
rect 24766 9279 24822 9288
rect 24780 9194 24808 9279
rect 24584 9172 24636 9178
rect 24688 9166 24808 9194
rect 24584 9114 24636 9120
rect 24400 8900 24452 8906
rect 24400 8842 24452 8848
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 24412 7274 24440 8842
rect 24596 8498 24624 9114
rect 24780 8974 24808 9166
rect 24768 8968 24820 8974
rect 24768 8910 24820 8916
rect 24768 8832 24820 8838
rect 24768 8774 24820 8780
rect 24584 8492 24636 8498
rect 24584 8434 24636 8440
rect 24780 8430 24808 8774
rect 24768 8424 24820 8430
rect 24768 8366 24820 8372
rect 24674 8120 24730 8129
rect 24674 8055 24676 8064
rect 24728 8055 24730 8064
rect 24676 8026 24728 8032
rect 24492 7744 24544 7750
rect 24492 7686 24544 7692
rect 24768 7744 24820 7750
rect 24768 7686 24820 7692
rect 24504 7410 24532 7686
rect 24780 7546 24808 7686
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 24492 7404 24544 7410
rect 24492 7346 24544 7352
rect 24400 7268 24452 7274
rect 24400 7210 24452 7216
rect 24214 7032 24270 7041
rect 24214 6967 24216 6976
rect 24268 6967 24270 6976
rect 24216 6938 24268 6944
rect 23756 6248 23808 6254
rect 23756 6190 23808 6196
rect 24228 5778 24256 6938
rect 24492 6452 24544 6458
rect 24492 6394 24544 6400
rect 24504 5817 24532 6394
rect 24768 6112 24820 6118
rect 24768 6054 24820 6060
rect 24490 5808 24546 5817
rect 24216 5772 24268 5778
rect 24490 5743 24546 5752
rect 24216 5714 24268 5720
rect 23400 5630 23704 5658
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 23020 5228 23072 5234
rect 23020 5170 23072 5176
rect 22376 5160 22428 5166
rect 22376 5102 22428 5108
rect 21732 4140 21784 4146
rect 21732 4082 21784 4088
rect 21824 4140 21876 4146
rect 21824 4082 21876 4088
rect 21836 4049 21864 4082
rect 21822 4040 21878 4049
rect 21822 3975 21878 3984
rect 22388 3942 22416 5102
rect 22836 5092 22888 5098
rect 22836 5034 22888 5040
rect 22652 4548 22704 4554
rect 22652 4490 22704 4496
rect 22664 4282 22692 4490
rect 22652 4276 22704 4282
rect 22652 4218 22704 4224
rect 22376 3936 22428 3942
rect 22848 3913 22876 5034
rect 23032 4282 23060 5170
rect 23112 4684 23164 4690
rect 23112 4626 23164 4632
rect 23020 4276 23072 4282
rect 23020 4218 23072 4224
rect 23020 4140 23072 4146
rect 23020 4082 23072 4088
rect 22376 3878 22428 3884
rect 22834 3904 22890 3913
rect 22834 3839 22890 3848
rect 21560 3590 21680 3618
rect 22744 3596 22796 3602
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21560 3398 21588 3590
rect 22744 3538 22796 3544
rect 21640 3528 21692 3534
rect 21640 3470 21692 3476
rect 21548 3392 21600 3398
rect 21548 3334 21600 3340
rect 21560 3126 21588 3334
rect 21652 3194 21680 3470
rect 21640 3188 21692 3194
rect 21640 3130 21692 3136
rect 21548 3120 21600 3126
rect 21548 3062 21600 3068
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 20168 2984 20220 2990
rect 20168 2926 20220 2932
rect 20812 2984 20864 2990
rect 20812 2926 20864 2932
rect 21916 2984 21968 2990
rect 21916 2926 21968 2932
rect 22468 2984 22520 2990
rect 22468 2926 22520 2932
rect 19352 2650 19380 2926
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 19248 2644 19300 2650
rect 19248 2586 19300 2592
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 19812 2514 19840 2790
rect 20180 2650 20208 2926
rect 20824 2774 20852 2926
rect 20732 2746 20852 2774
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 19800 2508 19852 2514
rect 19800 2450 19852 2456
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 19352 800 19380 2382
rect 20640 800 20668 2382
rect 20732 2378 20760 2746
rect 20720 2372 20772 2378
rect 20720 2314 20772 2320
rect 21364 2304 21416 2310
rect 21284 2264 21364 2292
rect 21284 800 21312 2264
rect 21364 2246 21416 2252
rect 21928 800 21956 2926
rect 22480 2378 22508 2926
rect 22756 2514 22784 3538
rect 22848 3194 22876 3839
rect 22928 3732 22980 3738
rect 22928 3674 22980 3680
rect 22836 3188 22888 3194
rect 22836 3130 22888 3136
rect 22940 2774 22968 3674
rect 23032 3482 23060 4082
rect 23124 3602 23152 4626
rect 23296 4140 23348 4146
rect 23296 4082 23348 4088
rect 23308 3738 23336 4082
rect 23400 4078 23428 5630
rect 24228 5302 24256 5714
rect 24504 5710 24532 5743
rect 24492 5704 24544 5710
rect 24492 5646 24544 5652
rect 24780 5642 24808 6054
rect 24872 5846 24900 9998
rect 25056 9178 25084 10406
rect 25148 10130 25176 11086
rect 25410 11047 25466 11056
rect 25228 10804 25280 10810
rect 25228 10746 25280 10752
rect 25136 10124 25188 10130
rect 25136 10066 25188 10072
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 25148 9518 25176 9862
rect 25136 9512 25188 9518
rect 25136 9454 25188 9460
rect 25240 9382 25268 10746
rect 25424 10742 25452 11047
rect 25412 10736 25464 10742
rect 25318 10704 25374 10713
rect 25412 10678 25464 10684
rect 25318 10639 25320 10648
rect 25372 10639 25374 10648
rect 25320 10610 25372 10616
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 25332 9722 25360 9998
rect 25412 9988 25464 9994
rect 25412 9930 25464 9936
rect 25320 9716 25372 9722
rect 25320 9658 25372 9664
rect 25424 9382 25452 9930
rect 25516 9625 25544 12406
rect 25608 11898 25636 12786
rect 25596 11892 25648 11898
rect 25596 11834 25648 11840
rect 25688 11892 25740 11898
rect 25688 11834 25740 11840
rect 25594 11792 25650 11801
rect 25594 11727 25650 11736
rect 25608 10146 25636 11727
rect 25700 11626 25728 11834
rect 25688 11620 25740 11626
rect 25688 11562 25740 11568
rect 25608 10118 25728 10146
rect 25792 10130 25820 16594
rect 25884 16250 25912 20352
rect 25976 20330 26004 20810
rect 25964 20324 26016 20330
rect 25964 20266 26016 20272
rect 26068 20058 26096 25230
rect 26160 22030 26188 25248
rect 26240 25230 26292 25236
rect 26238 24848 26294 24857
rect 26238 24783 26294 24792
rect 26148 22024 26200 22030
rect 26148 21966 26200 21972
rect 26160 21894 26188 21966
rect 26252 21894 26280 24783
rect 26344 24682 26372 32370
rect 26436 31958 26464 32438
rect 26700 32360 26752 32366
rect 26700 32302 26752 32308
rect 26608 32020 26660 32026
rect 26608 31962 26660 31968
rect 26424 31952 26476 31958
rect 26424 31894 26476 31900
rect 26620 31346 26648 31962
rect 26516 31340 26568 31346
rect 26516 31282 26568 31288
rect 26608 31340 26660 31346
rect 26608 31282 26660 31288
rect 26528 30938 26556 31282
rect 26712 31142 26740 32302
rect 26804 31657 26832 32914
rect 28092 32502 28120 33254
rect 28080 32496 28132 32502
rect 28080 32438 28132 32444
rect 27896 32428 27948 32434
rect 27896 32370 27948 32376
rect 27908 32026 27936 32370
rect 28080 32224 28132 32230
rect 28080 32166 28132 32172
rect 27896 32020 27948 32026
rect 27896 31962 27948 31968
rect 27988 31952 28040 31958
rect 27988 31894 28040 31900
rect 27344 31884 27396 31890
rect 27344 31826 27396 31832
rect 27252 31816 27304 31822
rect 27250 31784 27252 31793
rect 27304 31784 27306 31793
rect 27250 31719 27306 31728
rect 27356 31686 27384 31826
rect 27068 31680 27120 31686
rect 26790 31648 26846 31657
rect 27068 31622 27120 31628
rect 27344 31680 27396 31686
rect 27344 31622 27396 31628
rect 26790 31583 26846 31592
rect 26700 31136 26752 31142
rect 26700 31078 26752 31084
rect 26712 30938 26740 31078
rect 26516 30932 26568 30938
rect 26516 30874 26568 30880
rect 26700 30932 26752 30938
rect 26700 30874 26752 30880
rect 26516 30796 26568 30802
rect 26516 30738 26568 30744
rect 26424 30252 26476 30258
rect 26424 30194 26476 30200
rect 26436 29782 26464 30194
rect 26424 29776 26476 29782
rect 26424 29718 26476 29724
rect 26528 29646 26556 30738
rect 26516 29640 26568 29646
rect 26516 29582 26568 29588
rect 26422 29336 26478 29345
rect 26422 29271 26478 29280
rect 26436 29170 26464 29271
rect 26424 29164 26476 29170
rect 26424 29106 26476 29112
rect 26700 29028 26752 29034
rect 26700 28970 26752 28976
rect 26712 28762 26740 28970
rect 26700 28756 26752 28762
rect 26700 28698 26752 28704
rect 26516 28552 26568 28558
rect 26514 28520 26516 28529
rect 26568 28520 26570 28529
rect 26514 28455 26570 28464
rect 26516 28416 26568 28422
rect 26514 28384 26516 28393
rect 26568 28384 26570 28393
rect 26514 28319 26570 28328
rect 26516 27464 26568 27470
rect 26516 27406 26568 27412
rect 26424 25152 26476 25158
rect 26424 25094 26476 25100
rect 26332 24676 26384 24682
rect 26332 24618 26384 24624
rect 26436 24614 26464 25094
rect 26528 24818 26556 27406
rect 26804 27112 26832 31583
rect 27080 31346 27108 31622
rect 27250 31376 27306 31385
rect 27068 31340 27120 31346
rect 27068 31282 27120 31288
rect 27160 31340 27212 31346
rect 27250 31311 27252 31320
rect 27160 31282 27212 31288
rect 27304 31311 27306 31320
rect 27252 31282 27304 31288
rect 26974 31240 27030 31249
rect 26974 31175 26976 31184
rect 27028 31175 27030 31184
rect 26976 31146 27028 31152
rect 26884 30728 26936 30734
rect 26884 30670 26936 30676
rect 26896 30190 26924 30670
rect 26884 30184 26936 30190
rect 26884 30126 26936 30132
rect 26896 29646 26924 30126
rect 26976 30048 27028 30054
rect 26976 29990 27028 29996
rect 26884 29640 26936 29646
rect 26884 29582 26936 29588
rect 26988 29306 27016 29990
rect 26976 29300 27028 29306
rect 26976 29242 27028 29248
rect 27080 28762 27108 31282
rect 27172 30977 27200 31282
rect 27356 31260 27384 31622
rect 27436 31272 27488 31278
rect 27356 31232 27436 31260
rect 27436 31214 27488 31220
rect 27712 31272 27764 31278
rect 27712 31214 27764 31220
rect 27158 30968 27214 30977
rect 27158 30903 27214 30912
rect 27724 30870 27752 31214
rect 27896 31204 27948 31210
rect 27896 31146 27948 31152
rect 27908 31113 27936 31146
rect 27894 31104 27950 31113
rect 27894 31039 27950 31048
rect 27802 30968 27858 30977
rect 27802 30903 27858 30912
rect 27816 30870 27844 30903
rect 27528 30864 27580 30870
rect 27342 30832 27398 30841
rect 27712 30864 27764 30870
rect 27528 30806 27580 30812
rect 27618 30832 27674 30841
rect 27342 30767 27398 30776
rect 27068 28756 27120 28762
rect 27068 28698 27120 28704
rect 27356 28694 27384 30767
rect 27540 30394 27568 30806
rect 27712 30806 27764 30812
rect 27804 30864 27856 30870
rect 27804 30806 27856 30812
rect 27618 30767 27674 30776
rect 27632 30734 27660 30767
rect 27620 30728 27672 30734
rect 27620 30670 27672 30676
rect 27528 30388 27580 30394
rect 27528 30330 27580 30336
rect 27436 29844 27488 29850
rect 27436 29786 27488 29792
rect 27448 29306 27476 29786
rect 27816 29782 27844 30806
rect 27908 30734 27936 31039
rect 27896 30728 27948 30734
rect 27896 30670 27948 30676
rect 27894 29880 27950 29889
rect 27894 29815 27950 29824
rect 27908 29782 27936 29815
rect 27804 29776 27856 29782
rect 27804 29718 27856 29724
rect 27896 29776 27948 29782
rect 27896 29718 27948 29724
rect 27528 29572 27580 29578
rect 27528 29514 27580 29520
rect 27436 29300 27488 29306
rect 27436 29242 27488 29248
rect 27540 29170 27568 29514
rect 27528 29164 27580 29170
rect 27528 29106 27580 29112
rect 27436 29096 27488 29102
rect 27436 29038 27488 29044
rect 27344 28688 27396 28694
rect 27344 28630 27396 28636
rect 27356 27470 27384 28630
rect 27448 28558 27476 29038
rect 27540 28626 27568 29106
rect 27528 28620 27580 28626
rect 27528 28562 27580 28568
rect 27436 28552 27488 28558
rect 27436 28494 27488 28500
rect 27540 27554 27568 28562
rect 27896 28552 27948 28558
rect 27896 28494 27948 28500
rect 27540 27526 27844 27554
rect 27908 27538 27936 28494
rect 27344 27464 27396 27470
rect 27344 27406 27396 27412
rect 27712 27464 27764 27470
rect 27712 27406 27764 27412
rect 26620 27084 26832 27112
rect 26516 24812 26568 24818
rect 26516 24754 26568 24760
rect 26424 24608 26476 24614
rect 26424 24550 26476 24556
rect 26528 24426 26556 24754
rect 26344 24398 26556 24426
rect 26344 22642 26372 24398
rect 26422 24304 26478 24313
rect 26422 24239 26478 24248
rect 26436 24138 26464 24239
rect 26424 24132 26476 24138
rect 26424 24074 26476 24080
rect 26436 23798 26464 24074
rect 26424 23792 26476 23798
rect 26424 23734 26476 23740
rect 26424 22772 26476 22778
rect 26424 22714 26476 22720
rect 26332 22636 26384 22642
rect 26332 22578 26384 22584
rect 26148 21888 26200 21894
rect 26148 21830 26200 21836
rect 26240 21888 26292 21894
rect 26240 21830 26292 21836
rect 26056 20052 26108 20058
rect 26056 19994 26108 20000
rect 25964 18760 26016 18766
rect 25962 18728 25964 18737
rect 26016 18728 26018 18737
rect 25962 18663 26018 18672
rect 25964 18624 26016 18630
rect 25964 18566 26016 18572
rect 25976 18306 26004 18566
rect 26054 18320 26110 18329
rect 25976 18278 26054 18306
rect 26054 18255 26056 18264
rect 26108 18255 26110 18264
rect 26056 18226 26108 18232
rect 26160 17921 26188 21830
rect 26240 21072 26292 21078
rect 26240 21014 26292 21020
rect 26252 19990 26280 21014
rect 26240 19984 26292 19990
rect 26240 19926 26292 19932
rect 26344 19378 26372 22578
rect 26436 20602 26464 22714
rect 26516 22568 26568 22574
rect 26516 22510 26568 22516
rect 26528 22234 26556 22510
rect 26516 22228 26568 22234
rect 26516 22170 26568 22176
rect 26424 20596 26476 20602
rect 26424 20538 26476 20544
rect 26528 19786 26556 22170
rect 26620 21350 26648 27084
rect 26792 26988 26844 26994
rect 26792 26930 26844 26936
rect 26804 26586 26832 26930
rect 26792 26580 26844 26586
rect 26792 26522 26844 26528
rect 26700 26444 26752 26450
rect 26700 26386 26752 26392
rect 27620 26444 27672 26450
rect 27620 26386 27672 26392
rect 26712 25401 26740 26386
rect 27068 26376 27120 26382
rect 27068 26318 27120 26324
rect 26698 25392 26754 25401
rect 26698 25327 26754 25336
rect 26974 25392 27030 25401
rect 26974 25327 26976 25336
rect 27028 25327 27030 25336
rect 26976 25298 27028 25304
rect 26700 25288 26752 25294
rect 26700 25230 26752 25236
rect 26884 25288 26936 25294
rect 26884 25230 26936 25236
rect 26712 24410 26740 25230
rect 26896 24750 26924 25230
rect 26976 24948 27028 24954
rect 26976 24890 27028 24896
rect 26884 24744 26936 24750
rect 26884 24686 26936 24692
rect 26988 24410 27016 24890
rect 27080 24750 27108 26318
rect 27632 25129 27660 26386
rect 27724 26382 27752 27406
rect 27816 26382 27844 27526
rect 27896 27532 27948 27538
rect 27896 27474 27948 27480
rect 28000 26518 28028 31894
rect 28092 31822 28120 32166
rect 28080 31816 28132 31822
rect 28080 31758 28132 31764
rect 28264 31816 28316 31822
rect 28264 31758 28316 31764
rect 28080 31680 28132 31686
rect 28080 31622 28132 31628
rect 28092 31142 28120 31622
rect 28276 31346 28304 31758
rect 28264 31340 28316 31346
rect 28264 31282 28316 31288
rect 28264 31204 28316 31210
rect 28264 31146 28316 31152
rect 28080 31136 28132 31142
rect 28080 31078 28132 31084
rect 28092 30326 28120 31078
rect 28172 30660 28224 30666
rect 28172 30602 28224 30608
rect 28080 30320 28132 30326
rect 28080 30262 28132 30268
rect 28184 28994 28212 30602
rect 28276 29730 28304 31146
rect 28368 30870 28396 33526
rect 28448 33448 28500 33454
rect 28448 33390 28500 33396
rect 28460 33114 28488 33390
rect 28448 33108 28500 33114
rect 28448 33050 28500 33056
rect 28448 32360 28500 32366
rect 28448 32302 28500 32308
rect 28460 31482 28488 32302
rect 28540 32292 28592 32298
rect 28540 32234 28592 32240
rect 28552 31822 28580 32234
rect 28644 31822 28672 34156
rect 28920 34066 28948 34546
rect 29000 34400 29052 34406
rect 29000 34342 29052 34348
rect 28908 34060 28960 34066
rect 28908 34002 28960 34008
rect 28920 33522 28948 34002
rect 29012 33590 29040 34342
rect 29920 34060 29972 34066
rect 29920 34002 29972 34008
rect 29736 33924 29788 33930
rect 29736 33866 29788 33872
rect 29748 33658 29776 33866
rect 29736 33652 29788 33658
rect 29736 33594 29788 33600
rect 29000 33584 29052 33590
rect 29000 33526 29052 33532
rect 28908 33516 28960 33522
rect 28908 33458 28960 33464
rect 29552 33516 29604 33522
rect 29552 33458 29604 33464
rect 29644 33516 29696 33522
rect 29644 33458 29696 33464
rect 29000 33448 29052 33454
rect 29000 33390 29052 33396
rect 28908 32972 28960 32978
rect 29012 32960 29040 33390
rect 29092 33380 29144 33386
rect 29092 33322 29144 33328
rect 28960 32932 29040 32960
rect 28908 32914 28960 32920
rect 29104 32910 29132 33322
rect 29460 33312 29512 33318
rect 29460 33254 29512 33260
rect 29472 32978 29500 33254
rect 29564 33114 29592 33458
rect 29552 33108 29604 33114
rect 29552 33050 29604 33056
rect 29550 33008 29606 33017
rect 29460 32972 29512 32978
rect 29550 32943 29606 32952
rect 29460 32914 29512 32920
rect 29564 32910 29592 32943
rect 28816 32904 28868 32910
rect 29092 32904 29144 32910
rect 28816 32846 28868 32852
rect 28906 32872 28962 32881
rect 28828 32774 28856 32846
rect 29092 32846 29144 32852
rect 29552 32904 29604 32910
rect 29552 32846 29604 32852
rect 28906 32807 28962 32816
rect 28816 32768 28868 32774
rect 28920 32756 28948 32807
rect 28920 32728 29040 32756
rect 28816 32710 28868 32716
rect 29012 32570 29040 32728
rect 28908 32564 28960 32570
rect 28908 32506 28960 32512
rect 29000 32564 29052 32570
rect 29000 32506 29052 32512
rect 28816 32428 28868 32434
rect 28816 32370 28868 32376
rect 28828 31822 28856 32370
rect 28540 31816 28592 31822
rect 28540 31758 28592 31764
rect 28632 31816 28684 31822
rect 28632 31758 28684 31764
rect 28816 31816 28868 31822
rect 28816 31758 28868 31764
rect 28920 31782 28948 32506
rect 29012 31958 29040 32506
rect 29092 32428 29144 32434
rect 29092 32370 29144 32376
rect 29104 32337 29132 32370
rect 29368 32360 29420 32366
rect 29090 32328 29146 32337
rect 29368 32302 29420 32308
rect 29090 32263 29146 32272
rect 29380 32065 29408 32302
rect 29366 32056 29422 32065
rect 29366 31991 29422 32000
rect 29000 31952 29052 31958
rect 29000 31894 29052 31900
rect 29092 31884 29144 31890
rect 29092 31826 29144 31832
rect 29000 31816 29052 31822
rect 28920 31764 29000 31782
rect 28920 31758 29052 31764
rect 28552 31657 28580 31758
rect 28644 31686 28672 31758
rect 28632 31680 28684 31686
rect 28538 31648 28594 31657
rect 28632 31622 28684 31628
rect 28538 31583 28594 31592
rect 28448 31476 28500 31482
rect 28500 31436 28580 31464
rect 28448 31418 28500 31424
rect 28446 31376 28502 31385
rect 28446 31311 28448 31320
rect 28500 31311 28502 31320
rect 28448 31282 28500 31288
rect 28356 30864 28408 30870
rect 28356 30806 28408 30812
rect 28276 29702 28488 29730
rect 28552 29714 28580 31436
rect 28828 31414 28856 31758
rect 28920 31754 29040 31758
rect 28816 31408 28868 31414
rect 28816 31350 28868 31356
rect 28816 31272 28868 31278
rect 28816 31214 28868 31220
rect 28724 31136 28776 31142
rect 28724 31078 28776 31084
rect 28632 30796 28684 30802
rect 28632 30738 28684 30744
rect 28644 30666 28672 30738
rect 28632 30660 28684 30666
rect 28632 30602 28684 30608
rect 28276 29646 28304 29702
rect 28264 29640 28316 29646
rect 28264 29582 28316 29588
rect 28356 29640 28408 29646
rect 28356 29582 28408 29588
rect 28264 29504 28316 29510
rect 28264 29446 28316 29452
rect 28276 29170 28304 29446
rect 28368 29170 28396 29582
rect 28460 29170 28488 29702
rect 28540 29708 28592 29714
rect 28540 29650 28592 29656
rect 28540 29572 28592 29578
rect 28540 29514 28592 29520
rect 28552 29238 28580 29514
rect 28540 29232 28592 29238
rect 28540 29174 28592 29180
rect 28264 29164 28316 29170
rect 28264 29106 28316 29112
rect 28356 29164 28408 29170
rect 28356 29106 28408 29112
rect 28448 29164 28500 29170
rect 28448 29106 28500 29112
rect 28460 29050 28488 29106
rect 28092 28966 28212 28994
rect 28368 29022 28488 29050
rect 28092 27470 28120 28966
rect 28264 28960 28316 28966
rect 28264 28902 28316 28908
rect 28276 28558 28304 28902
rect 28264 28552 28316 28558
rect 28264 28494 28316 28500
rect 28172 27532 28224 27538
rect 28172 27474 28224 27480
rect 28080 27464 28132 27470
rect 28080 27406 28132 27412
rect 27988 26512 28040 26518
rect 27988 26454 28040 26460
rect 28184 26450 28212 27474
rect 28276 26772 28304 28494
rect 28368 26840 28396 29022
rect 28552 28422 28580 29174
rect 28540 28416 28592 28422
rect 28540 28358 28592 28364
rect 28644 27062 28672 30602
rect 28736 29102 28764 31078
rect 28724 29096 28776 29102
rect 28724 29038 28776 29044
rect 28828 29034 28856 31214
rect 28908 30864 28960 30870
rect 28908 30806 28960 30812
rect 28920 30326 28948 30806
rect 29000 30728 29052 30734
rect 29000 30670 29052 30676
rect 29012 30433 29040 30670
rect 28998 30424 29054 30433
rect 28998 30359 29054 30368
rect 28908 30320 28960 30326
rect 28908 30262 28960 30268
rect 28816 29028 28868 29034
rect 28816 28970 28868 28976
rect 28828 28558 28856 28970
rect 28816 28552 28868 28558
rect 28816 28494 28868 28500
rect 28724 27464 28776 27470
rect 28724 27406 28776 27412
rect 28632 27056 28684 27062
rect 28632 26998 28684 27004
rect 28368 26812 28488 26840
rect 28276 26744 28396 26772
rect 28172 26444 28224 26450
rect 28172 26386 28224 26392
rect 27712 26376 27764 26382
rect 27804 26376 27856 26382
rect 27712 26318 27764 26324
rect 27802 26344 27804 26353
rect 27896 26376 27948 26382
rect 27856 26344 27858 26353
rect 27724 26228 27752 26318
rect 27896 26318 27948 26324
rect 27988 26376 28040 26382
rect 27988 26318 28040 26324
rect 27802 26279 27858 26288
rect 27724 26200 27844 26228
rect 27908 26217 27936 26318
rect 27618 25120 27674 25129
rect 27618 25055 27674 25064
rect 27252 24812 27304 24818
rect 27252 24754 27304 24760
rect 27436 24812 27488 24818
rect 27436 24754 27488 24760
rect 27068 24744 27120 24750
rect 27068 24686 27120 24692
rect 27160 24676 27212 24682
rect 27160 24618 27212 24624
rect 26700 24404 26752 24410
rect 26700 24346 26752 24352
rect 26976 24404 27028 24410
rect 26976 24346 27028 24352
rect 26712 24206 26740 24346
rect 27172 24290 27200 24618
rect 26896 24262 27200 24290
rect 27264 24274 27292 24754
rect 27344 24608 27396 24614
rect 27344 24550 27396 24556
rect 27356 24410 27384 24550
rect 27344 24404 27396 24410
rect 27344 24346 27396 24352
rect 27252 24268 27304 24274
rect 26700 24200 26752 24206
rect 26700 24142 26752 24148
rect 26700 23656 26752 23662
rect 26700 23598 26752 23604
rect 26712 21690 26740 23598
rect 26792 22636 26844 22642
rect 26792 22578 26844 22584
rect 26700 21684 26752 21690
rect 26700 21626 26752 21632
rect 26608 21344 26660 21350
rect 26608 21286 26660 21292
rect 26608 20800 26660 20806
rect 26608 20742 26660 20748
rect 26620 19854 26648 20742
rect 26700 20460 26752 20466
rect 26700 20402 26752 20408
rect 26712 20058 26740 20402
rect 26700 20052 26752 20058
rect 26700 19994 26752 20000
rect 26608 19848 26660 19854
rect 26608 19790 26660 19796
rect 26516 19780 26568 19786
rect 26516 19722 26568 19728
rect 26332 19372 26384 19378
rect 26332 19314 26384 19320
rect 26528 18970 26556 19722
rect 26516 18964 26568 18970
rect 26516 18906 26568 18912
rect 26240 18896 26292 18902
rect 26240 18838 26292 18844
rect 26252 18154 26280 18838
rect 26516 18284 26568 18290
rect 26516 18226 26568 18232
rect 26240 18148 26292 18154
rect 26240 18090 26292 18096
rect 26424 18080 26476 18086
rect 26424 18022 26476 18028
rect 26146 17912 26202 17921
rect 26436 17882 26464 18022
rect 26146 17847 26202 17856
rect 26424 17876 26476 17882
rect 26424 17818 26476 17824
rect 26146 17776 26202 17785
rect 26146 17711 26202 17720
rect 26056 16584 26108 16590
rect 26056 16526 26108 16532
rect 25872 16244 25924 16250
rect 25872 16186 25924 16192
rect 25872 14408 25924 14414
rect 25872 14350 25924 14356
rect 25964 14408 26016 14414
rect 25964 14350 26016 14356
rect 25884 13190 25912 14350
rect 25976 14074 26004 14350
rect 25964 14068 26016 14074
rect 25964 14010 26016 14016
rect 26068 13954 26096 16526
rect 25976 13926 26096 13954
rect 25872 13184 25924 13190
rect 25872 13126 25924 13132
rect 25976 12918 26004 13926
rect 26056 13864 26108 13870
rect 26056 13806 26108 13812
rect 25964 12912 26016 12918
rect 25964 12854 26016 12860
rect 25872 12640 25924 12646
rect 25872 12582 25924 12588
rect 25884 11558 25912 12582
rect 26068 12238 26096 13806
rect 26160 13326 26188 17711
rect 26424 16584 26476 16590
rect 26424 16526 26476 16532
rect 26436 16250 26464 16526
rect 26332 16244 26384 16250
rect 26332 16186 26384 16192
rect 26424 16244 26476 16250
rect 26424 16186 26476 16192
rect 26240 15496 26292 15502
rect 26240 15438 26292 15444
rect 26252 14006 26280 15438
rect 26240 14000 26292 14006
rect 26240 13942 26292 13948
rect 26252 13326 26280 13942
rect 26344 13530 26372 16186
rect 26424 15428 26476 15434
rect 26424 15370 26476 15376
rect 26436 14278 26464 15370
rect 26424 14272 26476 14278
rect 26528 14249 26556 18226
rect 26620 17882 26648 19790
rect 26608 17876 26660 17882
rect 26608 17818 26660 17824
rect 26712 16794 26740 19994
rect 26804 18970 26832 22578
rect 26792 18964 26844 18970
rect 26792 18906 26844 18912
rect 26792 18216 26844 18222
rect 26792 18158 26844 18164
rect 26700 16788 26752 16794
rect 26700 16730 26752 16736
rect 26804 15348 26832 18158
rect 26896 17678 26924 24262
rect 27252 24210 27304 24216
rect 27448 24070 27476 24754
rect 27528 24608 27580 24614
rect 27528 24550 27580 24556
rect 27540 24342 27568 24550
rect 27528 24336 27580 24342
rect 27528 24278 27580 24284
rect 27528 24200 27580 24206
rect 27712 24200 27764 24206
rect 27580 24160 27660 24188
rect 27528 24142 27580 24148
rect 27436 24064 27488 24070
rect 27436 24006 27488 24012
rect 27528 24064 27580 24070
rect 27528 24006 27580 24012
rect 27252 23792 27304 23798
rect 27252 23734 27304 23740
rect 27068 22500 27120 22506
rect 27068 22442 27120 22448
rect 27080 22030 27108 22442
rect 27160 22228 27212 22234
rect 27160 22170 27212 22176
rect 27068 22024 27120 22030
rect 27068 21966 27120 21972
rect 26976 21888 27028 21894
rect 26976 21830 27028 21836
rect 26988 18086 27016 21830
rect 27080 21622 27108 21966
rect 27068 21616 27120 21622
rect 27068 21558 27120 21564
rect 27068 20392 27120 20398
rect 27068 20334 27120 20340
rect 27080 19417 27108 20334
rect 27172 19786 27200 22170
rect 27264 21554 27292 23734
rect 27540 22778 27568 24006
rect 27632 23100 27660 24160
rect 27712 24142 27764 24148
rect 27724 23866 27752 24142
rect 27712 23860 27764 23866
rect 27712 23802 27764 23808
rect 27816 23254 27844 26200
rect 27894 26208 27950 26217
rect 27894 26143 27950 26152
rect 28000 25770 28028 26318
rect 27988 25764 28040 25770
rect 27988 25706 28040 25712
rect 28184 24614 28212 26386
rect 28264 26240 28316 26246
rect 28264 26182 28316 26188
rect 28276 26042 28304 26182
rect 28264 26036 28316 26042
rect 28264 25978 28316 25984
rect 28368 25106 28396 26744
rect 28460 26500 28488 26812
rect 28540 26512 28592 26518
rect 28460 26472 28540 26500
rect 28540 26454 28592 26460
rect 28448 26376 28500 26382
rect 28448 26318 28500 26324
rect 28460 25430 28488 26318
rect 28552 25974 28580 26454
rect 28632 26308 28684 26314
rect 28632 26250 28684 26256
rect 28644 26217 28672 26250
rect 28630 26208 28686 26217
rect 28630 26143 28686 26152
rect 28540 25968 28592 25974
rect 28540 25910 28592 25916
rect 28448 25424 28500 25430
rect 28448 25366 28500 25372
rect 28276 25078 28396 25106
rect 27988 24608 28040 24614
rect 27988 24550 28040 24556
rect 28172 24608 28224 24614
rect 28172 24550 28224 24556
rect 28000 24274 28028 24550
rect 28184 24313 28212 24550
rect 28170 24304 28226 24313
rect 27988 24268 28040 24274
rect 28170 24239 28226 24248
rect 27988 24210 28040 24216
rect 28080 24200 28132 24206
rect 28080 24142 28132 24148
rect 27986 23896 28042 23905
rect 27986 23831 28042 23840
rect 28000 23730 28028 23831
rect 27988 23724 28040 23730
rect 27988 23666 28040 23672
rect 27804 23248 27856 23254
rect 27804 23190 27856 23196
rect 27632 23072 27844 23100
rect 27712 22976 27764 22982
rect 27712 22918 27764 22924
rect 27528 22772 27580 22778
rect 27528 22714 27580 22720
rect 27620 22772 27672 22778
rect 27620 22714 27672 22720
rect 27632 22522 27660 22714
rect 27448 22494 27660 22522
rect 27344 22432 27396 22438
rect 27344 22374 27396 22380
rect 27356 22234 27384 22374
rect 27344 22228 27396 22234
rect 27344 22170 27396 22176
rect 27448 21842 27476 22494
rect 27620 22432 27672 22438
rect 27620 22374 27672 22380
rect 27632 22094 27660 22374
rect 27540 22066 27660 22094
rect 27540 22030 27568 22066
rect 27528 22024 27580 22030
rect 27724 21978 27752 22918
rect 27816 22137 27844 23072
rect 28092 22438 28120 24142
rect 28276 24041 28304 25078
rect 28540 24812 28592 24818
rect 28540 24754 28592 24760
rect 28448 24608 28500 24614
rect 28448 24550 28500 24556
rect 28356 24404 28408 24410
rect 28356 24346 28408 24352
rect 28262 24032 28318 24041
rect 28262 23967 28318 23976
rect 28172 23588 28224 23594
rect 28172 23530 28224 23536
rect 28184 22506 28212 23530
rect 28172 22500 28224 22506
rect 28172 22442 28224 22448
rect 28080 22432 28132 22438
rect 28276 22386 28304 23967
rect 28368 23730 28396 24346
rect 28460 24206 28488 24550
rect 28552 24313 28580 24754
rect 28538 24304 28594 24313
rect 28736 24274 28764 27406
rect 28816 26376 28868 26382
rect 28814 26344 28816 26353
rect 28868 26344 28870 26353
rect 28814 26279 28870 26288
rect 29000 25696 29052 25702
rect 29000 25638 29052 25644
rect 29012 25362 29040 25638
rect 29000 25356 29052 25362
rect 29000 25298 29052 25304
rect 28908 24744 28960 24750
rect 28908 24686 28960 24692
rect 28538 24239 28594 24248
rect 28724 24268 28776 24274
rect 28724 24210 28776 24216
rect 28448 24200 28500 24206
rect 28448 24142 28500 24148
rect 28540 24200 28592 24206
rect 28540 24142 28592 24148
rect 28460 23769 28488 24142
rect 28446 23760 28502 23769
rect 28356 23724 28408 23730
rect 28552 23730 28580 24142
rect 28632 24132 28684 24138
rect 28632 24074 28684 24080
rect 28446 23695 28502 23704
rect 28540 23724 28592 23730
rect 28356 23666 28408 23672
rect 28540 23666 28592 23672
rect 28368 22982 28396 23666
rect 28356 22976 28408 22982
rect 28356 22918 28408 22924
rect 28644 22642 28672 24074
rect 28736 23866 28764 24210
rect 28724 23860 28776 23866
rect 28724 23802 28776 23808
rect 28920 23730 28948 24686
rect 29000 24200 29052 24206
rect 29000 24142 29052 24148
rect 29012 23866 29040 24142
rect 29000 23860 29052 23866
rect 29000 23802 29052 23808
rect 28724 23724 28776 23730
rect 28724 23666 28776 23672
rect 28908 23724 28960 23730
rect 28908 23666 28960 23672
rect 28448 22636 28500 22642
rect 28448 22578 28500 22584
rect 28632 22636 28684 22642
rect 28632 22578 28684 22584
rect 28460 22438 28488 22578
rect 28736 22574 28764 23666
rect 28920 23594 28948 23666
rect 28908 23588 28960 23594
rect 28908 23530 28960 23536
rect 28816 23520 28868 23526
rect 28816 23462 28868 23468
rect 28724 22568 28776 22574
rect 28724 22510 28776 22516
rect 28080 22374 28132 22380
rect 28184 22358 28304 22386
rect 28448 22432 28500 22438
rect 28448 22374 28500 22380
rect 27802 22128 27858 22137
rect 27802 22063 27858 22072
rect 27528 21966 27580 21972
rect 27356 21814 27476 21842
rect 27356 21554 27384 21814
rect 27252 21548 27304 21554
rect 27252 21490 27304 21496
rect 27344 21548 27396 21554
rect 27344 21490 27396 21496
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 27436 20460 27488 20466
rect 27540 20448 27568 21966
rect 27632 21962 27752 21978
rect 27620 21956 27752 21962
rect 27672 21950 27752 21956
rect 27620 21898 27672 21904
rect 27632 20874 27660 21898
rect 27896 21616 27948 21622
rect 27896 21558 27948 21564
rect 27986 21584 28042 21593
rect 27712 21548 27764 21554
rect 27712 21490 27764 21496
rect 27724 20874 27752 21490
rect 27620 20868 27672 20874
rect 27620 20810 27672 20816
rect 27712 20868 27764 20874
rect 27712 20810 27764 20816
rect 27618 20632 27674 20641
rect 27618 20567 27674 20576
rect 27488 20420 27568 20448
rect 27436 20402 27488 20408
rect 27250 20360 27306 20369
rect 27250 20295 27306 20304
rect 27264 19854 27292 20295
rect 27252 19848 27304 19854
rect 27252 19790 27304 19796
rect 27160 19780 27212 19786
rect 27160 19722 27212 19728
rect 27066 19408 27122 19417
rect 27066 19343 27122 19352
rect 27080 18290 27108 19343
rect 27172 18426 27200 19722
rect 27356 19514 27384 20402
rect 27252 19508 27304 19514
rect 27252 19450 27304 19456
rect 27344 19508 27396 19514
rect 27344 19450 27396 19456
rect 27264 19174 27292 19450
rect 27252 19168 27304 19174
rect 27252 19110 27304 19116
rect 27448 18970 27476 20402
rect 27528 20324 27580 20330
rect 27528 20266 27580 20272
rect 27540 20233 27568 20266
rect 27526 20224 27582 20233
rect 27526 20159 27582 20168
rect 27528 19848 27580 19854
rect 27528 19790 27580 19796
rect 27540 19428 27568 19790
rect 27632 19768 27660 20567
rect 27712 20460 27764 20466
rect 27712 20402 27764 20408
rect 27724 20058 27752 20402
rect 27804 20392 27856 20398
rect 27804 20334 27856 20340
rect 27816 20262 27844 20334
rect 27804 20256 27856 20262
rect 27804 20198 27856 20204
rect 27712 20052 27764 20058
rect 27712 19994 27764 20000
rect 27908 19854 27936 21558
rect 27986 21519 27988 21528
rect 28040 21519 28042 21528
rect 27988 21490 28040 21496
rect 27988 21344 28040 21350
rect 27988 21286 28040 21292
rect 28000 20262 28028 21286
rect 28080 20392 28132 20398
rect 28080 20334 28132 20340
rect 27988 20256 28040 20262
rect 27988 20198 28040 20204
rect 27896 19848 27948 19854
rect 27896 19790 27948 19796
rect 27712 19780 27764 19786
rect 27632 19740 27712 19768
rect 27712 19722 27764 19728
rect 27988 19780 28040 19786
rect 27988 19722 28040 19728
rect 27620 19440 27672 19446
rect 27540 19400 27620 19428
rect 27436 18964 27488 18970
rect 27436 18906 27488 18912
rect 27250 18728 27306 18737
rect 27250 18663 27306 18672
rect 27160 18420 27212 18426
rect 27160 18362 27212 18368
rect 27068 18284 27120 18290
rect 27068 18226 27120 18232
rect 27264 18222 27292 18663
rect 27436 18624 27488 18630
rect 27434 18592 27436 18601
rect 27488 18592 27490 18601
rect 27434 18527 27490 18536
rect 27448 18426 27476 18527
rect 27436 18420 27488 18426
rect 27436 18362 27488 18368
rect 27252 18216 27304 18222
rect 27252 18158 27304 18164
rect 26976 18080 27028 18086
rect 26976 18022 27028 18028
rect 26884 17672 26936 17678
rect 26884 17614 26936 17620
rect 27160 17536 27212 17542
rect 27160 17478 27212 17484
rect 27252 17536 27304 17542
rect 27252 17478 27304 17484
rect 27172 17202 27200 17478
rect 27264 17338 27292 17478
rect 27252 17332 27304 17338
rect 27252 17274 27304 17280
rect 27344 17332 27396 17338
rect 27344 17274 27396 17280
rect 27160 17196 27212 17202
rect 27160 17138 27212 17144
rect 27356 16697 27384 17274
rect 27342 16688 27398 16697
rect 27342 16623 27398 16632
rect 27540 16561 27568 19400
rect 27620 19382 27672 19388
rect 27804 19440 27856 19446
rect 27804 19382 27856 19388
rect 27710 19272 27766 19281
rect 27710 19207 27712 19216
rect 27764 19207 27766 19216
rect 27712 19178 27764 19184
rect 27620 18964 27672 18970
rect 27620 18906 27672 18912
rect 27632 18766 27660 18906
rect 27816 18902 27844 19382
rect 27804 18896 27856 18902
rect 27804 18838 27856 18844
rect 27620 18760 27672 18766
rect 27620 18702 27672 18708
rect 27896 18760 27948 18766
rect 27896 18702 27948 18708
rect 27632 18329 27660 18702
rect 27618 18320 27674 18329
rect 27618 18255 27674 18264
rect 27712 18284 27764 18290
rect 27632 18086 27660 18255
rect 27712 18226 27764 18232
rect 27620 18080 27672 18086
rect 27620 18022 27672 18028
rect 27618 17912 27674 17921
rect 27618 17847 27674 17856
rect 27632 17490 27660 17847
rect 27724 17610 27752 18226
rect 27712 17604 27764 17610
rect 27712 17546 27764 17552
rect 27632 17462 27752 17490
rect 27526 16552 27582 16561
rect 27526 16487 27582 16496
rect 27436 16448 27488 16454
rect 27436 16390 27488 16396
rect 27448 16114 27476 16390
rect 27540 16182 27568 16487
rect 27528 16176 27580 16182
rect 27580 16136 27660 16164
rect 27528 16118 27580 16124
rect 27436 16108 27488 16114
rect 27436 16050 27488 16056
rect 27252 15972 27304 15978
rect 27252 15914 27304 15920
rect 27264 15706 27292 15914
rect 27252 15700 27304 15706
rect 27252 15642 27304 15648
rect 26804 15320 26924 15348
rect 26608 14272 26660 14278
rect 26424 14214 26476 14220
rect 26514 14240 26570 14249
rect 26608 14214 26660 14220
rect 26514 14175 26570 14184
rect 26620 14090 26648 14214
rect 26436 14062 26648 14090
rect 26700 14068 26752 14074
rect 26332 13524 26384 13530
rect 26332 13466 26384 13472
rect 26148 13320 26200 13326
rect 26240 13320 26292 13326
rect 26148 13262 26200 13268
rect 26238 13288 26240 13297
rect 26292 13288 26294 13297
rect 26238 13223 26294 13232
rect 26436 12594 26464 14062
rect 26700 14010 26752 14016
rect 26712 13870 26740 14010
rect 26516 13864 26568 13870
rect 26516 13806 26568 13812
rect 26700 13864 26752 13870
rect 26700 13806 26752 13812
rect 26528 13308 26556 13806
rect 26608 13320 26660 13326
rect 26528 13280 26608 13308
rect 26608 13262 26660 13268
rect 26516 12912 26568 12918
rect 26516 12854 26568 12860
rect 26252 12566 26464 12594
rect 26056 12232 26108 12238
rect 26056 12174 26108 12180
rect 25964 11824 26016 11830
rect 26068 11812 26096 12174
rect 26016 11784 26096 11812
rect 25964 11766 26016 11772
rect 26252 11762 26280 12566
rect 26332 12232 26384 12238
rect 26332 12174 26384 12180
rect 26344 11830 26372 12174
rect 26424 12164 26476 12170
rect 26424 12106 26476 12112
rect 26332 11824 26384 11830
rect 26332 11766 26384 11772
rect 26240 11756 26292 11762
rect 26240 11698 26292 11704
rect 26056 11688 26108 11694
rect 26056 11630 26108 11636
rect 25964 11620 26016 11626
rect 25964 11562 26016 11568
rect 25872 11552 25924 11558
rect 25872 11494 25924 11500
rect 25596 10056 25648 10062
rect 25594 10024 25596 10033
rect 25648 10024 25650 10033
rect 25594 9959 25650 9968
rect 25596 9648 25648 9654
rect 25502 9616 25558 9625
rect 25596 9590 25648 9596
rect 25502 9551 25558 9560
rect 25228 9376 25280 9382
rect 25228 9318 25280 9324
rect 25412 9376 25464 9382
rect 25412 9318 25464 9324
rect 25148 9178 25360 9194
rect 25044 9172 25096 9178
rect 25044 9114 25096 9120
rect 25148 9172 25372 9178
rect 25148 9166 25320 9172
rect 25148 9110 25176 9166
rect 25320 9114 25372 9120
rect 25136 9104 25188 9110
rect 25042 9072 25098 9081
rect 25516 9058 25544 9551
rect 25136 9046 25188 9052
rect 25042 9007 25098 9016
rect 25424 9030 25544 9058
rect 25056 8974 25084 9007
rect 25424 8974 25452 9030
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 25412 8968 25464 8974
rect 25412 8910 25464 8916
rect 25320 8900 25372 8906
rect 25320 8842 25372 8848
rect 25228 8832 25280 8838
rect 24950 8800 25006 8809
rect 25228 8774 25280 8780
rect 24950 8735 25006 8744
rect 24964 8634 24992 8735
rect 24952 8628 25004 8634
rect 24952 8570 25004 8576
rect 25240 8498 25268 8774
rect 25228 8492 25280 8498
rect 25228 8434 25280 8440
rect 25044 7744 25096 7750
rect 25044 7686 25096 7692
rect 25056 7546 25084 7686
rect 25044 7540 25096 7546
rect 25044 7482 25096 7488
rect 25332 7342 25360 8842
rect 25504 8084 25556 8090
rect 25504 8026 25556 8032
rect 25320 7336 25372 7342
rect 25320 7278 25372 7284
rect 24952 6860 25004 6866
rect 24952 6802 25004 6808
rect 24964 6322 24992 6802
rect 25332 6662 25360 7278
rect 25516 7206 25544 8026
rect 25504 7200 25556 7206
rect 25504 7142 25556 7148
rect 25320 6656 25372 6662
rect 25320 6598 25372 6604
rect 24952 6316 25004 6322
rect 24952 6258 25004 6264
rect 25412 6316 25464 6322
rect 25412 6258 25464 6264
rect 25136 6112 25188 6118
rect 25136 6054 25188 6060
rect 24860 5840 24912 5846
rect 24860 5782 24912 5788
rect 24952 5840 25004 5846
rect 24952 5782 25004 5788
rect 24584 5636 24636 5642
rect 24584 5578 24636 5584
rect 24768 5636 24820 5642
rect 24768 5578 24820 5584
rect 24216 5296 24268 5302
rect 24216 5238 24268 5244
rect 23940 5228 23992 5234
rect 23940 5170 23992 5176
rect 23952 4214 23980 5170
rect 24596 4570 24624 5578
rect 24872 5302 24900 5782
rect 24964 5574 24992 5782
rect 25148 5710 25176 6054
rect 25424 5846 25452 6258
rect 25608 6186 25636 9590
rect 25700 9518 25728 10118
rect 25780 10124 25832 10130
rect 25780 10066 25832 10072
rect 25688 9512 25740 9518
rect 25688 9454 25740 9460
rect 25976 9382 26004 11562
rect 26068 11354 26096 11630
rect 26240 11552 26292 11558
rect 26240 11494 26292 11500
rect 26056 11348 26108 11354
rect 26056 11290 26108 11296
rect 26054 10840 26110 10849
rect 26054 10775 26056 10784
rect 26108 10775 26110 10784
rect 26056 10746 26108 10752
rect 26056 10668 26108 10674
rect 26056 10610 26108 10616
rect 26068 9874 26096 10610
rect 26252 9994 26280 11494
rect 26344 11150 26372 11766
rect 26436 11762 26464 12106
rect 26424 11756 26476 11762
rect 26424 11698 26476 11704
rect 26332 11144 26384 11150
rect 26332 11086 26384 11092
rect 26240 9988 26292 9994
rect 26240 9930 26292 9936
rect 26148 9920 26200 9926
rect 26068 9868 26148 9874
rect 26068 9862 26200 9868
rect 26068 9846 26188 9862
rect 25964 9376 26016 9382
rect 25964 9318 26016 9324
rect 26160 9178 26188 9846
rect 26240 9376 26292 9382
rect 26240 9318 26292 9324
rect 26252 9178 26280 9318
rect 26148 9172 26200 9178
rect 26148 9114 26200 9120
rect 26240 9172 26292 9178
rect 26240 9114 26292 9120
rect 26056 8968 26108 8974
rect 26056 8910 26108 8916
rect 25688 8832 25740 8838
rect 25688 8774 25740 8780
rect 25700 8498 25728 8774
rect 25688 8492 25740 8498
rect 25688 8434 25740 8440
rect 25780 8492 25832 8498
rect 25780 8434 25832 8440
rect 25792 7954 25820 8434
rect 26068 8090 26096 8910
rect 26160 8566 26188 9114
rect 26240 9036 26292 9042
rect 26240 8978 26292 8984
rect 26148 8560 26200 8566
rect 26148 8502 26200 8508
rect 26056 8084 26108 8090
rect 26056 8026 26108 8032
rect 26252 7954 26280 8978
rect 26344 8974 26372 11086
rect 26436 11082 26464 11698
rect 26528 11626 26556 12854
rect 26516 11620 26568 11626
rect 26516 11562 26568 11568
rect 26424 11076 26476 11082
rect 26424 11018 26476 11024
rect 26424 10736 26476 10742
rect 26424 10678 26476 10684
rect 26436 10062 26464 10678
rect 26620 10266 26648 13262
rect 26792 12912 26844 12918
rect 26792 12854 26844 12860
rect 26804 11354 26832 12854
rect 26896 12434 26924 15320
rect 27448 15065 27476 16050
rect 27528 15904 27580 15910
rect 27528 15846 27580 15852
rect 27434 15056 27490 15065
rect 27434 14991 27490 15000
rect 27252 14544 27304 14550
rect 27252 14486 27304 14492
rect 27066 14104 27122 14113
rect 27066 14039 27068 14048
rect 27120 14039 27122 14048
rect 27068 14010 27120 14016
rect 27264 14006 27292 14486
rect 27436 14408 27488 14414
rect 27436 14350 27488 14356
rect 27252 14000 27304 14006
rect 27252 13942 27304 13948
rect 27448 13938 27476 14350
rect 27436 13932 27488 13938
rect 27436 13874 27488 13880
rect 27252 13864 27304 13870
rect 27252 13806 27304 13812
rect 27160 13796 27212 13802
rect 27160 13738 27212 13744
rect 27172 13326 27200 13738
rect 27160 13320 27212 13326
rect 27160 13262 27212 13268
rect 26896 12406 27108 12434
rect 26882 11656 26938 11665
rect 26882 11591 26884 11600
rect 26936 11591 26938 11600
rect 26884 11562 26936 11568
rect 26792 11348 26844 11354
rect 26792 11290 26844 11296
rect 26804 11150 26832 11290
rect 26792 11144 26844 11150
rect 26792 11086 26844 11092
rect 26976 11144 27028 11150
rect 26976 11086 27028 11092
rect 26608 10260 26660 10266
rect 26608 10202 26660 10208
rect 26424 10056 26476 10062
rect 26424 9998 26476 10004
rect 26436 9518 26464 9998
rect 26514 9752 26570 9761
rect 26514 9687 26570 9696
rect 26424 9512 26476 9518
rect 26424 9454 26476 9460
rect 26436 9042 26464 9454
rect 26424 9036 26476 9042
rect 26424 8978 26476 8984
rect 26332 8968 26384 8974
rect 26332 8910 26384 8916
rect 26332 8832 26384 8838
rect 26528 8786 26556 9687
rect 26804 9654 26832 11086
rect 26884 9920 26936 9926
rect 26884 9862 26936 9868
rect 26792 9648 26844 9654
rect 26792 9590 26844 9596
rect 26896 9586 26924 9862
rect 26884 9580 26936 9586
rect 26884 9522 26936 9528
rect 26790 9208 26846 9217
rect 26896 9178 26924 9522
rect 26790 9143 26846 9152
rect 26884 9172 26936 9178
rect 26700 8900 26752 8906
rect 26700 8842 26752 8848
rect 26384 8780 26556 8786
rect 26332 8774 26556 8780
rect 26344 8758 26556 8774
rect 25780 7948 25832 7954
rect 25780 7890 25832 7896
rect 26240 7948 26292 7954
rect 26240 7890 26292 7896
rect 26344 7546 26372 8758
rect 26712 8498 26740 8842
rect 26700 8492 26752 8498
rect 26700 8434 26752 8440
rect 26424 8288 26476 8294
rect 26424 8230 26476 8236
rect 26436 8090 26464 8230
rect 26424 8084 26476 8090
rect 26424 8026 26476 8032
rect 26516 8084 26568 8090
rect 26516 8026 26568 8032
rect 26332 7540 26384 7546
rect 26332 7482 26384 7488
rect 26528 7410 26556 8026
rect 26804 8022 26832 9143
rect 26884 9114 26936 9120
rect 26988 8294 27016 11086
rect 27080 10010 27108 12406
rect 27172 10130 27200 13262
rect 27264 12850 27292 13806
rect 27252 12844 27304 12850
rect 27448 12832 27476 13874
rect 27540 13462 27568 15846
rect 27632 13954 27660 16136
rect 27724 16114 27752 17462
rect 27908 17377 27936 18702
rect 28000 18630 28028 19722
rect 27988 18624 28040 18630
rect 27988 18566 28040 18572
rect 28000 18290 28028 18566
rect 27988 18284 28040 18290
rect 27988 18226 28040 18232
rect 27988 18080 28040 18086
rect 27988 18022 28040 18028
rect 27894 17368 27950 17377
rect 27894 17303 27950 17312
rect 27804 17060 27856 17066
rect 27804 17002 27856 17008
rect 27712 16108 27764 16114
rect 27712 16050 27764 16056
rect 27712 14884 27764 14890
rect 27712 14826 27764 14832
rect 27724 14346 27752 14826
rect 27816 14618 27844 17002
rect 28000 16522 28028 18022
rect 28092 16794 28120 20334
rect 28184 18902 28212 22358
rect 28540 21888 28592 21894
rect 28540 21830 28592 21836
rect 28356 21344 28408 21350
rect 28356 21286 28408 21292
rect 28368 21010 28396 21286
rect 28356 21004 28408 21010
rect 28356 20946 28408 20952
rect 28356 20868 28408 20874
rect 28356 20810 28408 20816
rect 28264 20460 28316 20466
rect 28264 20402 28316 20408
rect 28276 19990 28304 20402
rect 28264 19984 28316 19990
rect 28264 19926 28316 19932
rect 28368 19334 28396 20810
rect 28448 20256 28500 20262
rect 28448 20198 28500 20204
rect 28460 19922 28488 20198
rect 28448 19916 28500 19922
rect 28448 19858 28500 19864
rect 28368 19306 28488 19334
rect 28264 19168 28316 19174
rect 28264 19110 28316 19116
rect 28172 18896 28224 18902
rect 28172 18838 28224 18844
rect 28184 18358 28212 18838
rect 28172 18352 28224 18358
rect 28172 18294 28224 18300
rect 28172 17196 28224 17202
rect 28172 17138 28224 17144
rect 28080 16788 28132 16794
rect 28080 16730 28132 16736
rect 28184 16658 28212 17138
rect 28276 16794 28304 19110
rect 28356 18692 28408 18698
rect 28356 18634 28408 18640
rect 28368 18601 28396 18634
rect 28354 18592 28410 18601
rect 28354 18527 28410 18536
rect 28460 17610 28488 19306
rect 28552 17882 28580 21830
rect 28736 20874 28764 22510
rect 28724 20868 28776 20874
rect 28724 20810 28776 20816
rect 28828 20806 28856 23462
rect 28908 23248 28960 23254
rect 28908 23190 28960 23196
rect 28920 22642 28948 23190
rect 28998 23080 29054 23089
rect 28998 23015 29054 23024
rect 29012 22642 29040 23015
rect 28908 22636 28960 22642
rect 28908 22578 28960 22584
rect 29000 22636 29052 22642
rect 29000 22578 29052 22584
rect 29000 21616 29052 21622
rect 28998 21584 29000 21593
rect 29052 21584 29054 21593
rect 29104 21554 29132 31826
rect 29656 31482 29684 33458
rect 29736 33108 29788 33114
rect 29736 33050 29788 33056
rect 29748 32570 29776 33050
rect 29932 32978 29960 34002
rect 30196 33992 30248 33998
rect 30196 33934 30248 33940
rect 30208 33658 30236 33934
rect 30484 33930 30512 36042
rect 31116 34740 31168 34746
rect 31116 34682 31168 34688
rect 30472 33924 30524 33930
rect 30524 33884 30604 33912
rect 30472 33866 30524 33872
rect 30196 33652 30248 33658
rect 30196 33594 30248 33600
rect 30104 33448 30156 33454
rect 30104 33390 30156 33396
rect 29920 32972 29972 32978
rect 29920 32914 29972 32920
rect 29736 32564 29788 32570
rect 29736 32506 29788 32512
rect 29920 32564 29972 32570
rect 29920 32506 29972 32512
rect 29736 32360 29788 32366
rect 29736 32302 29788 32308
rect 29644 31476 29696 31482
rect 29644 31418 29696 31424
rect 29276 31340 29328 31346
rect 29276 31282 29328 31288
rect 29288 30394 29316 31282
rect 29552 30728 29604 30734
rect 29552 30670 29604 30676
rect 29276 30388 29328 30394
rect 29276 30330 29328 30336
rect 29288 28490 29316 30330
rect 29564 30190 29592 30670
rect 29552 30184 29604 30190
rect 29552 30126 29604 30132
rect 29748 29306 29776 32302
rect 29932 30394 29960 32506
rect 30116 32298 30144 33390
rect 30196 32972 30248 32978
rect 30196 32914 30248 32920
rect 30208 32502 30236 32914
rect 30576 32881 30604 33884
rect 30748 33380 30800 33386
rect 30748 33322 30800 33328
rect 30562 32872 30618 32881
rect 30472 32836 30524 32842
rect 30562 32807 30618 32816
rect 30472 32778 30524 32784
rect 30288 32768 30340 32774
rect 30288 32710 30340 32716
rect 30196 32496 30248 32502
rect 30196 32438 30248 32444
rect 30012 32292 30064 32298
rect 30012 32234 30064 32240
rect 30104 32292 30156 32298
rect 30104 32234 30156 32240
rect 30024 31822 30052 32234
rect 30012 31816 30064 31822
rect 30012 31758 30064 31764
rect 30104 30660 30156 30666
rect 30104 30602 30156 30608
rect 29920 30388 29972 30394
rect 29920 30330 29972 30336
rect 29736 29300 29788 29306
rect 29736 29242 29788 29248
rect 29644 28756 29696 28762
rect 29644 28698 29696 28704
rect 29276 28484 29328 28490
rect 29276 28426 29328 28432
rect 29184 28416 29236 28422
rect 29184 28358 29236 28364
rect 29196 28014 29224 28358
rect 29184 28008 29236 28014
rect 29184 27950 29236 27956
rect 29288 26568 29316 28426
rect 29656 27470 29684 28698
rect 29748 28558 29776 29242
rect 29920 28756 29972 28762
rect 29920 28698 29972 28704
rect 29932 28558 29960 28698
rect 29736 28552 29788 28558
rect 29736 28494 29788 28500
rect 29920 28552 29972 28558
rect 29920 28494 29972 28500
rect 29748 27538 29776 28494
rect 29828 28484 29880 28490
rect 29828 28426 29880 28432
rect 30012 28484 30064 28490
rect 30012 28426 30064 28432
rect 29840 28098 29868 28426
rect 29840 28070 29960 28098
rect 29932 27878 29960 28070
rect 29920 27872 29972 27878
rect 29920 27814 29972 27820
rect 29736 27532 29788 27538
rect 29736 27474 29788 27480
rect 29644 27464 29696 27470
rect 29644 27406 29696 27412
rect 29932 26858 29960 27814
rect 30024 27130 30052 28426
rect 30116 28150 30144 30602
rect 30208 30190 30236 32438
rect 30300 31754 30328 32710
rect 30484 32026 30512 32778
rect 30472 32020 30524 32026
rect 30472 31962 30524 31968
rect 30300 31726 30512 31754
rect 30484 30802 30512 31726
rect 30472 30796 30524 30802
rect 30472 30738 30524 30744
rect 30380 30728 30432 30734
rect 30380 30670 30432 30676
rect 30288 30592 30340 30598
rect 30288 30534 30340 30540
rect 30300 30258 30328 30534
rect 30288 30252 30340 30258
rect 30288 30194 30340 30200
rect 30196 30184 30248 30190
rect 30196 30126 30248 30132
rect 30104 28144 30156 28150
rect 30104 28086 30156 28092
rect 30208 28014 30236 30126
rect 30392 29492 30420 30670
rect 30576 30666 30604 32807
rect 30654 31784 30710 31793
rect 30760 31754 30788 33322
rect 31024 33312 31076 33318
rect 31024 33254 31076 33260
rect 30932 32836 30984 32842
rect 30932 32778 30984 32784
rect 30944 32745 30972 32778
rect 30930 32736 30986 32745
rect 30930 32671 30986 32680
rect 30710 31728 30788 31754
rect 30654 31719 30656 31728
rect 30708 31726 30788 31728
rect 30708 31719 30710 31726
rect 30656 31690 30708 31696
rect 30748 31340 30800 31346
rect 30748 31282 30800 31288
rect 30840 31340 30892 31346
rect 30840 31282 30892 31288
rect 30760 30977 30788 31282
rect 30746 30968 30802 30977
rect 30746 30903 30802 30912
rect 30748 30728 30800 30734
rect 30746 30696 30748 30705
rect 30800 30696 30802 30705
rect 30564 30660 30616 30666
rect 30746 30631 30802 30640
rect 30564 30602 30616 30608
rect 30472 30252 30524 30258
rect 30472 30194 30524 30200
rect 30564 30252 30616 30258
rect 30564 30194 30616 30200
rect 30484 30161 30512 30194
rect 30470 30152 30526 30161
rect 30470 30087 30526 30096
rect 30470 29880 30526 29889
rect 30470 29815 30526 29824
rect 30484 29646 30512 29815
rect 30472 29640 30524 29646
rect 30472 29582 30524 29588
rect 30392 29464 30512 29492
rect 30380 29164 30432 29170
rect 30380 29106 30432 29112
rect 30286 29064 30342 29073
rect 30286 28999 30342 29008
rect 30196 28008 30248 28014
rect 30196 27950 30248 27956
rect 30300 27878 30328 28999
rect 30392 28422 30420 29106
rect 30380 28416 30432 28422
rect 30380 28358 30432 28364
rect 30104 27872 30156 27878
rect 30104 27814 30156 27820
rect 30288 27872 30340 27878
rect 30288 27814 30340 27820
rect 30012 27124 30064 27130
rect 30012 27066 30064 27072
rect 30012 26920 30064 26926
rect 30012 26862 30064 26868
rect 29920 26852 29972 26858
rect 29920 26794 29972 26800
rect 29734 26752 29790 26761
rect 29734 26687 29790 26696
rect 29748 26586 29776 26687
rect 29736 26580 29788 26586
rect 29288 26540 29408 26568
rect 29276 26444 29328 26450
rect 29276 26386 29328 26392
rect 29288 25906 29316 26386
rect 29380 26042 29408 26540
rect 29736 26522 29788 26528
rect 29932 26382 29960 26794
rect 29920 26376 29972 26382
rect 29920 26318 29972 26324
rect 29736 26308 29788 26314
rect 29736 26250 29788 26256
rect 29368 26036 29420 26042
rect 29368 25978 29420 25984
rect 29276 25900 29328 25906
rect 29276 25842 29328 25848
rect 29368 25900 29420 25906
rect 29368 25842 29420 25848
rect 29552 25900 29604 25906
rect 29552 25842 29604 25848
rect 29380 25809 29408 25842
rect 29366 25800 29422 25809
rect 29366 25735 29422 25744
rect 29184 23792 29236 23798
rect 29184 23734 29236 23740
rect 28998 21519 29054 21528
rect 29092 21548 29144 21554
rect 29012 21146 29040 21519
rect 29092 21490 29144 21496
rect 29000 21140 29052 21146
rect 29000 21082 29052 21088
rect 28908 20936 28960 20942
rect 28906 20904 28908 20913
rect 29092 20936 29144 20942
rect 28960 20904 28962 20913
rect 29092 20878 29144 20884
rect 28906 20839 28962 20848
rect 28816 20800 28868 20806
rect 28816 20742 28868 20748
rect 29000 20800 29052 20806
rect 29000 20742 29052 20748
rect 28724 20528 28776 20534
rect 28722 20496 28724 20505
rect 28776 20496 28778 20505
rect 29012 20466 29040 20742
rect 28722 20431 28778 20440
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 28632 20392 28684 20398
rect 28632 20334 28684 20340
rect 28644 18698 28672 20334
rect 28722 19952 28778 19961
rect 28722 19887 28778 19896
rect 28736 19718 28764 19887
rect 28908 19848 28960 19854
rect 28908 19790 28960 19796
rect 28724 19712 28776 19718
rect 28724 19654 28776 19660
rect 28724 19372 28776 19378
rect 28724 19314 28776 19320
rect 28736 18970 28764 19314
rect 28920 19009 28948 19790
rect 29000 19508 29052 19514
rect 29000 19450 29052 19456
rect 28906 19000 28962 19009
rect 28724 18964 28776 18970
rect 28906 18935 28962 18944
rect 28724 18906 28776 18912
rect 29012 18766 29040 19450
rect 29104 19310 29132 20878
rect 29092 19304 29144 19310
rect 29092 19246 29144 19252
rect 28724 18760 28776 18766
rect 28722 18728 28724 18737
rect 29000 18760 29052 18766
rect 28776 18728 28778 18737
rect 28632 18692 28684 18698
rect 29000 18702 29052 18708
rect 28722 18663 28778 18672
rect 28632 18634 28684 18640
rect 28540 17876 28592 17882
rect 28540 17818 28592 17824
rect 28540 17672 28592 17678
rect 28540 17614 28592 17620
rect 28448 17604 28500 17610
rect 28448 17546 28500 17552
rect 28354 17368 28410 17377
rect 28354 17303 28410 17312
rect 28368 16998 28396 17303
rect 28356 16992 28408 16998
rect 28356 16934 28408 16940
rect 28264 16788 28316 16794
rect 28264 16730 28316 16736
rect 28172 16652 28224 16658
rect 28172 16594 28224 16600
rect 28080 16584 28132 16590
rect 28080 16526 28132 16532
rect 27988 16516 28040 16522
rect 27988 16458 28040 16464
rect 28000 16114 28028 16458
rect 28092 16250 28120 16526
rect 28080 16244 28132 16250
rect 28080 16186 28132 16192
rect 27988 16108 28040 16114
rect 27988 16050 28040 16056
rect 27896 15904 27948 15910
rect 27896 15846 27948 15852
rect 27988 15904 28040 15910
rect 27988 15846 28040 15852
rect 28080 15904 28132 15910
rect 28080 15846 28132 15852
rect 27804 14612 27856 14618
rect 27804 14554 27856 14560
rect 27802 14512 27858 14521
rect 27802 14447 27858 14456
rect 27712 14340 27764 14346
rect 27712 14282 27764 14288
rect 27724 14113 27752 14282
rect 27710 14104 27766 14113
rect 27710 14039 27766 14048
rect 27632 13926 27752 13954
rect 27620 13864 27672 13870
rect 27620 13806 27672 13812
rect 27528 13456 27580 13462
rect 27528 13398 27580 13404
rect 27528 12844 27580 12850
rect 27448 12804 27528 12832
rect 27252 12786 27304 12792
rect 27528 12786 27580 12792
rect 27160 10124 27212 10130
rect 27160 10066 27212 10072
rect 27080 9982 27200 10010
rect 27068 9648 27120 9654
rect 27068 9590 27120 9596
rect 27080 9518 27108 9590
rect 27068 9512 27120 9518
rect 27068 9454 27120 9460
rect 27068 8968 27120 8974
rect 27068 8910 27120 8916
rect 27080 8634 27108 8910
rect 27068 8628 27120 8634
rect 27068 8570 27120 8576
rect 27172 8480 27200 9982
rect 27264 9217 27292 12786
rect 27540 12714 27568 12786
rect 27528 12708 27580 12714
rect 27528 12650 27580 12656
rect 27632 11558 27660 13806
rect 27724 13190 27752 13926
rect 27816 13802 27844 14447
rect 27804 13796 27856 13802
rect 27804 13738 27856 13744
rect 27804 13252 27856 13258
rect 27804 13194 27856 13200
rect 27712 13184 27764 13190
rect 27712 13126 27764 13132
rect 27816 12968 27844 13194
rect 27724 12940 27844 12968
rect 27724 12850 27752 12940
rect 27908 12866 27936 15846
rect 28000 14657 28028 15846
rect 27986 14648 28042 14657
rect 27986 14583 28042 14592
rect 28092 14498 28120 15846
rect 28000 14470 28120 14498
rect 28000 13326 28028 14470
rect 28080 14408 28132 14414
rect 28078 14376 28080 14385
rect 28132 14376 28134 14385
rect 28078 14311 28134 14320
rect 28080 13932 28132 13938
rect 28080 13874 28132 13880
rect 28092 13734 28120 13874
rect 28080 13728 28132 13734
rect 28080 13670 28132 13676
rect 27988 13320 28040 13326
rect 27988 13262 28040 13268
rect 27712 12844 27764 12850
rect 27712 12786 27764 12792
rect 27816 12838 27936 12866
rect 28092 12850 28120 13670
rect 28080 12844 28132 12850
rect 27816 12646 27844 12838
rect 28080 12786 28132 12792
rect 27896 12776 27948 12782
rect 27896 12718 27948 12724
rect 27804 12640 27856 12646
rect 27804 12582 27856 12588
rect 27908 12628 27936 12718
rect 28080 12708 28132 12714
rect 28080 12650 28132 12656
rect 27988 12640 28040 12646
rect 27908 12600 27988 12628
rect 27908 12238 27936 12600
rect 27988 12582 28040 12588
rect 28092 12374 28120 12650
rect 28080 12368 28132 12374
rect 28080 12310 28132 12316
rect 27896 12232 27948 12238
rect 27896 12174 27948 12180
rect 27988 11756 28040 11762
rect 27988 11698 28040 11704
rect 27620 11552 27672 11558
rect 27620 11494 27672 11500
rect 27710 11520 27766 11529
rect 27710 11455 27766 11464
rect 27724 11150 27752 11455
rect 28000 11354 28028 11698
rect 28078 11384 28134 11393
rect 27988 11348 28040 11354
rect 28078 11319 28134 11328
rect 27988 11290 28040 11296
rect 27988 11212 28040 11218
rect 27988 11154 28040 11160
rect 27712 11144 27764 11150
rect 27712 11086 27764 11092
rect 27896 11144 27948 11150
rect 27896 11086 27948 11092
rect 27620 10668 27672 10674
rect 27620 10610 27672 10616
rect 27632 10577 27660 10610
rect 27618 10568 27674 10577
rect 27618 10503 27674 10512
rect 27724 10266 27752 11086
rect 27908 10810 27936 11086
rect 27804 10804 27856 10810
rect 27804 10746 27856 10752
rect 27896 10804 27948 10810
rect 27896 10746 27948 10752
rect 27712 10260 27764 10266
rect 27712 10202 27764 10208
rect 27816 10198 27844 10746
rect 28000 10674 28028 11154
rect 27988 10668 28040 10674
rect 27988 10610 28040 10616
rect 27804 10192 27856 10198
rect 27804 10134 27856 10140
rect 27620 10056 27672 10062
rect 27620 9998 27672 10004
rect 27344 9988 27396 9994
rect 27344 9930 27396 9936
rect 27356 9518 27384 9930
rect 27436 9580 27488 9586
rect 27436 9522 27488 9528
rect 27344 9512 27396 9518
rect 27344 9454 27396 9460
rect 27250 9208 27306 9217
rect 27250 9143 27306 9152
rect 27356 8974 27384 9454
rect 27344 8968 27396 8974
rect 27344 8910 27396 8916
rect 27172 8452 27292 8480
rect 27068 8424 27120 8430
rect 27264 8401 27292 8452
rect 27356 8430 27384 8910
rect 27448 8566 27476 9522
rect 27632 9382 27660 9998
rect 27896 9920 27948 9926
rect 27896 9862 27948 9868
rect 27908 9654 27936 9862
rect 27896 9648 27948 9654
rect 27896 9590 27948 9596
rect 27908 9518 27936 9590
rect 27896 9512 27948 9518
rect 27896 9454 27948 9460
rect 27620 9376 27672 9382
rect 27620 9318 27672 9324
rect 27804 9376 27856 9382
rect 27804 9318 27856 9324
rect 27632 9178 27660 9318
rect 27710 9208 27766 9217
rect 27620 9172 27672 9178
rect 27710 9143 27712 9152
rect 27620 9114 27672 9120
rect 27764 9143 27766 9152
rect 27712 9114 27764 9120
rect 27528 9036 27580 9042
rect 27528 8978 27580 8984
rect 27436 8560 27488 8566
rect 27436 8502 27488 8508
rect 27344 8424 27396 8430
rect 27068 8366 27120 8372
rect 27250 8392 27306 8401
rect 26976 8288 27028 8294
rect 26976 8230 27028 8236
rect 26792 8016 26844 8022
rect 26792 7958 26844 7964
rect 27080 7954 27108 8366
rect 27344 8366 27396 8372
rect 27250 8327 27306 8336
rect 26608 7948 26660 7954
rect 26608 7890 26660 7896
rect 27068 7948 27120 7954
rect 27068 7890 27120 7896
rect 27160 7948 27212 7954
rect 27160 7890 27212 7896
rect 26620 7410 26648 7890
rect 27080 7410 27108 7890
rect 27172 7857 27200 7890
rect 27158 7848 27214 7857
rect 27158 7783 27214 7792
rect 26516 7404 26568 7410
rect 26516 7346 26568 7352
rect 26608 7404 26660 7410
rect 26608 7346 26660 7352
rect 27068 7404 27120 7410
rect 27068 7346 27120 7352
rect 27080 7274 27108 7346
rect 27264 7342 27292 8327
rect 27448 8090 27476 8502
rect 27540 8498 27568 8978
rect 27724 8566 27752 9114
rect 27712 8560 27764 8566
rect 27712 8502 27764 8508
rect 27528 8492 27580 8498
rect 27528 8434 27580 8440
rect 27436 8084 27488 8090
rect 27436 8026 27488 8032
rect 27448 7410 27476 8026
rect 27540 8022 27568 8434
rect 27816 8294 27844 9318
rect 27804 8288 27856 8294
rect 27804 8230 27856 8236
rect 27528 8016 27580 8022
rect 27528 7958 27580 7964
rect 27436 7404 27488 7410
rect 27540 7392 27568 7958
rect 27816 7886 27844 8230
rect 27804 7880 27856 7886
rect 27804 7822 27856 7828
rect 27620 7404 27672 7410
rect 27540 7364 27620 7392
rect 27436 7346 27488 7352
rect 27620 7346 27672 7352
rect 27252 7336 27304 7342
rect 27252 7278 27304 7284
rect 27816 7274 27844 7822
rect 27068 7268 27120 7274
rect 27068 7210 27120 7216
rect 27804 7268 27856 7274
rect 27804 7210 27856 7216
rect 28000 7206 28028 10610
rect 28092 10538 28120 11319
rect 28080 10532 28132 10538
rect 28080 10474 28132 10480
rect 28080 10260 28132 10266
rect 28080 10202 28132 10208
rect 28092 7818 28120 10202
rect 28184 8022 28212 16594
rect 28448 16516 28500 16522
rect 28276 16476 28448 16504
rect 28276 16114 28304 16476
rect 28448 16458 28500 16464
rect 28264 16108 28316 16114
rect 28264 16050 28316 16056
rect 28356 16108 28408 16114
rect 28356 16050 28408 16056
rect 28368 15910 28396 16050
rect 28448 15972 28500 15978
rect 28448 15914 28500 15920
rect 28356 15904 28408 15910
rect 28356 15846 28408 15852
rect 28264 14408 28316 14414
rect 28264 14350 28316 14356
rect 28276 14074 28304 14350
rect 28264 14068 28316 14074
rect 28264 14010 28316 14016
rect 28460 14006 28488 15914
rect 28552 14770 28580 17614
rect 28644 16726 28672 18634
rect 28816 18624 28868 18630
rect 28816 18566 28868 18572
rect 28828 17882 28856 18566
rect 28816 17876 28868 17882
rect 28816 17818 28868 17824
rect 28998 17776 29054 17785
rect 28998 17711 29054 17720
rect 28724 17672 28776 17678
rect 28724 17614 28776 17620
rect 28816 17672 28868 17678
rect 28816 17614 28868 17620
rect 28736 17241 28764 17614
rect 28828 17338 28856 17614
rect 28816 17332 28868 17338
rect 28816 17274 28868 17280
rect 28722 17232 28778 17241
rect 28722 17167 28778 17176
rect 28906 17232 28962 17241
rect 29012 17218 29040 17711
rect 29092 17604 29144 17610
rect 29092 17546 29144 17552
rect 28962 17190 29040 17218
rect 28906 17167 28962 17176
rect 28724 17128 28776 17134
rect 28724 17070 28776 17076
rect 28632 16720 28684 16726
rect 28632 16662 28684 16668
rect 28632 16584 28684 16590
rect 28630 16552 28632 16561
rect 28684 16552 28686 16561
rect 28630 16487 28686 16496
rect 28736 15706 28764 17070
rect 29000 17060 29052 17066
rect 29000 17002 29052 17008
rect 28814 16688 28870 16697
rect 28814 16623 28870 16632
rect 28724 15700 28776 15706
rect 28724 15642 28776 15648
rect 28552 14742 28672 14770
rect 28538 14648 28594 14657
rect 28538 14583 28540 14592
rect 28592 14583 28594 14592
rect 28540 14554 28592 14560
rect 28644 14464 28672 14742
rect 28644 14436 28708 14464
rect 28540 14340 28592 14346
rect 28680 14328 28708 14436
rect 28540 14282 28592 14288
rect 28644 14300 28708 14328
rect 28552 14006 28580 14282
rect 28448 14000 28500 14006
rect 28448 13942 28500 13948
rect 28540 14000 28592 14006
rect 28540 13942 28592 13948
rect 28264 13456 28316 13462
rect 28264 13398 28316 13404
rect 28276 12850 28304 13398
rect 28356 13184 28408 13190
rect 28356 13126 28408 13132
rect 28368 12850 28396 13126
rect 28264 12844 28316 12850
rect 28264 12786 28316 12792
rect 28356 12844 28408 12850
rect 28356 12786 28408 12792
rect 28264 12708 28316 12714
rect 28264 12650 28316 12656
rect 28356 12708 28408 12714
rect 28356 12650 28408 12656
rect 28276 11354 28304 12650
rect 28368 11937 28396 12650
rect 28354 11928 28410 11937
rect 28354 11863 28410 11872
rect 28460 11762 28488 13942
rect 28540 12232 28592 12238
rect 28540 12174 28592 12180
rect 28448 11756 28500 11762
rect 28448 11698 28500 11704
rect 28356 11552 28408 11558
rect 28356 11494 28408 11500
rect 28264 11348 28316 11354
rect 28264 11290 28316 11296
rect 28368 11150 28396 11494
rect 28356 11144 28408 11150
rect 28356 11086 28408 11092
rect 28368 10810 28396 11086
rect 28552 11014 28580 12174
rect 28644 11558 28672 14300
rect 28724 14000 28776 14006
rect 28724 13942 28776 13948
rect 28736 12850 28764 13942
rect 28828 13938 28856 16623
rect 28908 15904 28960 15910
rect 28908 15846 28960 15852
rect 28920 15502 28948 15846
rect 28908 15496 28960 15502
rect 28908 15438 28960 15444
rect 28908 15360 28960 15366
rect 28908 15302 28960 15308
rect 28920 14550 28948 15302
rect 29012 15026 29040 17002
rect 29104 16794 29132 17546
rect 29092 16788 29144 16794
rect 29092 16730 29144 16736
rect 29092 15496 29144 15502
rect 29092 15438 29144 15444
rect 29104 15337 29132 15438
rect 29090 15328 29146 15337
rect 29090 15263 29146 15272
rect 29000 15020 29052 15026
rect 29000 14962 29052 14968
rect 29012 14618 29040 14962
rect 29000 14612 29052 14618
rect 29000 14554 29052 14560
rect 28908 14544 28960 14550
rect 28906 14512 28908 14521
rect 28960 14512 28962 14521
rect 28906 14447 28962 14456
rect 29012 14414 29040 14554
rect 28908 14408 28960 14414
rect 28906 14376 28908 14385
rect 29000 14408 29052 14414
rect 28960 14376 28962 14385
rect 29000 14350 29052 14356
rect 28906 14311 28962 14320
rect 28906 14104 28962 14113
rect 28906 14039 28962 14048
rect 28816 13932 28868 13938
rect 28816 13874 28868 13880
rect 28920 12986 28948 14039
rect 29012 13802 29040 14350
rect 29000 13796 29052 13802
rect 29000 13738 29052 13744
rect 29196 13734 29224 23734
rect 29276 23588 29328 23594
rect 29276 23530 29328 23536
rect 29288 23322 29316 23530
rect 29276 23316 29328 23322
rect 29276 23258 29328 23264
rect 29276 23044 29328 23050
rect 29276 22986 29328 22992
rect 29288 22545 29316 22986
rect 29460 22636 29512 22642
rect 29460 22578 29512 22584
rect 29274 22536 29330 22545
rect 29274 22471 29330 22480
rect 29472 20369 29500 22578
rect 29458 20360 29514 20369
rect 29458 20295 29514 20304
rect 29368 19372 29420 19378
rect 29368 19314 29420 19320
rect 29460 19372 29512 19378
rect 29460 19314 29512 19320
rect 29276 19236 29328 19242
rect 29276 19178 29328 19184
rect 29288 18902 29316 19178
rect 29276 18896 29328 18902
rect 29276 18838 29328 18844
rect 29288 18630 29316 18838
rect 29380 18766 29408 19314
rect 29368 18760 29420 18766
rect 29368 18702 29420 18708
rect 29276 18624 29328 18630
rect 29276 18566 29328 18572
rect 29380 18154 29408 18702
rect 29368 18148 29420 18154
rect 29368 18090 29420 18096
rect 29276 17672 29328 17678
rect 29276 17614 29328 17620
rect 29288 16998 29316 17614
rect 29276 16992 29328 16998
rect 29276 16934 29328 16940
rect 29288 16046 29316 16934
rect 29276 16040 29328 16046
rect 29276 15982 29328 15988
rect 29276 15360 29328 15366
rect 29276 15302 29328 15308
rect 29184 13728 29236 13734
rect 29090 13696 29146 13705
rect 29184 13670 29236 13676
rect 29090 13631 29146 13640
rect 29104 12986 29132 13631
rect 29288 13258 29316 15302
rect 29276 13252 29328 13258
rect 29276 13194 29328 13200
rect 29184 13184 29236 13190
rect 29184 13126 29236 13132
rect 28908 12980 28960 12986
rect 28908 12922 28960 12928
rect 29092 12980 29144 12986
rect 29092 12922 29144 12928
rect 29196 12850 29224 13126
rect 29288 12918 29316 13194
rect 29276 12912 29328 12918
rect 29276 12854 29328 12860
rect 28724 12844 28776 12850
rect 28724 12786 28776 12792
rect 28816 12844 28868 12850
rect 28816 12786 28868 12792
rect 29184 12844 29236 12850
rect 29184 12786 29236 12792
rect 28736 12102 28764 12786
rect 28828 12646 28856 12786
rect 28816 12640 28868 12646
rect 28816 12582 28868 12588
rect 29092 12640 29144 12646
rect 29092 12582 29144 12588
rect 28724 12096 28776 12102
rect 28724 12038 28776 12044
rect 28632 11552 28684 11558
rect 28632 11494 28684 11500
rect 28828 11150 28856 12582
rect 28816 11144 28868 11150
rect 28816 11086 28868 11092
rect 28540 11008 28592 11014
rect 28540 10950 28592 10956
rect 28356 10804 28408 10810
rect 28356 10746 28408 10752
rect 28540 10736 28592 10742
rect 28540 10678 28592 10684
rect 28264 10668 28316 10674
rect 28264 10610 28316 10616
rect 28276 9926 28304 10610
rect 28448 10056 28500 10062
rect 28448 9998 28500 10004
rect 28264 9920 28316 9926
rect 28264 9862 28316 9868
rect 28460 9586 28488 9998
rect 28448 9580 28500 9586
rect 28448 9522 28500 9528
rect 28262 9480 28318 9489
rect 28262 9415 28318 9424
rect 28276 8974 28304 9415
rect 28356 9172 28408 9178
rect 28356 9114 28408 9120
rect 28264 8968 28316 8974
rect 28264 8910 28316 8916
rect 28264 8356 28316 8362
rect 28368 8344 28396 9114
rect 28460 8362 28488 9522
rect 28552 9110 28580 10678
rect 28828 10674 28856 11086
rect 29104 11014 29132 12582
rect 29184 11144 29236 11150
rect 29184 11086 29236 11092
rect 29092 11008 29144 11014
rect 29092 10950 29144 10956
rect 29196 10674 29224 11086
rect 28816 10668 28868 10674
rect 28816 10610 28868 10616
rect 29184 10668 29236 10674
rect 29184 10610 29236 10616
rect 28906 10568 28962 10577
rect 28906 10503 28962 10512
rect 28632 10056 28684 10062
rect 28920 10044 28948 10503
rect 29184 10260 29236 10266
rect 29184 10202 29236 10208
rect 29092 10056 29144 10062
rect 28920 10016 29092 10044
rect 28632 9998 28684 10004
rect 29092 9998 29144 10004
rect 28644 9722 28672 9998
rect 28632 9716 28684 9722
rect 28632 9658 28684 9664
rect 28644 9382 28672 9658
rect 29092 9648 29144 9654
rect 29090 9616 29092 9625
rect 29144 9616 29146 9625
rect 29090 9551 29146 9560
rect 28906 9480 28962 9489
rect 28906 9415 28962 9424
rect 28632 9376 28684 9382
rect 28632 9318 28684 9324
rect 28920 9110 28948 9415
rect 29000 9376 29052 9382
rect 29000 9318 29052 9324
rect 28540 9104 28592 9110
rect 28540 9046 28592 9052
rect 28908 9104 28960 9110
rect 28908 9046 28960 9052
rect 28552 8838 28580 9046
rect 28724 8968 28776 8974
rect 28724 8910 28776 8916
rect 28632 8900 28684 8906
rect 28632 8842 28684 8848
rect 28540 8832 28592 8838
rect 28540 8774 28592 8780
rect 28644 8634 28672 8842
rect 28736 8634 28764 8910
rect 28908 8832 28960 8838
rect 28908 8774 28960 8780
rect 28814 8664 28870 8673
rect 28632 8628 28684 8634
rect 28632 8570 28684 8576
rect 28724 8628 28776 8634
rect 28814 8599 28816 8608
rect 28724 8570 28776 8576
rect 28868 8599 28870 8608
rect 28816 8570 28868 8576
rect 28920 8498 28948 8774
rect 29012 8566 29040 9318
rect 29104 8906 29132 9551
rect 29196 9042 29224 10202
rect 29184 9036 29236 9042
rect 29184 8978 29236 8984
rect 29092 8900 29144 8906
rect 29092 8842 29144 8848
rect 29000 8560 29052 8566
rect 29000 8502 29052 8508
rect 28908 8492 28960 8498
rect 28908 8434 28960 8440
rect 29092 8492 29144 8498
rect 29196 8480 29224 8978
rect 29144 8452 29224 8480
rect 29092 8434 29144 8440
rect 28998 8392 29054 8401
rect 28316 8316 28396 8344
rect 28448 8356 28500 8362
rect 28264 8298 28316 8304
rect 28998 8327 29000 8336
rect 28448 8298 28500 8304
rect 29052 8327 29054 8336
rect 29000 8298 29052 8304
rect 28276 8090 28304 8298
rect 28632 8288 28684 8294
rect 28632 8230 28684 8236
rect 28644 8090 28672 8230
rect 28264 8084 28316 8090
rect 28264 8026 28316 8032
rect 28632 8084 28684 8090
rect 28632 8026 28684 8032
rect 28172 8016 28224 8022
rect 28172 7958 28224 7964
rect 29012 7954 29040 8298
rect 29000 7948 29052 7954
rect 29000 7890 29052 7896
rect 28816 7880 28868 7886
rect 28816 7822 28868 7828
rect 29184 7880 29236 7886
rect 29184 7822 29236 7828
rect 28080 7812 28132 7818
rect 28080 7754 28132 7760
rect 27988 7200 28040 7206
rect 27988 7142 28040 7148
rect 25964 6860 26016 6866
rect 25964 6802 26016 6808
rect 25596 6180 25648 6186
rect 25596 6122 25648 6128
rect 25504 5908 25556 5914
rect 25504 5850 25556 5856
rect 25412 5840 25464 5846
rect 25412 5782 25464 5788
rect 25136 5704 25188 5710
rect 25136 5646 25188 5652
rect 25424 5642 25452 5782
rect 25516 5642 25544 5850
rect 25688 5704 25740 5710
rect 25688 5646 25740 5652
rect 25780 5704 25832 5710
rect 25780 5646 25832 5652
rect 25412 5636 25464 5642
rect 25412 5578 25464 5584
rect 25504 5636 25556 5642
rect 25504 5578 25556 5584
rect 25700 5574 25728 5646
rect 24952 5568 25004 5574
rect 24952 5510 25004 5516
rect 25044 5568 25096 5574
rect 25044 5510 25096 5516
rect 25136 5568 25188 5574
rect 25136 5510 25188 5516
rect 25688 5568 25740 5574
rect 25688 5510 25740 5516
rect 25056 5302 25084 5510
rect 24860 5296 24912 5302
rect 24860 5238 24912 5244
rect 25044 5296 25096 5302
rect 25044 5238 25096 5244
rect 24872 4706 24900 5238
rect 24780 4690 24900 4706
rect 24768 4684 24900 4690
rect 24820 4678 24900 4684
rect 24768 4626 24820 4632
rect 24596 4542 24808 4570
rect 24780 4486 24808 4542
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 23940 4208 23992 4214
rect 23940 4150 23992 4156
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23388 4072 23440 4078
rect 23388 4014 23440 4020
rect 23296 3732 23348 3738
rect 23296 3674 23348 3680
rect 23112 3596 23164 3602
rect 23112 3538 23164 3544
rect 23032 3454 23152 3482
rect 23124 3058 23152 3454
rect 23112 3052 23164 3058
rect 23112 2994 23164 3000
rect 23124 2774 23152 2994
rect 23400 2990 23428 4014
rect 23492 3126 23520 4082
rect 23952 3126 23980 4150
rect 24780 3534 24808 4422
rect 24872 3602 24900 4678
rect 25148 4554 25176 5510
rect 25700 5166 25728 5510
rect 25792 5370 25820 5646
rect 25976 5574 26004 6802
rect 28092 6662 28120 7754
rect 28264 7744 28316 7750
rect 28264 7686 28316 7692
rect 28276 7274 28304 7686
rect 28264 7268 28316 7274
rect 28264 7210 28316 7216
rect 28276 6934 28304 7210
rect 28828 7206 28856 7822
rect 29196 7449 29224 7822
rect 29182 7440 29238 7449
rect 29182 7375 29184 7384
rect 29236 7375 29238 7384
rect 29184 7346 29236 7352
rect 28816 7200 28868 7206
rect 28816 7142 28868 7148
rect 28264 6928 28316 6934
rect 28264 6870 28316 6876
rect 29000 6860 29052 6866
rect 29000 6802 29052 6808
rect 28080 6656 28132 6662
rect 28080 6598 28132 6604
rect 26516 6452 26568 6458
rect 26516 6394 26568 6400
rect 26884 6452 26936 6458
rect 26884 6394 26936 6400
rect 26240 6384 26292 6390
rect 26240 6326 26292 6332
rect 26252 6254 26280 6326
rect 26240 6248 26292 6254
rect 26240 6190 26292 6196
rect 26252 5710 26280 6190
rect 26424 5908 26476 5914
rect 26424 5850 26476 5856
rect 26240 5704 26292 5710
rect 26240 5646 26292 5652
rect 26436 5642 26464 5850
rect 26528 5642 26556 6394
rect 26896 6322 26924 6394
rect 26792 6316 26844 6322
rect 26792 6258 26844 6264
rect 26884 6316 26936 6322
rect 26884 6258 26936 6264
rect 27344 6316 27396 6322
rect 27344 6258 27396 6264
rect 28724 6316 28776 6322
rect 28724 6258 28776 6264
rect 26700 5840 26752 5846
rect 26700 5782 26752 5788
rect 26424 5636 26476 5642
rect 26424 5578 26476 5584
rect 26516 5636 26568 5642
rect 26516 5578 26568 5584
rect 25964 5568 26016 5574
rect 25964 5510 26016 5516
rect 25780 5364 25832 5370
rect 25780 5306 25832 5312
rect 25688 5160 25740 5166
rect 25688 5102 25740 5108
rect 26148 5160 26200 5166
rect 26148 5102 26200 5108
rect 26160 4622 26188 5102
rect 26712 4622 26740 5782
rect 26804 5370 26832 6258
rect 26896 5710 26924 6258
rect 27356 6118 27384 6258
rect 27252 6112 27304 6118
rect 27252 6054 27304 6060
rect 27344 6112 27396 6118
rect 27344 6054 27396 6060
rect 27264 5778 27292 6054
rect 27252 5772 27304 5778
rect 27252 5714 27304 5720
rect 26884 5704 26936 5710
rect 26884 5646 26936 5652
rect 27356 5642 27384 6054
rect 28736 5953 28764 6258
rect 28722 5944 28778 5953
rect 28722 5879 28724 5888
rect 28776 5879 28778 5888
rect 28724 5850 28776 5856
rect 27344 5636 27396 5642
rect 27344 5578 27396 5584
rect 28080 5568 28132 5574
rect 28080 5510 28132 5516
rect 26792 5364 26844 5370
rect 26792 5306 26844 5312
rect 28092 5166 28120 5510
rect 28172 5296 28224 5302
rect 28172 5238 28224 5244
rect 28080 5160 28132 5166
rect 28080 5102 28132 5108
rect 26148 4616 26200 4622
rect 26148 4558 26200 4564
rect 26700 4616 26752 4622
rect 26700 4558 26752 4564
rect 25136 4548 25188 4554
rect 25136 4490 25188 4496
rect 28184 4146 28212 5238
rect 29012 5234 29040 6802
rect 29288 6798 29316 12854
rect 29472 12442 29500 19314
rect 29564 17785 29592 25842
rect 29644 24336 29696 24342
rect 29644 24278 29696 24284
rect 29656 23798 29684 24278
rect 29644 23792 29696 23798
rect 29644 23734 29696 23740
rect 29642 23080 29698 23089
rect 29642 23015 29698 23024
rect 29656 22778 29684 23015
rect 29644 22772 29696 22778
rect 29644 22714 29696 22720
rect 29644 22092 29696 22098
rect 29644 22034 29696 22040
rect 29656 21078 29684 22034
rect 29748 21350 29776 26250
rect 29828 23112 29880 23118
rect 29828 23054 29880 23060
rect 29840 22137 29868 23054
rect 29920 22636 29972 22642
rect 29920 22578 29972 22584
rect 29932 22409 29960 22578
rect 30024 22545 30052 26862
rect 30010 22536 30066 22545
rect 30010 22471 30066 22480
rect 30012 22432 30064 22438
rect 29918 22400 29974 22409
rect 30012 22374 30064 22380
rect 29918 22335 29974 22344
rect 30024 22234 30052 22374
rect 30012 22228 30064 22234
rect 30012 22170 30064 22176
rect 29826 22128 29882 22137
rect 29826 22063 29882 22072
rect 29736 21344 29788 21350
rect 29736 21286 29788 21292
rect 29644 21072 29696 21078
rect 29644 21014 29696 21020
rect 29840 20777 29868 22063
rect 30012 21888 30064 21894
rect 29932 21848 30012 21876
rect 29932 20942 29960 21848
rect 30012 21830 30064 21836
rect 29920 20936 29972 20942
rect 29920 20878 29972 20884
rect 30012 20936 30064 20942
rect 30012 20878 30064 20884
rect 29826 20768 29882 20777
rect 29826 20703 29882 20712
rect 29736 20528 29788 20534
rect 29734 20496 29736 20505
rect 29788 20496 29790 20505
rect 29734 20431 29790 20440
rect 29828 20460 29880 20466
rect 29644 19236 29696 19242
rect 29644 19178 29696 19184
rect 29550 17776 29606 17785
rect 29550 17711 29606 17720
rect 29552 16244 29604 16250
rect 29552 16186 29604 16192
rect 29564 15314 29592 16186
rect 29656 15434 29684 19178
rect 29644 15428 29696 15434
rect 29644 15370 29696 15376
rect 29564 15286 29684 15314
rect 29656 14550 29684 15286
rect 29644 14544 29696 14550
rect 29644 14486 29696 14492
rect 29552 13932 29604 13938
rect 29552 13874 29604 13880
rect 29460 12436 29512 12442
rect 29460 12378 29512 12384
rect 29564 12322 29592 13874
rect 29380 12294 29592 12322
rect 29380 7546 29408 12294
rect 29460 12096 29512 12102
rect 29460 12038 29512 12044
rect 29472 11762 29500 12038
rect 29460 11756 29512 11762
rect 29460 11698 29512 11704
rect 29472 11150 29500 11698
rect 29552 11688 29604 11694
rect 29552 11630 29604 11636
rect 29564 11354 29592 11630
rect 29552 11348 29604 11354
rect 29552 11290 29604 11296
rect 29550 11248 29606 11257
rect 29550 11183 29606 11192
rect 29460 11144 29512 11150
rect 29460 11086 29512 11092
rect 29460 11008 29512 11014
rect 29458 10976 29460 10985
rect 29512 10976 29514 10985
rect 29458 10911 29514 10920
rect 29564 10248 29592 11183
rect 29656 10742 29684 14486
rect 29748 12986 29776 20431
rect 29828 20402 29880 20408
rect 29840 20262 29868 20402
rect 29828 20256 29880 20262
rect 29828 20198 29880 20204
rect 29932 20074 29960 20878
rect 30024 20466 30052 20878
rect 30012 20460 30064 20466
rect 30012 20402 30064 20408
rect 29840 20046 29960 20074
rect 29840 15502 29868 20046
rect 29920 19984 29972 19990
rect 29920 19926 29972 19932
rect 29932 19378 29960 19926
rect 30024 19378 30052 20402
rect 30116 19990 30144 27814
rect 30392 27674 30420 28358
rect 30380 27668 30432 27674
rect 30380 27610 30432 27616
rect 30288 24744 30340 24750
rect 30288 24686 30340 24692
rect 30196 23248 30248 23254
rect 30196 23190 30248 23196
rect 30208 22778 30236 23190
rect 30196 22772 30248 22778
rect 30196 22714 30248 22720
rect 30208 22030 30236 22714
rect 30300 22624 30328 24686
rect 30392 23730 30420 27610
rect 30484 27033 30512 29464
rect 30576 28014 30604 30194
rect 30748 29504 30800 29510
rect 30748 29446 30800 29452
rect 30760 29306 30788 29446
rect 30748 29300 30800 29306
rect 30748 29242 30800 29248
rect 30656 28484 30708 28490
rect 30656 28426 30708 28432
rect 30564 28008 30616 28014
rect 30564 27950 30616 27956
rect 30576 27538 30604 27950
rect 30668 27878 30696 28426
rect 30852 28150 30880 31282
rect 30944 29578 30972 32671
rect 31036 31822 31064 33254
rect 31128 32502 31156 34682
rect 31220 33017 31248 41006
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 35594 40284 35902 40293
rect 35594 40282 35600 40284
rect 35656 40282 35680 40284
rect 35736 40282 35760 40284
rect 35816 40282 35840 40284
rect 35896 40282 35902 40284
rect 35656 40230 35658 40282
rect 35838 40230 35840 40282
rect 35594 40228 35600 40230
rect 35656 40228 35680 40230
rect 35736 40228 35760 40230
rect 35816 40228 35840 40230
rect 35896 40228 35902 40230
rect 35594 40219 35902 40228
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 35594 39196 35902 39205
rect 35594 39194 35600 39196
rect 35656 39194 35680 39196
rect 35736 39194 35760 39196
rect 35816 39194 35840 39196
rect 35896 39194 35902 39196
rect 35656 39142 35658 39194
rect 35838 39142 35840 39194
rect 35594 39140 35600 39142
rect 35656 39140 35680 39142
rect 35736 39140 35760 39142
rect 35816 39140 35840 39142
rect 35896 39140 35902 39142
rect 35594 39131 35902 39140
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 35594 38108 35902 38117
rect 35594 38106 35600 38108
rect 35656 38106 35680 38108
rect 35736 38106 35760 38108
rect 35816 38106 35840 38108
rect 35896 38106 35902 38108
rect 35656 38054 35658 38106
rect 35838 38054 35840 38106
rect 35594 38052 35600 38054
rect 35656 38052 35680 38054
rect 35736 38052 35760 38054
rect 35816 38052 35840 38054
rect 35896 38052 35902 38054
rect 35594 38043 35902 38052
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35594 37020 35902 37029
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 32036 33992 32088 33998
rect 32036 33934 32088 33940
rect 31392 33856 31444 33862
rect 31392 33798 31444 33804
rect 31404 33522 31432 33798
rect 31392 33516 31444 33522
rect 31392 33458 31444 33464
rect 31944 33516 31996 33522
rect 31944 33458 31996 33464
rect 31206 33008 31262 33017
rect 31206 32943 31262 32952
rect 31116 32496 31168 32502
rect 31116 32438 31168 32444
rect 31404 32434 31432 33458
rect 31668 32768 31720 32774
rect 31668 32710 31720 32716
rect 31392 32428 31444 32434
rect 31392 32370 31444 32376
rect 31484 32428 31536 32434
rect 31484 32370 31536 32376
rect 31404 31958 31432 32370
rect 31392 31952 31444 31958
rect 31392 31894 31444 31900
rect 31024 31816 31076 31822
rect 31024 31758 31076 31764
rect 31392 31816 31444 31822
rect 31392 31758 31444 31764
rect 31036 30161 31064 31758
rect 31208 30728 31260 30734
rect 31260 30676 31340 30682
rect 31208 30670 31340 30676
rect 31220 30654 31340 30670
rect 31116 30592 31168 30598
rect 31116 30534 31168 30540
rect 31128 30258 31156 30534
rect 31312 30258 31340 30654
rect 31116 30252 31168 30258
rect 31116 30194 31168 30200
rect 31300 30252 31352 30258
rect 31300 30194 31352 30200
rect 31022 30152 31078 30161
rect 31022 30087 31078 30096
rect 31022 30016 31078 30025
rect 31022 29951 31078 29960
rect 31036 29782 31064 29951
rect 31024 29776 31076 29782
rect 31024 29718 31076 29724
rect 30932 29572 30984 29578
rect 30932 29514 30984 29520
rect 30840 28144 30892 28150
rect 30840 28086 30892 28092
rect 30748 28076 30800 28082
rect 30748 28018 30800 28024
rect 30656 27872 30708 27878
rect 30656 27814 30708 27820
rect 30760 27606 30788 28018
rect 30748 27600 30800 27606
rect 30748 27542 30800 27548
rect 30564 27532 30616 27538
rect 30564 27474 30616 27480
rect 30470 27024 30526 27033
rect 30470 26959 30526 26968
rect 30746 27024 30802 27033
rect 30746 26959 30748 26968
rect 30800 26959 30802 26968
rect 30748 26930 30800 26936
rect 30748 26376 30800 26382
rect 30748 26318 30800 26324
rect 30760 25702 30788 26318
rect 30852 26042 30880 28086
rect 31208 27668 31260 27674
rect 31208 27610 31260 27616
rect 30932 27600 30984 27606
rect 30932 27542 30984 27548
rect 30944 26353 30972 27542
rect 31024 27532 31076 27538
rect 31024 27474 31076 27480
rect 31036 27130 31064 27474
rect 31114 27432 31170 27441
rect 31220 27402 31248 27610
rect 31114 27367 31170 27376
rect 31208 27396 31260 27402
rect 31128 27130 31156 27367
rect 31208 27338 31260 27344
rect 31024 27124 31076 27130
rect 31024 27066 31076 27072
rect 31116 27124 31168 27130
rect 31116 27066 31168 27072
rect 31022 26888 31078 26897
rect 31022 26823 31078 26832
rect 30930 26344 30986 26353
rect 30930 26279 30986 26288
rect 30840 26036 30892 26042
rect 30840 25978 30892 25984
rect 30932 25900 30984 25906
rect 31036 25888 31064 26823
rect 31128 26246 31156 27066
rect 31208 26308 31260 26314
rect 31208 26250 31260 26256
rect 31116 26240 31168 26246
rect 31116 26182 31168 26188
rect 31128 25974 31156 26182
rect 31116 25968 31168 25974
rect 31116 25910 31168 25916
rect 30984 25860 31064 25888
rect 30932 25842 30984 25848
rect 30748 25696 30800 25702
rect 30748 25638 30800 25644
rect 30656 25492 30708 25498
rect 30656 25434 30708 25440
rect 30668 24818 30696 25434
rect 30760 25294 30788 25638
rect 30944 25362 30972 25842
rect 30932 25356 30984 25362
rect 30932 25298 30984 25304
rect 30748 25288 30800 25294
rect 30748 25230 30800 25236
rect 30656 24812 30708 24818
rect 30656 24754 30708 24760
rect 30840 24812 30892 24818
rect 30840 24754 30892 24760
rect 30380 23724 30432 23730
rect 30380 23666 30432 23672
rect 30380 22636 30432 22642
rect 30300 22596 30380 22624
rect 30432 22596 30512 22624
rect 30380 22578 30432 22584
rect 30288 22500 30340 22506
rect 30288 22442 30340 22448
rect 30196 22024 30248 22030
rect 30196 21966 30248 21972
rect 30196 21344 30248 21350
rect 30196 21286 30248 21292
rect 30104 19984 30156 19990
rect 30104 19926 30156 19932
rect 30102 19816 30158 19825
rect 30102 19751 30158 19760
rect 29920 19372 29972 19378
rect 29920 19314 29972 19320
rect 30012 19372 30064 19378
rect 30012 19314 30064 19320
rect 29932 19174 29960 19314
rect 29920 19168 29972 19174
rect 29920 19110 29972 19116
rect 29920 18760 29972 18766
rect 29918 18728 29920 18737
rect 29972 18728 29974 18737
rect 29918 18663 29974 18672
rect 29920 18624 29972 18630
rect 29920 18566 29972 18572
rect 29932 15570 29960 18566
rect 30024 18222 30052 19314
rect 30116 19310 30144 19751
rect 30208 19394 30236 21286
rect 30300 20874 30328 22442
rect 30484 22098 30512 22596
rect 30564 22568 30616 22574
rect 30564 22510 30616 22516
rect 30472 22092 30524 22098
rect 30472 22034 30524 22040
rect 30576 22030 30604 22510
rect 30564 22024 30616 22030
rect 30564 21966 30616 21972
rect 30472 20936 30524 20942
rect 30470 20904 30472 20913
rect 30524 20904 30526 20913
rect 30288 20868 30340 20874
rect 30470 20839 30526 20848
rect 30288 20810 30340 20816
rect 30300 19514 30328 20810
rect 30472 20800 30524 20806
rect 30472 20742 30524 20748
rect 30484 20602 30512 20742
rect 30472 20596 30524 20602
rect 30472 20538 30524 20544
rect 30484 19786 30512 20538
rect 30668 20262 30696 24754
rect 30852 20534 30880 24754
rect 30944 24410 30972 25298
rect 31024 25152 31076 25158
rect 31024 25094 31076 25100
rect 30932 24404 30984 24410
rect 30932 24346 30984 24352
rect 30932 23724 30984 23730
rect 30932 23666 30984 23672
rect 30944 21350 30972 23666
rect 31036 23594 31064 25094
rect 31116 24064 31168 24070
rect 31116 24006 31168 24012
rect 31128 23866 31156 24006
rect 31116 23860 31168 23866
rect 31116 23802 31168 23808
rect 31024 23588 31076 23594
rect 31024 23530 31076 23536
rect 31220 23118 31248 26250
rect 31312 25974 31340 30194
rect 31404 30122 31432 31758
rect 31496 31686 31524 32370
rect 31680 32298 31708 32710
rect 31956 32570 31984 33458
rect 32048 32978 32076 33934
rect 32680 33924 32732 33930
rect 32680 33866 32732 33872
rect 32496 33856 32548 33862
rect 32496 33798 32548 33804
rect 32036 32972 32088 32978
rect 32036 32914 32088 32920
rect 32220 32904 32272 32910
rect 32220 32846 32272 32852
rect 31944 32564 31996 32570
rect 31944 32506 31996 32512
rect 31668 32292 31720 32298
rect 31668 32234 31720 32240
rect 31680 32026 31708 32234
rect 31852 32224 31904 32230
rect 31852 32166 31904 32172
rect 31668 32020 31720 32026
rect 31668 31962 31720 31968
rect 31576 31884 31628 31890
rect 31864 31872 31892 32166
rect 32126 32056 32182 32065
rect 32232 32026 32260 32846
rect 32508 32842 32536 33798
rect 32692 33658 32720 33866
rect 34060 33856 34112 33862
rect 34060 33798 34112 33804
rect 32680 33652 32732 33658
rect 32680 33594 32732 33600
rect 34072 33522 34100 33798
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 32956 33516 33008 33522
rect 32956 33458 33008 33464
rect 34060 33516 34112 33522
rect 34060 33458 34112 33464
rect 34244 33516 34296 33522
rect 34244 33458 34296 33464
rect 32496 32836 32548 32842
rect 32496 32778 32548 32784
rect 32404 32768 32456 32774
rect 32324 32728 32404 32756
rect 32126 31991 32128 32000
rect 32180 31991 32182 32000
rect 32220 32020 32272 32026
rect 32128 31962 32180 31968
rect 32220 31962 32272 31968
rect 31628 31844 31892 31872
rect 31576 31826 31628 31832
rect 32220 31816 32272 31822
rect 32220 31758 32272 31764
rect 31576 31748 31628 31754
rect 31576 31690 31628 31696
rect 32036 31748 32088 31754
rect 32036 31690 32088 31696
rect 31484 31680 31536 31686
rect 31484 31622 31536 31628
rect 31392 30116 31444 30122
rect 31392 30058 31444 30064
rect 31390 30016 31446 30025
rect 31390 29951 31446 29960
rect 31404 28150 31432 29951
rect 31496 29306 31524 31622
rect 31588 31278 31616 31690
rect 31576 31272 31628 31278
rect 31576 31214 31628 31220
rect 31576 31136 31628 31142
rect 31576 31078 31628 31084
rect 31588 30734 31616 31078
rect 32048 30734 32076 31690
rect 32128 30796 32180 30802
rect 32128 30738 32180 30744
rect 31576 30728 31628 30734
rect 31576 30670 31628 30676
rect 32036 30728 32088 30734
rect 32036 30670 32088 30676
rect 31668 30660 31720 30666
rect 31668 30602 31720 30608
rect 31574 30424 31630 30433
rect 31574 30359 31630 30368
rect 31588 30054 31616 30359
rect 31680 30054 31708 30602
rect 31760 30320 31812 30326
rect 31758 30288 31760 30297
rect 31944 30320 31996 30326
rect 31812 30288 31814 30297
rect 31944 30262 31996 30268
rect 31758 30223 31814 30232
rect 31760 30184 31812 30190
rect 31760 30126 31812 30132
rect 31576 30048 31628 30054
rect 31576 29990 31628 29996
rect 31668 30048 31720 30054
rect 31668 29990 31720 29996
rect 31772 29714 31800 30126
rect 31760 29708 31812 29714
rect 31760 29650 31812 29656
rect 31852 29708 31904 29714
rect 31852 29650 31904 29656
rect 31484 29300 31536 29306
rect 31484 29242 31536 29248
rect 31772 29238 31800 29650
rect 31864 29510 31892 29650
rect 31956 29510 31984 30262
rect 32048 30122 32076 30670
rect 32140 30258 32168 30738
rect 32128 30252 32180 30258
rect 32128 30194 32180 30200
rect 32036 30116 32088 30122
rect 32036 30058 32088 30064
rect 32232 30025 32260 31758
rect 32324 30666 32352 32728
rect 32508 32745 32536 32778
rect 32404 32710 32456 32716
rect 32494 32736 32550 32745
rect 32494 32671 32550 32680
rect 32404 32428 32456 32434
rect 32404 32370 32456 32376
rect 32416 32026 32444 32370
rect 32404 32020 32456 32026
rect 32404 31962 32456 31968
rect 32968 31958 32996 33458
rect 33140 33312 33192 33318
rect 33140 33254 33192 33260
rect 33048 32496 33100 32502
rect 33048 32438 33100 32444
rect 32496 31952 32548 31958
rect 32496 31894 32548 31900
rect 32956 31952 33008 31958
rect 32956 31894 33008 31900
rect 32312 30660 32364 30666
rect 32312 30602 32364 30608
rect 32312 30252 32364 30258
rect 32312 30194 32364 30200
rect 32218 30016 32274 30025
rect 32218 29951 32274 29960
rect 31852 29504 31904 29510
rect 31852 29446 31904 29452
rect 31944 29504 31996 29510
rect 31944 29446 31996 29452
rect 31760 29232 31812 29238
rect 31760 29174 31812 29180
rect 31392 28144 31444 28150
rect 31392 28086 31444 28092
rect 31404 27402 31432 28086
rect 31668 28008 31720 28014
rect 31668 27950 31720 27956
rect 31484 27940 31536 27946
rect 31484 27882 31536 27888
rect 31392 27396 31444 27402
rect 31392 27338 31444 27344
rect 31404 26382 31432 27338
rect 31392 26376 31444 26382
rect 31392 26318 31444 26324
rect 31300 25968 31352 25974
rect 31300 25910 31352 25916
rect 31392 25968 31444 25974
rect 31392 25910 31444 25916
rect 31208 23112 31260 23118
rect 31208 23054 31260 23060
rect 31300 23112 31352 23118
rect 31300 23054 31352 23060
rect 31116 23044 31168 23050
rect 31116 22986 31168 22992
rect 31022 22264 31078 22273
rect 31022 22199 31078 22208
rect 30932 21344 30984 21350
rect 30932 21286 30984 21292
rect 30840 20528 30892 20534
rect 30760 20488 30840 20516
rect 30656 20256 30708 20262
rect 30656 20198 30708 20204
rect 30472 19780 30524 19786
rect 30472 19722 30524 19728
rect 30288 19508 30340 19514
rect 30288 19450 30340 19456
rect 30208 19366 30420 19394
rect 30392 19334 30420 19366
rect 30104 19304 30156 19310
rect 30104 19246 30156 19252
rect 30196 19304 30248 19310
rect 30196 19246 30248 19252
rect 30300 19306 30420 19334
rect 30104 19168 30156 19174
rect 30104 19110 30156 19116
rect 30116 18442 30144 19110
rect 30208 18630 30236 19246
rect 30300 18766 30328 19306
rect 30564 18964 30616 18970
rect 30564 18906 30616 18912
rect 30288 18760 30340 18766
rect 30288 18702 30340 18708
rect 30196 18624 30248 18630
rect 30196 18566 30248 18572
rect 30116 18414 30236 18442
rect 30012 18216 30064 18222
rect 30012 18158 30064 18164
rect 30012 16516 30064 16522
rect 30012 16458 30064 16464
rect 30024 16250 30052 16458
rect 30012 16244 30064 16250
rect 30012 16186 30064 16192
rect 30024 15638 30052 16186
rect 30012 15632 30064 15638
rect 30012 15574 30064 15580
rect 29920 15564 29972 15570
rect 29920 15506 29972 15512
rect 30208 15502 30236 18414
rect 30300 16153 30328 18702
rect 30470 18184 30526 18193
rect 30470 18119 30526 18128
rect 30380 17128 30432 17134
rect 30380 17070 30432 17076
rect 30392 16425 30420 17070
rect 30378 16416 30434 16425
rect 30378 16351 30434 16360
rect 30378 16280 30434 16289
rect 30484 16250 30512 18119
rect 30378 16215 30434 16224
rect 30472 16244 30524 16250
rect 30392 16182 30420 16215
rect 30472 16186 30524 16192
rect 30380 16176 30432 16182
rect 30286 16144 30342 16153
rect 30380 16118 30432 16124
rect 30286 16079 30342 16088
rect 30300 15910 30328 16079
rect 30288 15904 30340 15910
rect 30288 15846 30340 15852
rect 29828 15496 29880 15502
rect 29828 15438 29880 15444
rect 30196 15496 30248 15502
rect 30196 15438 30248 15444
rect 30208 15366 30236 15438
rect 30196 15360 30248 15366
rect 30196 15302 30248 15308
rect 30288 15360 30340 15366
rect 30288 15302 30340 15308
rect 30380 15360 30432 15366
rect 30380 15302 30432 15308
rect 30300 15094 30328 15302
rect 30288 15088 30340 15094
rect 30288 15030 30340 15036
rect 30300 13870 30328 15030
rect 30392 14278 30420 15302
rect 30484 14414 30512 16186
rect 30576 16114 30604 18906
rect 30668 16289 30696 20198
rect 30760 19224 30788 20488
rect 30840 20470 30892 20476
rect 30932 20324 30984 20330
rect 30932 20266 30984 20272
rect 30840 20256 30892 20262
rect 30840 20198 30892 20204
rect 30852 19378 30880 20198
rect 30944 19417 30972 20266
rect 31036 19514 31064 22199
rect 31024 19508 31076 19514
rect 31024 19450 31076 19456
rect 30930 19408 30986 19417
rect 30840 19372 30892 19378
rect 30930 19343 30986 19352
rect 31024 19372 31076 19378
rect 30840 19314 30892 19320
rect 30840 19236 30892 19242
rect 30760 19196 30840 19224
rect 30760 16454 30788 19196
rect 30840 19178 30892 19184
rect 30944 18834 30972 19343
rect 31024 19314 31076 19320
rect 31036 18902 31064 19314
rect 31024 18896 31076 18902
rect 31024 18838 31076 18844
rect 30932 18828 30984 18834
rect 30932 18770 30984 18776
rect 30932 18692 30984 18698
rect 31036 18680 31064 18838
rect 30984 18652 31064 18680
rect 30932 18634 30984 18640
rect 30932 17808 30984 17814
rect 30932 17750 30984 17756
rect 30748 16448 30800 16454
rect 30748 16390 30800 16396
rect 30654 16280 30710 16289
rect 30654 16215 30710 16224
rect 30564 16108 30616 16114
rect 30564 16050 30616 16056
rect 30472 14408 30524 14414
rect 30470 14376 30472 14385
rect 30524 14376 30526 14385
rect 30470 14311 30526 14320
rect 30576 14278 30604 16050
rect 30380 14272 30432 14278
rect 30380 14214 30432 14220
rect 30564 14272 30616 14278
rect 30564 14214 30616 14220
rect 30288 13864 30340 13870
rect 30288 13806 30340 13812
rect 30196 13320 30248 13326
rect 30196 13262 30248 13268
rect 30288 13320 30340 13326
rect 30288 13262 30340 13268
rect 30208 13025 30236 13262
rect 30194 13016 30250 13025
rect 29736 12980 29788 12986
rect 29736 12922 29788 12928
rect 30104 12980 30156 12986
rect 30194 12951 30250 12960
rect 30104 12922 30156 12928
rect 29920 12912 29972 12918
rect 29920 12854 29972 12860
rect 29736 12776 29788 12782
rect 29734 12744 29736 12753
rect 29788 12744 29790 12753
rect 29734 12679 29790 12688
rect 29734 12336 29790 12345
rect 29734 12271 29790 12280
rect 29748 11098 29776 12271
rect 29932 12238 29960 12854
rect 30116 12850 30144 12922
rect 30104 12844 30156 12850
rect 30104 12786 30156 12792
rect 30012 12708 30064 12714
rect 30012 12650 30064 12656
rect 30024 12306 30052 12650
rect 30012 12300 30064 12306
rect 30012 12242 30064 12248
rect 29920 12232 29972 12238
rect 29920 12174 29972 12180
rect 29748 11070 29960 11098
rect 30024 11082 30052 12242
rect 30104 12232 30156 12238
rect 30104 12174 30156 12180
rect 30116 11762 30144 12174
rect 30208 11830 30236 12951
rect 30300 12782 30328 13262
rect 30288 12776 30340 12782
rect 30288 12718 30340 12724
rect 30392 12646 30420 14214
rect 30576 13938 30604 14214
rect 30564 13932 30616 13938
rect 30564 13874 30616 13880
rect 30472 13524 30524 13530
rect 30472 13466 30524 13472
rect 30484 12850 30512 13466
rect 30472 12844 30524 12850
rect 30472 12786 30524 12792
rect 30484 12753 30512 12786
rect 30470 12744 30526 12753
rect 30470 12679 30526 12688
rect 30380 12640 30432 12646
rect 30380 12582 30432 12588
rect 30472 12640 30524 12646
rect 30472 12582 30524 12588
rect 30484 12481 30512 12582
rect 30470 12472 30526 12481
rect 30470 12407 30526 12416
rect 30196 11824 30248 11830
rect 30196 11766 30248 11772
rect 30104 11756 30156 11762
rect 30104 11698 30156 11704
rect 29828 11008 29880 11014
rect 29748 10968 29828 10996
rect 29644 10736 29696 10742
rect 29644 10678 29696 10684
rect 29472 10220 29592 10248
rect 29368 7540 29420 7546
rect 29368 7482 29420 7488
rect 29276 6792 29328 6798
rect 29276 6734 29328 6740
rect 29184 6452 29236 6458
rect 29184 6394 29236 6400
rect 29196 5710 29224 6394
rect 29380 6390 29408 7482
rect 29472 6730 29500 10220
rect 29550 10160 29606 10169
rect 29550 10095 29552 10104
rect 29604 10095 29606 10104
rect 29552 10066 29604 10072
rect 29748 9674 29776 10968
rect 29828 10950 29880 10956
rect 29828 10668 29880 10674
rect 29828 10610 29880 10616
rect 29840 10062 29868 10610
rect 29828 10056 29880 10062
rect 29828 9998 29880 10004
rect 29656 9646 29776 9674
rect 29840 9654 29868 9998
rect 29828 9648 29880 9654
rect 29656 8480 29684 9646
rect 29828 9590 29880 9596
rect 29828 9512 29880 9518
rect 29828 9454 29880 9460
rect 29734 9072 29790 9081
rect 29734 9007 29790 9016
rect 29748 8974 29776 9007
rect 29736 8968 29788 8974
rect 29736 8910 29788 8916
rect 29748 8673 29776 8910
rect 29734 8664 29790 8673
rect 29734 8599 29790 8608
rect 29840 8566 29868 9454
rect 29828 8560 29880 8566
rect 29828 8502 29880 8508
rect 29736 8492 29788 8498
rect 29656 8452 29736 8480
rect 29656 7886 29684 8452
rect 29736 8434 29788 8440
rect 29828 8288 29880 8294
rect 29828 8230 29880 8236
rect 29840 7886 29868 8230
rect 29644 7880 29696 7886
rect 29644 7822 29696 7828
rect 29828 7880 29880 7886
rect 29828 7822 29880 7828
rect 29550 7576 29606 7585
rect 29550 7511 29606 7520
rect 29564 7478 29592 7511
rect 29552 7472 29604 7478
rect 29552 7414 29604 7420
rect 29460 6724 29512 6730
rect 29460 6666 29512 6672
rect 29368 6384 29420 6390
rect 29368 6326 29420 6332
rect 29472 6118 29500 6666
rect 29564 6458 29592 7414
rect 29932 6798 29960 11070
rect 30012 11076 30064 11082
rect 30012 11018 30064 11024
rect 30116 10062 30144 11698
rect 30208 11218 30236 11766
rect 30576 11694 30604 13874
rect 30564 11688 30616 11694
rect 30564 11630 30616 11636
rect 30196 11212 30248 11218
rect 30196 11154 30248 11160
rect 30104 10056 30156 10062
rect 30024 10016 30104 10044
rect 30024 8430 30052 10016
rect 30104 9998 30156 10004
rect 30104 9444 30156 9450
rect 30104 9386 30156 9392
rect 30116 8974 30144 9386
rect 30104 8968 30156 8974
rect 30104 8910 30156 8916
rect 30012 8424 30064 8430
rect 30012 8366 30064 8372
rect 30208 8294 30236 11154
rect 30564 11144 30616 11150
rect 30564 11086 30616 11092
rect 30288 11076 30340 11082
rect 30288 11018 30340 11024
rect 30300 10674 30328 11018
rect 30472 11008 30524 11014
rect 30472 10950 30524 10956
rect 30288 10668 30340 10674
rect 30288 10610 30340 10616
rect 30484 9926 30512 10950
rect 30472 9920 30524 9926
rect 30472 9862 30524 9868
rect 30380 9580 30432 9586
rect 30380 9522 30432 9528
rect 30288 9444 30340 9450
rect 30288 9386 30340 9392
rect 30196 8288 30248 8294
rect 30196 8230 30248 8236
rect 30300 8090 30328 9386
rect 30392 9382 30420 9522
rect 30380 9376 30432 9382
rect 30380 9318 30432 9324
rect 30472 9376 30524 9382
rect 30472 9318 30524 9324
rect 30484 9110 30512 9318
rect 30576 9110 30604 11086
rect 30668 10418 30696 16215
rect 30760 16114 30788 16390
rect 30748 16108 30800 16114
rect 30748 16050 30800 16056
rect 30840 15904 30892 15910
rect 30840 15846 30892 15852
rect 30852 15502 30880 15846
rect 30840 15496 30892 15502
rect 30840 15438 30892 15444
rect 30748 15428 30800 15434
rect 30748 15370 30800 15376
rect 30760 13870 30788 15370
rect 30748 13864 30800 13870
rect 30748 13806 30800 13812
rect 30748 13728 30800 13734
rect 30748 13670 30800 13676
rect 30760 12238 30788 13670
rect 30944 13190 30972 17750
rect 31024 17672 31076 17678
rect 31024 17614 31076 17620
rect 31036 16046 31064 17614
rect 31128 16164 31156 22986
rect 31220 20398 31248 23054
rect 31312 22438 31340 23054
rect 31404 22642 31432 25910
rect 31496 23730 31524 27882
rect 31576 27124 31628 27130
rect 31576 27066 31628 27072
rect 31588 26382 31616 27066
rect 31576 26376 31628 26382
rect 31680 26353 31708 27950
rect 31864 27826 31892 29446
rect 31956 28626 31984 29446
rect 32220 29028 32272 29034
rect 32220 28970 32272 28976
rect 31944 28620 31996 28626
rect 31944 28562 31996 28568
rect 31956 27946 31984 28562
rect 32232 28558 32260 28970
rect 32220 28552 32272 28558
rect 32220 28494 32272 28500
rect 31944 27940 31996 27946
rect 31944 27882 31996 27888
rect 32128 27872 32180 27878
rect 31864 27798 32076 27826
rect 32128 27814 32180 27820
rect 31852 27600 31904 27606
rect 31852 27542 31904 27548
rect 31864 27112 31892 27542
rect 31864 27084 31984 27112
rect 31956 26994 31984 27084
rect 31760 26988 31812 26994
rect 31760 26930 31812 26936
rect 31944 26988 31996 26994
rect 31944 26930 31996 26936
rect 31772 26586 31800 26930
rect 31760 26580 31812 26586
rect 31760 26522 31812 26528
rect 31956 26450 31984 26930
rect 32048 26926 32076 27798
rect 32140 27538 32168 27814
rect 32324 27606 32352 30194
rect 32508 30161 32536 31894
rect 32956 31816 33008 31822
rect 32956 31758 33008 31764
rect 32772 31748 32824 31754
rect 32772 31690 32824 31696
rect 32784 31346 32812 31690
rect 32772 31340 32824 31346
rect 32772 31282 32824 31288
rect 32680 30796 32732 30802
rect 32680 30738 32732 30744
rect 32588 30660 32640 30666
rect 32588 30602 32640 30608
rect 32494 30152 32550 30161
rect 32494 30087 32550 30096
rect 32404 29164 32456 29170
rect 32508 29152 32536 30087
rect 32456 29124 32536 29152
rect 32404 29106 32456 29112
rect 32404 28756 32456 28762
rect 32404 28698 32456 28704
rect 32416 28082 32444 28698
rect 32508 28218 32536 29124
rect 32600 28762 32628 30602
rect 32692 30394 32720 30738
rect 32680 30388 32732 30394
rect 32680 30330 32732 30336
rect 32680 30048 32732 30054
rect 32680 29990 32732 29996
rect 32692 29170 32720 29990
rect 32772 29640 32824 29646
rect 32772 29582 32824 29588
rect 32864 29640 32916 29646
rect 32864 29582 32916 29588
rect 32784 29306 32812 29582
rect 32772 29300 32824 29306
rect 32772 29242 32824 29248
rect 32876 29186 32904 29582
rect 32680 29164 32732 29170
rect 32680 29106 32732 29112
rect 32784 29158 32904 29186
rect 32588 28756 32640 28762
rect 32588 28698 32640 28704
rect 32680 28620 32732 28626
rect 32680 28562 32732 28568
rect 32588 28552 32640 28558
rect 32588 28494 32640 28500
rect 32496 28212 32548 28218
rect 32496 28154 32548 28160
rect 32404 28076 32456 28082
rect 32404 28018 32456 28024
rect 32416 27860 32444 28018
rect 32508 27962 32536 28154
rect 32600 28082 32628 28494
rect 32588 28076 32640 28082
rect 32588 28018 32640 28024
rect 32508 27934 32628 27962
rect 32416 27832 32536 27860
rect 32312 27600 32364 27606
rect 32312 27542 32364 27548
rect 32128 27532 32180 27538
rect 32128 27474 32180 27480
rect 32128 27396 32180 27402
rect 32404 27396 32456 27402
rect 32128 27338 32180 27344
rect 32232 27356 32404 27384
rect 32140 27062 32168 27338
rect 32128 27056 32180 27062
rect 32128 26998 32180 27004
rect 32036 26920 32088 26926
rect 32036 26862 32088 26868
rect 31944 26444 31996 26450
rect 31944 26386 31996 26392
rect 31852 26376 31904 26382
rect 31576 26318 31628 26324
rect 31666 26344 31722 26353
rect 31666 26279 31722 26288
rect 31850 26344 31852 26353
rect 31904 26344 31906 26353
rect 31850 26279 31906 26288
rect 31852 26240 31904 26246
rect 31852 26182 31904 26188
rect 31576 25900 31628 25906
rect 31576 25842 31628 25848
rect 31484 23724 31536 23730
rect 31484 23666 31536 23672
rect 31484 23588 31536 23594
rect 31484 23530 31536 23536
rect 31392 22636 31444 22642
rect 31392 22578 31444 22584
rect 31300 22432 31352 22438
rect 31300 22374 31352 22380
rect 31300 21344 31352 21350
rect 31300 21286 31352 21292
rect 31208 20392 31260 20398
rect 31208 20334 31260 20340
rect 31220 19854 31248 20334
rect 31208 19848 31260 19854
rect 31208 19790 31260 19796
rect 31208 19168 31260 19174
rect 31208 19110 31260 19116
rect 31220 18766 31248 19110
rect 31208 18760 31260 18766
rect 31208 18702 31260 18708
rect 31312 17814 31340 21286
rect 31404 19922 31432 22578
rect 31496 21622 31524 23530
rect 31588 23526 31616 25842
rect 31864 25294 31892 26182
rect 31956 25702 31984 26386
rect 32048 26382 32076 26862
rect 32036 26376 32088 26382
rect 32036 26318 32088 26324
rect 31944 25696 31996 25702
rect 31944 25638 31996 25644
rect 32128 25696 32180 25702
rect 32128 25638 32180 25644
rect 31944 25492 31996 25498
rect 31944 25434 31996 25440
rect 31956 25401 31984 25434
rect 31942 25392 31998 25401
rect 31942 25327 31998 25336
rect 32140 25294 32168 25638
rect 31760 25288 31812 25294
rect 31760 25230 31812 25236
rect 31852 25288 31904 25294
rect 31852 25230 31904 25236
rect 32128 25288 32180 25294
rect 32128 25230 32180 25236
rect 31772 24818 31800 25230
rect 32128 25152 32180 25158
rect 32128 25094 32180 25100
rect 31760 24812 31812 24818
rect 31760 24754 31812 24760
rect 31576 23520 31628 23526
rect 31576 23462 31628 23468
rect 31772 23118 31800 24754
rect 31852 24744 31904 24750
rect 31852 24686 31904 24692
rect 31760 23112 31812 23118
rect 31760 23054 31812 23060
rect 31668 22976 31720 22982
rect 31588 22924 31668 22930
rect 31588 22918 31720 22924
rect 31588 22902 31708 22918
rect 31588 22574 31616 22902
rect 31772 22642 31800 23054
rect 31864 22817 31892 24686
rect 31944 24676 31996 24682
rect 31944 24618 31996 24624
rect 31850 22808 31906 22817
rect 31850 22743 31852 22752
rect 31904 22743 31906 22752
rect 31852 22714 31904 22720
rect 31668 22636 31720 22642
rect 31668 22578 31720 22584
rect 31760 22636 31812 22642
rect 31760 22578 31812 22584
rect 31852 22636 31904 22642
rect 31852 22578 31904 22584
rect 31576 22568 31628 22574
rect 31576 22510 31628 22516
rect 31680 22234 31708 22578
rect 31864 22409 31892 22578
rect 31850 22400 31906 22409
rect 31850 22335 31906 22344
rect 31668 22228 31720 22234
rect 31668 22170 31720 22176
rect 31484 21616 31536 21622
rect 31484 21558 31536 21564
rect 31852 21548 31904 21554
rect 31852 21490 31904 21496
rect 31668 21344 31720 21350
rect 31668 21286 31720 21292
rect 31484 20460 31536 20466
rect 31484 20402 31536 20408
rect 31576 20460 31628 20466
rect 31576 20402 31628 20408
rect 31496 20330 31524 20402
rect 31484 20324 31536 20330
rect 31484 20266 31536 20272
rect 31588 20262 31616 20402
rect 31680 20346 31708 21286
rect 31864 20942 31892 21490
rect 31852 20936 31904 20942
rect 31852 20878 31904 20884
rect 31760 20528 31812 20534
rect 31758 20496 31760 20505
rect 31812 20496 31814 20505
rect 31864 20466 31892 20878
rect 31758 20431 31814 20440
rect 31852 20460 31904 20466
rect 31852 20402 31904 20408
rect 31760 20392 31812 20398
rect 31680 20340 31760 20346
rect 31680 20334 31812 20340
rect 31680 20318 31800 20334
rect 31576 20256 31628 20262
rect 31576 20198 31628 20204
rect 31392 19916 31444 19922
rect 31392 19858 31444 19864
rect 31300 17808 31352 17814
rect 31300 17750 31352 17756
rect 31300 17604 31352 17610
rect 31404 17592 31432 19858
rect 31680 19854 31708 20318
rect 31760 20256 31812 20262
rect 31760 20198 31812 20204
rect 31484 19848 31536 19854
rect 31484 19790 31536 19796
rect 31668 19848 31720 19854
rect 31668 19790 31720 19796
rect 31496 18766 31524 19790
rect 31576 19712 31628 19718
rect 31628 19660 31708 19666
rect 31576 19654 31708 19660
rect 31588 19638 31708 19654
rect 31680 19514 31708 19638
rect 31668 19508 31720 19514
rect 31668 19450 31720 19456
rect 31668 18896 31720 18902
rect 31668 18838 31720 18844
rect 31484 18760 31536 18766
rect 31484 18702 31536 18708
rect 31496 18086 31524 18702
rect 31576 18420 31628 18426
rect 31576 18362 31628 18368
rect 31484 18080 31536 18086
rect 31484 18022 31536 18028
rect 31496 17678 31524 18022
rect 31484 17672 31536 17678
rect 31484 17614 31536 17620
rect 31352 17564 31432 17592
rect 31300 17546 31352 17552
rect 31312 17513 31340 17546
rect 31298 17504 31354 17513
rect 31298 17439 31354 17448
rect 31392 16584 31444 16590
rect 31392 16526 31444 16532
rect 31300 16176 31352 16182
rect 31128 16136 31300 16164
rect 31024 16040 31076 16046
rect 31024 15982 31076 15988
rect 31024 15496 31076 15502
rect 31024 15438 31076 15444
rect 31036 15162 31064 15438
rect 31024 15156 31076 15162
rect 31024 15098 31076 15104
rect 31024 14476 31076 14482
rect 31024 14418 31076 14424
rect 30932 13184 30984 13190
rect 30932 13126 30984 13132
rect 30838 13016 30894 13025
rect 30838 12951 30894 12960
rect 30852 12850 30880 12951
rect 30944 12918 30972 13126
rect 30932 12912 30984 12918
rect 30932 12854 30984 12860
rect 30840 12844 30892 12850
rect 30840 12786 30892 12792
rect 30944 12442 30972 12854
rect 30932 12436 30984 12442
rect 30932 12378 30984 12384
rect 30748 12232 30800 12238
rect 30748 12174 30800 12180
rect 30760 11082 30788 12174
rect 30840 12164 30892 12170
rect 30840 12106 30892 12112
rect 30852 11150 30880 12106
rect 30932 11348 30984 11354
rect 30932 11290 30984 11296
rect 30944 11257 30972 11290
rect 30930 11248 30986 11257
rect 30930 11183 30986 11192
rect 30840 11144 30892 11150
rect 30840 11086 30892 11092
rect 30748 11076 30800 11082
rect 30748 11018 30800 11024
rect 30840 10668 30892 10674
rect 30840 10610 30892 10616
rect 30668 10390 30788 10418
rect 30656 10260 30708 10266
rect 30656 10202 30708 10208
rect 30472 9104 30524 9110
rect 30472 9046 30524 9052
rect 30564 9104 30616 9110
rect 30564 9046 30616 9052
rect 30380 8900 30432 8906
rect 30380 8842 30432 8848
rect 30392 8537 30420 8842
rect 30378 8528 30434 8537
rect 30378 8463 30434 8472
rect 30576 8480 30604 9046
rect 30668 8974 30696 10202
rect 30760 10062 30788 10390
rect 30748 10056 30800 10062
rect 30748 9998 30800 10004
rect 30760 9722 30788 9998
rect 30852 9761 30880 10610
rect 30932 10260 30984 10266
rect 31036 10248 31064 14418
rect 31128 11014 31156 16136
rect 31300 16118 31352 16124
rect 31404 16114 31432 16526
rect 31496 16114 31524 17614
rect 31588 16697 31616 18362
rect 31574 16688 31630 16697
rect 31574 16623 31630 16632
rect 31392 16108 31444 16114
rect 31392 16050 31444 16056
rect 31484 16108 31536 16114
rect 31484 16050 31536 16056
rect 31300 15972 31352 15978
rect 31300 15914 31352 15920
rect 31208 15496 31260 15502
rect 31206 15464 31208 15473
rect 31260 15464 31262 15473
rect 31206 15399 31262 15408
rect 31208 12708 31260 12714
rect 31208 12650 31260 12656
rect 31220 11898 31248 12650
rect 31312 12434 31340 15914
rect 31404 13938 31432 16050
rect 31496 15473 31524 16050
rect 31576 16040 31628 16046
rect 31576 15982 31628 15988
rect 31588 15502 31616 15982
rect 31576 15496 31628 15502
rect 31482 15464 31538 15473
rect 31576 15438 31628 15444
rect 31482 15399 31538 15408
rect 31496 15366 31524 15399
rect 31484 15360 31536 15366
rect 31484 15302 31536 15308
rect 31484 14952 31536 14958
rect 31484 14894 31536 14900
rect 31392 13932 31444 13938
rect 31392 13874 31444 13880
rect 31496 13326 31524 14894
rect 31576 13932 31628 13938
rect 31576 13874 31628 13880
rect 31484 13320 31536 13326
rect 31484 13262 31536 13268
rect 31392 13252 31444 13258
rect 31392 13194 31444 13200
rect 31404 12918 31432 13194
rect 31484 13184 31536 13190
rect 31484 13126 31536 13132
rect 31392 12912 31444 12918
rect 31392 12854 31444 12860
rect 31312 12406 31432 12434
rect 31300 12096 31352 12102
rect 31300 12038 31352 12044
rect 31208 11892 31260 11898
rect 31208 11834 31260 11840
rect 31116 11008 31168 11014
rect 31116 10950 31168 10956
rect 31220 10810 31248 11834
rect 31208 10804 31260 10810
rect 31208 10746 31260 10752
rect 31116 10668 31168 10674
rect 31116 10610 31168 10616
rect 31128 10470 31156 10610
rect 31206 10568 31262 10577
rect 31206 10503 31262 10512
rect 31116 10464 31168 10470
rect 31116 10406 31168 10412
rect 30984 10220 31064 10248
rect 30932 10202 30984 10208
rect 31116 10192 31168 10198
rect 31116 10134 31168 10140
rect 30932 9920 30984 9926
rect 30932 9862 30984 9868
rect 30838 9752 30894 9761
rect 30748 9716 30800 9722
rect 30838 9687 30894 9696
rect 30748 9658 30800 9664
rect 30748 9444 30800 9450
rect 30748 9386 30800 9392
rect 30656 8968 30708 8974
rect 30656 8910 30708 8916
rect 30656 8492 30708 8498
rect 30576 8452 30656 8480
rect 30656 8434 30708 8440
rect 30380 8288 30432 8294
rect 30380 8230 30432 8236
rect 30392 8090 30420 8230
rect 30288 8084 30340 8090
rect 30288 8026 30340 8032
rect 30380 8084 30432 8090
rect 30380 8026 30432 8032
rect 30300 7886 30328 8026
rect 30288 7880 30340 7886
rect 30288 7822 30340 7828
rect 30300 7546 30328 7822
rect 30196 7540 30248 7546
rect 30196 7482 30248 7488
rect 30288 7540 30340 7546
rect 30288 7482 30340 7488
rect 30208 6798 30236 7482
rect 30668 7410 30696 8434
rect 30760 8430 30788 9386
rect 30748 8424 30800 8430
rect 30748 8366 30800 8372
rect 30760 8090 30788 8366
rect 30748 8084 30800 8090
rect 30748 8026 30800 8032
rect 30852 7750 30880 9687
rect 30944 9654 30972 9862
rect 30932 9648 30984 9654
rect 30932 9590 30984 9596
rect 31024 9580 31076 9586
rect 31024 9522 31076 9528
rect 30932 8832 30984 8838
rect 30932 8774 30984 8780
rect 30944 8430 30972 8774
rect 30932 8424 30984 8430
rect 30932 8366 30984 8372
rect 31036 8294 31064 9522
rect 31128 9178 31156 10134
rect 31116 9172 31168 9178
rect 31116 9114 31168 9120
rect 31128 9081 31156 9114
rect 31114 9072 31170 9081
rect 31114 9007 31170 9016
rect 31128 8974 31156 9007
rect 31220 8974 31248 10503
rect 31116 8968 31168 8974
rect 31116 8910 31168 8916
rect 31208 8968 31260 8974
rect 31208 8910 31260 8916
rect 31220 8634 31248 8910
rect 31208 8628 31260 8634
rect 31208 8570 31260 8576
rect 31024 8288 31076 8294
rect 31024 8230 31076 8236
rect 31036 7886 31064 8230
rect 31024 7880 31076 7886
rect 31024 7822 31076 7828
rect 30840 7744 30892 7750
rect 30840 7686 30892 7692
rect 31036 7410 31064 7822
rect 30656 7404 30708 7410
rect 30656 7346 30708 7352
rect 31024 7404 31076 7410
rect 31024 7346 31076 7352
rect 31220 7206 31248 8570
rect 31312 7750 31340 12038
rect 31404 10538 31432 12406
rect 31392 10532 31444 10538
rect 31392 10474 31444 10480
rect 31404 10198 31432 10474
rect 31392 10192 31444 10198
rect 31392 10134 31444 10140
rect 31392 10056 31444 10062
rect 31392 9998 31444 10004
rect 31404 9926 31432 9998
rect 31392 9920 31444 9926
rect 31392 9862 31444 9868
rect 31392 9648 31444 9654
rect 31392 9590 31444 9596
rect 31404 7954 31432 9590
rect 31496 9178 31524 13126
rect 31588 10577 31616 13874
rect 31680 11880 31708 18838
rect 31772 18766 31800 20198
rect 31760 18760 31812 18766
rect 31760 18702 31812 18708
rect 31852 18692 31904 18698
rect 31852 18634 31904 18640
rect 31864 18358 31892 18634
rect 31852 18352 31904 18358
rect 31852 18294 31904 18300
rect 31850 17912 31906 17921
rect 31850 17847 31906 17856
rect 31864 17678 31892 17847
rect 31852 17672 31904 17678
rect 31852 17614 31904 17620
rect 31956 17202 31984 24618
rect 32036 23180 32088 23186
rect 32036 23122 32088 23128
rect 32048 22778 32076 23122
rect 32036 22772 32088 22778
rect 32036 22714 32088 22720
rect 32140 22658 32168 25094
rect 32048 22630 32168 22658
rect 32048 20466 32076 22630
rect 32128 22500 32180 22506
rect 32128 22442 32180 22448
rect 32140 22098 32168 22442
rect 32128 22092 32180 22098
rect 32128 22034 32180 22040
rect 32232 22030 32260 27356
rect 32404 27338 32456 27344
rect 32310 27024 32366 27033
rect 32310 26959 32366 26968
rect 32324 26790 32352 26959
rect 32508 26897 32536 27832
rect 32600 27606 32628 27934
rect 32588 27600 32640 27606
rect 32588 27542 32640 27548
rect 32600 27470 32628 27542
rect 32588 27464 32640 27470
rect 32588 27406 32640 27412
rect 32588 26920 32640 26926
rect 32494 26888 32550 26897
rect 32588 26862 32640 26868
rect 32494 26823 32550 26832
rect 32312 26784 32364 26790
rect 32312 26726 32364 26732
rect 32324 26625 32352 26726
rect 32310 26616 32366 26625
rect 32310 26551 32366 26560
rect 32494 26616 32550 26625
rect 32494 26551 32550 26560
rect 32508 26518 32536 26551
rect 32496 26512 32548 26518
rect 32496 26454 32548 26460
rect 32600 26382 32628 26862
rect 32404 26376 32456 26382
rect 32496 26376 32548 26382
rect 32404 26318 32456 26324
rect 32494 26344 32496 26353
rect 32588 26376 32640 26382
rect 32548 26344 32550 26353
rect 32416 26194 32444 26318
rect 32588 26318 32640 26324
rect 32494 26279 32550 26288
rect 32416 26166 32628 26194
rect 32496 25900 32548 25906
rect 32496 25842 32548 25848
rect 32404 25152 32456 25158
rect 32404 25094 32456 25100
rect 32416 24857 32444 25094
rect 32508 24993 32536 25842
rect 32600 25158 32628 26166
rect 32588 25152 32640 25158
rect 32588 25094 32640 25100
rect 32494 24984 32550 24993
rect 32494 24919 32550 24928
rect 32402 24848 32458 24857
rect 32402 24783 32458 24792
rect 32496 24404 32548 24410
rect 32496 24346 32548 24352
rect 32312 23656 32364 23662
rect 32310 23624 32312 23633
rect 32364 23624 32366 23633
rect 32310 23559 32366 23568
rect 32312 23520 32364 23526
rect 32312 23462 32364 23468
rect 32220 22024 32272 22030
rect 32220 21966 32272 21972
rect 32232 21350 32260 21966
rect 32220 21344 32272 21350
rect 32220 21286 32272 21292
rect 32220 20936 32272 20942
rect 32220 20878 32272 20884
rect 32036 20460 32088 20466
rect 32036 20402 32088 20408
rect 32232 20262 32260 20878
rect 32220 20256 32272 20262
rect 32220 20198 32272 20204
rect 32220 18624 32272 18630
rect 32220 18566 32272 18572
rect 32128 18080 32180 18086
rect 32128 18022 32180 18028
rect 32140 17678 32168 18022
rect 32128 17672 32180 17678
rect 32128 17614 32180 17620
rect 31944 17196 31996 17202
rect 31944 17138 31996 17144
rect 31944 16448 31996 16454
rect 31944 16390 31996 16396
rect 31852 15700 31904 15706
rect 31852 15642 31904 15648
rect 31864 15434 31892 15642
rect 31760 15428 31812 15434
rect 31760 15370 31812 15376
rect 31852 15428 31904 15434
rect 31852 15370 31904 15376
rect 31772 15162 31800 15370
rect 31760 15156 31812 15162
rect 31760 15098 31812 15104
rect 31864 15042 31892 15370
rect 31772 15014 31892 15042
rect 31772 13530 31800 15014
rect 31850 13560 31906 13569
rect 31760 13524 31812 13530
rect 31850 13495 31906 13504
rect 31760 13466 31812 13472
rect 31864 13462 31892 13495
rect 31852 13456 31904 13462
rect 31852 13398 31904 13404
rect 31852 13320 31904 13326
rect 31852 13262 31904 13268
rect 31864 12850 31892 13262
rect 31956 13258 31984 16390
rect 32128 15360 32180 15366
rect 32128 15302 32180 15308
rect 32036 14000 32088 14006
rect 32036 13942 32088 13948
rect 31944 13252 31996 13258
rect 31944 13194 31996 13200
rect 31760 12844 31812 12850
rect 31760 12786 31812 12792
rect 31852 12844 31904 12850
rect 31852 12786 31904 12792
rect 31772 12102 31800 12786
rect 31760 12096 31812 12102
rect 31760 12038 31812 12044
rect 31680 11852 31800 11880
rect 31668 11076 31720 11082
rect 31668 11018 31720 11024
rect 31574 10568 31630 10577
rect 31574 10503 31630 10512
rect 31574 9344 31630 9353
rect 31574 9279 31630 9288
rect 31484 9172 31536 9178
rect 31484 9114 31536 9120
rect 31496 8906 31524 9114
rect 31484 8900 31536 8906
rect 31484 8842 31536 8848
rect 31588 8498 31616 9279
rect 31576 8492 31628 8498
rect 31496 8452 31576 8480
rect 31496 7954 31524 8452
rect 31576 8434 31628 8440
rect 31576 8084 31628 8090
rect 31576 8026 31628 8032
rect 31392 7948 31444 7954
rect 31392 7890 31444 7896
rect 31484 7948 31536 7954
rect 31484 7890 31536 7896
rect 31300 7744 31352 7750
rect 31300 7686 31352 7692
rect 31404 7478 31432 7890
rect 31392 7472 31444 7478
rect 31392 7414 31444 7420
rect 31588 7342 31616 8026
rect 31680 7342 31708 11018
rect 31772 10266 31800 11852
rect 31852 11688 31904 11694
rect 31852 11630 31904 11636
rect 31864 10674 31892 11630
rect 31944 11552 31996 11558
rect 31944 11494 31996 11500
rect 31852 10668 31904 10674
rect 31852 10610 31904 10616
rect 31956 10538 31984 11494
rect 31944 10532 31996 10538
rect 31944 10474 31996 10480
rect 31760 10260 31812 10266
rect 31760 10202 31812 10208
rect 31772 8498 31800 10202
rect 32048 10062 32076 13942
rect 32140 13734 32168 15302
rect 32232 14006 32260 18566
rect 32220 14000 32272 14006
rect 32220 13942 32272 13948
rect 32128 13728 32180 13734
rect 32128 13670 32180 13676
rect 32218 13696 32274 13705
rect 32218 13631 32274 13640
rect 32128 13524 32180 13530
rect 32128 13466 32180 13472
rect 32140 11014 32168 13466
rect 32232 12850 32260 13631
rect 32220 12844 32272 12850
rect 32220 12786 32272 12792
rect 32220 11212 32272 11218
rect 32220 11154 32272 11160
rect 32128 11008 32180 11014
rect 32128 10950 32180 10956
rect 32232 10742 32260 11154
rect 32220 10736 32272 10742
rect 32220 10678 32272 10684
rect 32324 10674 32352 23462
rect 32404 22636 32456 22642
rect 32404 22578 32456 22584
rect 32416 21894 32444 22578
rect 32404 21888 32456 21894
rect 32404 21830 32456 21836
rect 32508 21010 32536 24346
rect 32692 22574 32720 28562
rect 32784 28014 32812 29158
rect 32864 29028 32916 29034
rect 32864 28970 32916 28976
rect 32772 28008 32824 28014
rect 32772 27950 32824 27956
rect 32784 27577 32812 27950
rect 32770 27568 32826 27577
rect 32770 27503 32826 27512
rect 32772 27464 32824 27470
rect 32772 27406 32824 27412
rect 32784 27334 32812 27406
rect 32772 27328 32824 27334
rect 32770 27296 32772 27305
rect 32824 27296 32826 27305
rect 32770 27231 32826 27240
rect 32772 26308 32824 26314
rect 32772 26250 32824 26256
rect 32680 22568 32732 22574
rect 32680 22510 32732 22516
rect 32692 22094 32720 22510
rect 32600 22066 32720 22094
rect 32496 21004 32548 21010
rect 32496 20946 32548 20952
rect 32600 20466 32628 22066
rect 32784 21536 32812 26250
rect 32876 25362 32904 28970
rect 32968 28626 32996 31758
rect 33060 29714 33088 32438
rect 33152 32026 33180 33254
rect 34256 33114 34284 33458
rect 38752 33448 38804 33454
rect 38752 33390 38804 33396
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 33232 33108 33284 33114
rect 33232 33050 33284 33056
rect 34244 33108 34296 33114
rect 34244 33050 34296 33056
rect 33140 32020 33192 32026
rect 33140 31962 33192 31968
rect 33244 31822 33272 33050
rect 34336 33040 34388 33046
rect 34336 32982 34388 32988
rect 33692 32904 33744 32910
rect 33692 32846 33744 32852
rect 33704 32502 33732 32846
rect 34348 32570 34376 32982
rect 37280 32904 37332 32910
rect 35806 32872 35862 32881
rect 35862 32842 36032 32858
rect 37280 32846 37332 32852
rect 35862 32836 36044 32842
rect 35862 32830 35992 32836
rect 35806 32807 35862 32816
rect 35992 32778 36044 32784
rect 36452 32836 36504 32842
rect 36452 32778 36504 32784
rect 34428 32768 34480 32774
rect 34428 32710 34480 32716
rect 34610 32736 34666 32745
rect 34336 32564 34388 32570
rect 34336 32506 34388 32512
rect 33692 32496 33744 32502
rect 33692 32438 33744 32444
rect 33968 32428 34020 32434
rect 33968 32370 34020 32376
rect 34152 32428 34204 32434
rect 34152 32370 34204 32376
rect 33232 31816 33284 31822
rect 33232 31758 33284 31764
rect 33784 31408 33836 31414
rect 33784 31350 33836 31356
rect 33324 31136 33376 31142
rect 33324 31078 33376 31084
rect 33600 31136 33652 31142
rect 33600 31078 33652 31084
rect 33336 30666 33364 31078
rect 33612 30938 33640 31078
rect 33600 30932 33652 30938
rect 33600 30874 33652 30880
rect 33692 30796 33744 30802
rect 33692 30738 33744 30744
rect 33324 30660 33376 30666
rect 33324 30602 33376 30608
rect 33140 30252 33192 30258
rect 33140 30194 33192 30200
rect 33048 29708 33100 29714
rect 33048 29650 33100 29656
rect 33048 29572 33100 29578
rect 33048 29514 33100 29520
rect 33060 29170 33088 29514
rect 33048 29164 33100 29170
rect 33048 29106 33100 29112
rect 32956 28620 33008 28626
rect 32956 28562 33008 28568
rect 32956 27532 33008 27538
rect 32956 27474 33008 27480
rect 32968 27334 32996 27474
rect 32956 27328 33008 27334
rect 32956 27270 33008 27276
rect 32864 25356 32916 25362
rect 32864 25298 32916 25304
rect 32968 24750 32996 27270
rect 33060 25294 33088 29106
rect 33152 28966 33180 30194
rect 33336 29646 33364 30602
rect 33600 30592 33652 30598
rect 33600 30534 33652 30540
rect 33506 30288 33562 30297
rect 33506 30223 33562 30232
rect 33414 30152 33470 30161
rect 33414 30087 33416 30096
rect 33468 30087 33470 30096
rect 33416 30058 33468 30064
rect 33428 29753 33456 30058
rect 33414 29744 33470 29753
rect 33520 29714 33548 30223
rect 33612 30054 33640 30534
rect 33704 30433 33732 30738
rect 33690 30424 33746 30433
rect 33690 30359 33746 30368
rect 33704 30326 33732 30359
rect 33692 30320 33744 30326
rect 33692 30262 33744 30268
rect 33600 30048 33652 30054
rect 33600 29990 33652 29996
rect 33612 29782 33640 29990
rect 33600 29776 33652 29782
rect 33600 29718 33652 29724
rect 33414 29679 33470 29688
rect 33508 29708 33560 29714
rect 33508 29650 33560 29656
rect 33324 29640 33376 29646
rect 33324 29582 33376 29588
rect 33232 29504 33284 29510
rect 33232 29446 33284 29452
rect 33140 28960 33192 28966
rect 33140 28902 33192 28908
rect 33140 27464 33192 27470
rect 33140 27406 33192 27412
rect 33152 26246 33180 27406
rect 33244 26761 33272 29446
rect 33520 29345 33548 29650
rect 33796 29510 33824 31350
rect 33876 30728 33928 30734
rect 33874 30696 33876 30705
rect 33928 30696 33930 30705
rect 33874 30631 33930 30640
rect 33876 29844 33928 29850
rect 33876 29786 33928 29792
rect 33888 29753 33916 29786
rect 33874 29744 33930 29753
rect 33874 29679 33930 29688
rect 33980 29646 34008 32370
rect 34164 31822 34192 32370
rect 34440 32366 34468 32710
rect 34610 32671 34666 32680
rect 34624 32502 34652 32671
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 36464 32570 36492 32778
rect 36452 32564 36504 32570
rect 36452 32506 36504 32512
rect 34612 32496 34664 32502
rect 34612 32438 34664 32444
rect 34428 32360 34480 32366
rect 34428 32302 34480 32308
rect 34624 32026 34652 32438
rect 37292 32434 37320 32846
rect 37280 32428 37332 32434
rect 37280 32370 37332 32376
rect 38200 32428 38252 32434
rect 38200 32370 38252 32376
rect 35992 32360 36044 32366
rect 34794 32328 34850 32337
rect 35992 32302 36044 32308
rect 36084 32360 36136 32366
rect 36084 32302 36136 32308
rect 37464 32360 37516 32366
rect 37464 32302 37516 32308
rect 37556 32360 37608 32366
rect 37556 32302 37608 32308
rect 37832 32360 37884 32366
rect 37832 32302 37884 32308
rect 34794 32263 34850 32272
rect 34808 32230 34836 32263
rect 34796 32224 34848 32230
rect 34796 32166 34848 32172
rect 34612 32020 34664 32026
rect 34612 31962 34664 31968
rect 34808 31890 34836 32166
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 36004 31890 36032 32302
rect 36096 32026 36124 32302
rect 37372 32292 37424 32298
rect 37372 32234 37424 32240
rect 36084 32020 36136 32026
rect 36084 31962 36136 31968
rect 36728 31952 36780 31958
rect 36728 31894 36780 31900
rect 34796 31884 34848 31890
rect 34796 31826 34848 31832
rect 34888 31884 34940 31890
rect 34888 31826 34940 31832
rect 35992 31884 36044 31890
rect 35992 31826 36044 31832
rect 36176 31884 36228 31890
rect 36176 31826 36228 31832
rect 34152 31816 34204 31822
rect 34152 31758 34204 31764
rect 34244 31680 34296 31686
rect 34244 31622 34296 31628
rect 34256 31414 34284 31622
rect 34900 31482 34928 31826
rect 35440 31680 35492 31686
rect 35440 31622 35492 31628
rect 35992 31680 36044 31686
rect 35992 31622 36044 31628
rect 35452 31482 35480 31622
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35594 31515 35902 31524
rect 34888 31476 34940 31482
rect 34888 31418 34940 31424
rect 35440 31476 35492 31482
rect 35440 31418 35492 31424
rect 34244 31408 34296 31414
rect 34244 31350 34296 31356
rect 34796 31408 34848 31414
rect 34796 31350 34848 31356
rect 34336 31340 34388 31346
rect 34336 31282 34388 31288
rect 34152 31136 34204 31142
rect 34152 31078 34204 31084
rect 34060 30184 34112 30190
rect 34060 30126 34112 30132
rect 34072 29889 34100 30126
rect 34164 30122 34192 31078
rect 34348 30734 34376 31282
rect 34808 31142 34836 31350
rect 36004 31346 36032 31622
rect 36188 31414 36216 31826
rect 36740 31822 36768 31894
rect 36728 31816 36780 31822
rect 36728 31758 36780 31764
rect 36544 31748 36596 31754
rect 36544 31690 36596 31696
rect 36176 31408 36228 31414
rect 36176 31350 36228 31356
rect 35992 31340 36044 31346
rect 35992 31282 36044 31288
rect 36360 31340 36412 31346
rect 36360 31282 36412 31288
rect 36452 31340 36504 31346
rect 36452 31282 36504 31288
rect 35440 31272 35492 31278
rect 35440 31214 35492 31220
rect 34796 31136 34848 31142
rect 34796 31078 34848 31084
rect 34610 30968 34666 30977
rect 34610 30903 34666 30912
rect 34704 30932 34756 30938
rect 34624 30870 34652 30903
rect 34704 30874 34756 30880
rect 34612 30864 34664 30870
rect 34612 30806 34664 30812
rect 34336 30728 34388 30734
rect 34336 30670 34388 30676
rect 34244 30592 34296 30598
rect 34244 30534 34296 30540
rect 34152 30116 34204 30122
rect 34152 30058 34204 30064
rect 34058 29880 34114 29889
rect 34058 29815 34114 29824
rect 33968 29640 34020 29646
rect 33968 29582 34020 29588
rect 33784 29504 33836 29510
rect 33784 29446 33836 29452
rect 33966 29472 34022 29481
rect 33966 29407 34022 29416
rect 33506 29336 33562 29345
rect 33506 29271 33562 29280
rect 33692 29300 33744 29306
rect 33692 29242 33744 29248
rect 33508 29232 33560 29238
rect 33704 29209 33732 29242
rect 33508 29174 33560 29180
rect 33690 29200 33746 29209
rect 33520 29073 33548 29174
rect 33690 29135 33692 29144
rect 33744 29135 33746 29144
rect 33874 29200 33930 29209
rect 33874 29135 33930 29144
rect 33692 29106 33744 29112
rect 33506 29064 33562 29073
rect 33888 29034 33916 29135
rect 33506 28999 33562 29008
rect 33876 29028 33928 29034
rect 33876 28970 33928 28976
rect 33600 28960 33652 28966
rect 33600 28902 33652 28908
rect 33612 28558 33640 28902
rect 33600 28552 33652 28558
rect 33600 28494 33652 28500
rect 33508 28484 33560 28490
rect 33508 28426 33560 28432
rect 33692 28484 33744 28490
rect 33692 28426 33744 28432
rect 33416 28416 33468 28422
rect 33416 28358 33468 28364
rect 33230 26752 33286 26761
rect 33230 26687 33286 26696
rect 33140 26240 33192 26246
rect 33140 26182 33192 26188
rect 33048 25288 33100 25294
rect 33048 25230 33100 25236
rect 32956 24744 33008 24750
rect 32956 24686 33008 24692
rect 33152 24698 33180 26182
rect 33244 24834 33272 26687
rect 33324 25288 33376 25294
rect 33324 25230 33376 25236
rect 33336 24954 33364 25230
rect 33324 24948 33376 24954
rect 33324 24890 33376 24896
rect 33244 24806 33364 24834
rect 33152 24670 33272 24698
rect 33140 24608 33192 24614
rect 33140 24550 33192 24556
rect 33152 23769 33180 24550
rect 33138 23760 33194 23769
rect 32956 23724 33008 23730
rect 33138 23695 33140 23704
rect 32956 23666 33008 23672
rect 33192 23695 33194 23704
rect 33140 23666 33192 23672
rect 32864 22976 32916 22982
rect 32864 22918 32916 22924
rect 32876 22642 32904 22918
rect 32864 22636 32916 22642
rect 32864 22578 32916 22584
rect 32864 22500 32916 22506
rect 32864 22442 32916 22448
rect 32876 22166 32904 22442
rect 32864 22160 32916 22166
rect 32864 22102 32916 22108
rect 32968 22098 32996 23666
rect 33048 23520 33100 23526
rect 33048 23462 33100 23468
rect 33060 23186 33088 23462
rect 33244 23304 33272 24670
rect 33152 23276 33272 23304
rect 33048 23180 33100 23186
rect 33048 23122 33100 23128
rect 33048 22636 33100 22642
rect 33048 22578 33100 22584
rect 33060 22438 33088 22578
rect 33048 22432 33100 22438
rect 33048 22374 33100 22380
rect 33152 22386 33180 23276
rect 33230 23216 33286 23225
rect 33336 23202 33364 24806
rect 33286 23174 33364 23202
rect 33428 23186 33456 28358
rect 33520 26382 33548 28426
rect 33600 26512 33652 26518
rect 33598 26480 33600 26489
rect 33652 26480 33654 26489
rect 33598 26415 33654 26424
rect 33508 26376 33560 26382
rect 33508 26318 33560 26324
rect 33612 25430 33640 26415
rect 33600 25424 33652 25430
rect 33600 25366 33652 25372
rect 33704 25294 33732 28426
rect 33784 27464 33836 27470
rect 33784 27406 33836 27412
rect 33692 25288 33744 25294
rect 33690 25256 33692 25265
rect 33744 25256 33746 25265
rect 33690 25191 33746 25200
rect 33600 25152 33652 25158
rect 33600 25094 33652 25100
rect 33508 24404 33560 24410
rect 33508 24346 33560 24352
rect 33520 23866 33548 24346
rect 33612 23866 33640 25094
rect 33508 23860 33560 23866
rect 33508 23802 33560 23808
rect 33600 23860 33652 23866
rect 33600 23802 33652 23808
rect 33796 23746 33824 27406
rect 33888 26518 33916 28970
rect 33876 26512 33928 26518
rect 33876 26454 33928 26460
rect 33876 26376 33928 26382
rect 33876 26318 33928 26324
rect 33888 25906 33916 26318
rect 33980 26042 34008 29407
rect 34072 29034 34100 29815
rect 34164 29646 34192 30058
rect 34256 29782 34284 30534
rect 34348 30054 34376 30670
rect 34336 30048 34388 30054
rect 34336 29990 34388 29996
rect 34244 29776 34296 29782
rect 34244 29718 34296 29724
rect 34152 29640 34204 29646
rect 34152 29582 34204 29588
rect 34244 29640 34296 29646
rect 34244 29582 34296 29588
rect 34152 29504 34204 29510
rect 34150 29472 34152 29481
rect 34204 29472 34206 29481
rect 34150 29407 34206 29416
rect 34152 29164 34204 29170
rect 34152 29106 34204 29112
rect 34164 29034 34192 29106
rect 34060 29028 34112 29034
rect 34060 28970 34112 28976
rect 34152 29028 34204 29034
rect 34152 28970 34204 28976
rect 34164 28762 34192 28970
rect 34256 28966 34284 29582
rect 34348 29238 34376 29990
rect 34716 29646 34744 30874
rect 34704 29640 34756 29646
rect 34704 29582 34756 29588
rect 34336 29232 34388 29238
rect 34336 29174 34388 29180
rect 34520 29232 34572 29238
rect 34520 29174 34572 29180
rect 34610 29200 34666 29209
rect 34244 28960 34296 28966
rect 34244 28902 34296 28908
rect 34152 28756 34204 28762
rect 34152 28698 34204 28704
rect 34256 28558 34284 28902
rect 34244 28552 34296 28558
rect 34244 28494 34296 28500
rect 34348 28490 34376 29174
rect 34428 28960 34480 28966
rect 34428 28902 34480 28908
rect 34440 28762 34468 28902
rect 34428 28756 34480 28762
rect 34428 28698 34480 28704
rect 34336 28484 34388 28490
rect 34336 28426 34388 28432
rect 34244 28416 34296 28422
rect 34164 28376 34244 28404
rect 34060 26852 34112 26858
rect 34060 26794 34112 26800
rect 33968 26036 34020 26042
rect 33968 25978 34020 25984
rect 33876 25900 33928 25906
rect 33876 25842 33928 25848
rect 33612 23718 33824 23746
rect 33416 23180 33468 23186
rect 33230 23151 33232 23160
rect 33284 23151 33286 23160
rect 33232 23122 33284 23128
rect 33416 23122 33468 23128
rect 33232 23044 33284 23050
rect 33232 22986 33284 22992
rect 33508 23044 33560 23050
rect 33508 22986 33560 22992
rect 33244 22930 33272 22986
rect 33244 22902 33456 22930
rect 33428 22642 33456 22902
rect 33416 22636 33468 22642
rect 33416 22578 33468 22584
rect 33520 22409 33548 22986
rect 33506 22400 33562 22409
rect 33152 22358 33272 22386
rect 33140 22228 33192 22234
rect 33140 22170 33192 22176
rect 32956 22092 33008 22098
rect 32956 22034 33008 22040
rect 32692 21508 32812 21536
rect 32496 20460 32548 20466
rect 32496 20402 32548 20408
rect 32588 20460 32640 20466
rect 32588 20402 32640 20408
rect 32404 19712 32456 19718
rect 32404 19654 32456 19660
rect 32416 18290 32444 19654
rect 32404 18284 32456 18290
rect 32404 18226 32456 18232
rect 32416 13530 32444 18226
rect 32508 15638 32536 20402
rect 32600 19446 32628 20402
rect 32588 19440 32640 19446
rect 32588 19382 32640 19388
rect 32692 17678 32720 21508
rect 32772 21412 32824 21418
rect 32772 21354 32824 21360
rect 32784 18970 32812 21354
rect 32864 20936 32916 20942
rect 32864 20878 32916 20884
rect 32876 20466 32904 20878
rect 32864 20460 32916 20466
rect 32864 20402 32916 20408
rect 32864 20256 32916 20262
rect 32864 20198 32916 20204
rect 32772 18964 32824 18970
rect 32772 18906 32824 18912
rect 32876 18698 32904 20198
rect 32864 18692 32916 18698
rect 32864 18634 32916 18640
rect 32772 17876 32824 17882
rect 32772 17818 32824 17824
rect 32680 17672 32732 17678
rect 32784 17649 32812 17818
rect 32680 17614 32732 17620
rect 32770 17640 32826 17649
rect 32692 17270 32720 17614
rect 32770 17575 32826 17584
rect 32680 17264 32732 17270
rect 32680 17206 32732 17212
rect 32588 17196 32640 17202
rect 32588 17138 32640 17144
rect 32600 16697 32628 17138
rect 32586 16688 32642 16697
rect 32586 16623 32642 16632
rect 32772 15904 32824 15910
rect 32772 15846 32824 15852
rect 32496 15632 32548 15638
rect 32496 15574 32548 15580
rect 32404 13524 32456 13530
rect 32404 13466 32456 13472
rect 32402 13424 32458 13433
rect 32402 13359 32458 13368
rect 32312 10668 32364 10674
rect 32312 10610 32364 10616
rect 32128 10600 32180 10606
rect 32128 10542 32180 10548
rect 32036 10056 32088 10062
rect 32036 9998 32088 10004
rect 32140 9994 32168 10542
rect 32128 9988 32180 9994
rect 32128 9930 32180 9936
rect 32126 9616 32182 9625
rect 32126 9551 32128 9560
rect 32180 9551 32182 9560
rect 32128 9522 32180 9528
rect 32416 9042 32444 13359
rect 32508 13326 32536 15574
rect 32784 15570 32812 15846
rect 32772 15564 32824 15570
rect 32772 15506 32824 15512
rect 32772 13932 32824 13938
rect 32772 13874 32824 13880
rect 32588 13728 32640 13734
rect 32588 13670 32640 13676
rect 32496 13320 32548 13326
rect 32496 13262 32548 13268
rect 32496 13184 32548 13190
rect 32496 13126 32548 13132
rect 32508 12850 32536 13126
rect 32496 12844 32548 12850
rect 32496 12786 32548 12792
rect 32600 10674 32628 13670
rect 32784 13462 32812 13874
rect 32876 13462 32904 18634
rect 32968 17678 32996 22034
rect 33048 21548 33100 21554
rect 33048 21490 33100 21496
rect 33060 21010 33088 21490
rect 33048 21004 33100 21010
rect 33048 20946 33100 20952
rect 33048 20256 33100 20262
rect 33048 20198 33100 20204
rect 33060 19854 33088 20198
rect 33048 19848 33100 19854
rect 33048 19790 33100 19796
rect 33152 18306 33180 22170
rect 33244 22166 33272 22358
rect 33506 22335 33562 22344
rect 33232 22160 33284 22166
rect 33232 22102 33284 22108
rect 33244 21690 33272 22102
rect 33612 22094 33640 23718
rect 33692 23656 33744 23662
rect 33692 23598 33744 23604
rect 33704 23186 33732 23598
rect 33692 23180 33744 23186
rect 33692 23122 33744 23128
rect 33968 23112 34020 23118
rect 33968 23054 34020 23060
rect 33692 22976 33744 22982
rect 33692 22918 33744 22924
rect 33428 22066 33640 22094
rect 33232 21684 33284 21690
rect 33232 21626 33284 21632
rect 33232 21344 33284 21350
rect 33232 21286 33284 21292
rect 33244 20398 33272 21286
rect 33232 20392 33284 20398
rect 33232 20334 33284 20340
rect 33324 19780 33376 19786
rect 33324 19722 33376 19728
rect 33336 19446 33364 19722
rect 33324 19440 33376 19446
rect 33324 19382 33376 19388
rect 33152 18278 33272 18306
rect 33140 18148 33192 18154
rect 33140 18090 33192 18096
rect 33048 17740 33100 17746
rect 33048 17682 33100 17688
rect 32956 17672 33008 17678
rect 32956 17614 33008 17620
rect 32956 17536 33008 17542
rect 32956 17478 33008 17484
rect 32968 16726 32996 17478
rect 32956 16720 33008 16726
rect 32956 16662 33008 16668
rect 33060 15706 33088 17682
rect 33048 15700 33100 15706
rect 33048 15642 33100 15648
rect 33048 15360 33100 15366
rect 33048 15302 33100 15308
rect 32956 14340 33008 14346
rect 32956 14282 33008 14288
rect 32968 14074 32996 14282
rect 32956 14068 33008 14074
rect 32956 14010 33008 14016
rect 32956 13864 33008 13870
rect 32956 13806 33008 13812
rect 32772 13456 32824 13462
rect 32772 13398 32824 13404
rect 32864 13456 32916 13462
rect 32864 13398 32916 13404
rect 32784 13326 32812 13398
rect 32772 13320 32824 13326
rect 32772 13262 32824 13268
rect 32968 12986 32996 13806
rect 33060 13258 33088 15302
rect 33152 15094 33180 18090
rect 33244 16114 33272 18278
rect 33336 17678 33364 19382
rect 33324 17672 33376 17678
rect 33324 17614 33376 17620
rect 33336 16182 33364 17614
rect 33324 16176 33376 16182
rect 33324 16118 33376 16124
rect 33232 16108 33284 16114
rect 33232 16050 33284 16056
rect 33232 15428 33284 15434
rect 33232 15370 33284 15376
rect 33140 15088 33192 15094
rect 33140 15030 33192 15036
rect 33244 13802 33272 15370
rect 33324 14884 33376 14890
rect 33324 14826 33376 14832
rect 33232 13796 33284 13802
rect 33232 13738 33284 13744
rect 33244 13462 33272 13738
rect 33232 13456 33284 13462
rect 33232 13398 33284 13404
rect 33232 13320 33284 13326
rect 33232 13262 33284 13268
rect 33048 13252 33100 13258
rect 33048 13194 33100 13200
rect 32956 12980 33008 12986
rect 32956 12922 33008 12928
rect 33244 12850 33272 13262
rect 32956 12844 33008 12850
rect 32956 12786 33008 12792
rect 33232 12844 33284 12850
rect 33232 12786 33284 12792
rect 32864 11756 32916 11762
rect 32864 11698 32916 11704
rect 32876 11150 32904 11698
rect 32864 11144 32916 11150
rect 32862 11112 32864 11121
rect 32916 11112 32918 11121
rect 32862 11047 32918 11056
rect 32680 11008 32732 11014
rect 32680 10950 32732 10956
rect 32772 11008 32824 11014
rect 32772 10950 32824 10956
rect 32588 10668 32640 10674
rect 32588 10610 32640 10616
rect 32692 10062 32720 10950
rect 32784 10266 32812 10950
rect 32864 10804 32916 10810
rect 32864 10746 32916 10752
rect 32876 10674 32904 10746
rect 32968 10674 32996 12786
rect 33232 12232 33284 12238
rect 33232 12174 33284 12180
rect 33048 11892 33100 11898
rect 33048 11834 33100 11840
rect 33060 11218 33088 11834
rect 33048 11212 33100 11218
rect 33048 11154 33100 11160
rect 32864 10668 32916 10674
rect 32864 10610 32916 10616
rect 32956 10668 33008 10674
rect 32956 10610 33008 10616
rect 32772 10260 32824 10266
rect 32772 10202 32824 10208
rect 32680 10056 32732 10062
rect 32680 9998 32732 10004
rect 32968 9994 32996 10610
rect 33060 10062 33088 11154
rect 33244 11064 33272 12174
rect 33336 11218 33364 14826
rect 33428 11558 33456 22066
rect 33508 20800 33560 20806
rect 33508 20742 33560 20748
rect 33520 17814 33548 20742
rect 33600 20460 33652 20466
rect 33600 20402 33652 20408
rect 33612 18358 33640 20402
rect 33704 19990 33732 22918
rect 33876 22636 33928 22642
rect 33876 22578 33928 22584
rect 33784 21684 33836 21690
rect 33784 21626 33836 21632
rect 33796 20942 33824 21626
rect 33784 20936 33836 20942
rect 33784 20878 33836 20884
rect 33888 20874 33916 22578
rect 33980 21894 34008 23054
rect 34072 22234 34100 26794
rect 34164 24886 34192 28376
rect 34244 28358 34296 28364
rect 34428 27532 34480 27538
rect 34428 27474 34480 27480
rect 34440 26994 34468 27474
rect 34428 26988 34480 26994
rect 34428 26930 34480 26936
rect 34440 26790 34468 26930
rect 34428 26784 34480 26790
rect 34428 26726 34480 26732
rect 34532 26586 34560 29174
rect 34610 29135 34612 29144
rect 34664 29135 34666 29144
rect 34612 29106 34664 29112
rect 34808 29050 34836 31078
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35452 30274 35480 31214
rect 36372 30938 36400 31282
rect 36360 30932 36412 30938
rect 36360 30874 36412 30880
rect 36084 30864 36136 30870
rect 36084 30806 36136 30812
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 35452 30246 35756 30274
rect 35348 30048 35400 30054
rect 35348 29990 35400 29996
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35256 29844 35308 29850
rect 35360 29832 35388 29990
rect 35308 29804 35388 29832
rect 35256 29786 35308 29792
rect 34888 29776 34940 29782
rect 34888 29718 34940 29724
rect 35164 29776 35216 29782
rect 35164 29718 35216 29724
rect 34624 29022 34836 29050
rect 34520 26580 34572 26586
rect 34520 26522 34572 26528
rect 34428 26376 34480 26382
rect 34428 26318 34480 26324
rect 34440 25906 34468 26318
rect 34532 25906 34560 26522
rect 34336 25900 34388 25906
rect 34336 25842 34388 25848
rect 34428 25900 34480 25906
rect 34428 25842 34480 25848
rect 34520 25900 34572 25906
rect 34520 25842 34572 25848
rect 34348 25362 34376 25842
rect 34428 25764 34480 25770
rect 34428 25706 34480 25712
rect 34336 25356 34388 25362
rect 34256 25316 34336 25344
rect 34152 24880 34204 24886
rect 34152 24822 34204 24828
rect 34164 23594 34192 24822
rect 34152 23588 34204 23594
rect 34152 23530 34204 23536
rect 34164 23322 34192 23530
rect 34152 23316 34204 23322
rect 34152 23258 34204 23264
rect 34256 23050 34284 25316
rect 34336 25298 34388 25304
rect 34336 23724 34388 23730
rect 34336 23666 34388 23672
rect 34244 23044 34296 23050
rect 34244 22986 34296 22992
rect 34060 22228 34112 22234
rect 34060 22170 34112 22176
rect 33968 21888 34020 21894
rect 33968 21830 34020 21836
rect 34152 21684 34204 21690
rect 34152 21626 34204 21632
rect 33968 21480 34020 21486
rect 33968 21422 34020 21428
rect 33876 20868 33928 20874
rect 33876 20810 33928 20816
rect 33784 20392 33836 20398
rect 33784 20334 33836 20340
rect 33692 19984 33744 19990
rect 33692 19926 33744 19932
rect 33692 19712 33744 19718
rect 33692 19654 33744 19660
rect 33600 18352 33652 18358
rect 33600 18294 33652 18300
rect 33508 17808 33560 17814
rect 33508 17750 33560 17756
rect 33508 17604 33560 17610
rect 33508 17546 33560 17552
rect 33600 17604 33652 17610
rect 33600 17546 33652 17552
rect 33520 17338 33548 17546
rect 33508 17332 33560 17338
rect 33508 17274 33560 17280
rect 33520 12782 33548 17274
rect 33612 17202 33640 17546
rect 33600 17196 33652 17202
rect 33600 17138 33652 17144
rect 33598 17096 33654 17105
rect 33598 17031 33600 17040
rect 33652 17031 33654 17040
rect 33600 17002 33652 17008
rect 33600 16516 33652 16522
rect 33600 16458 33652 16464
rect 33612 14482 33640 16458
rect 33600 14476 33652 14482
rect 33600 14418 33652 14424
rect 33600 13864 33652 13870
rect 33600 13806 33652 13812
rect 33508 12776 33560 12782
rect 33508 12718 33560 12724
rect 33508 12300 33560 12306
rect 33508 12242 33560 12248
rect 33520 12209 33548 12242
rect 33506 12200 33562 12209
rect 33506 12135 33562 12144
rect 33520 11830 33548 12135
rect 33612 11898 33640 13806
rect 33704 12889 33732 19654
rect 33796 19530 33824 20334
rect 33888 19922 33916 20810
rect 33980 20602 34008 21422
rect 33968 20596 34020 20602
rect 33968 20538 34020 20544
rect 33968 20256 34020 20262
rect 33968 20198 34020 20204
rect 33876 19916 33928 19922
rect 33876 19858 33928 19864
rect 33888 19718 33916 19858
rect 33876 19712 33928 19718
rect 33876 19654 33928 19660
rect 33796 19502 33916 19530
rect 33784 18284 33836 18290
rect 33784 18226 33836 18232
rect 33796 17678 33824 18226
rect 33784 17672 33836 17678
rect 33784 17614 33836 17620
rect 33888 16232 33916 19502
rect 33980 19446 34008 20198
rect 34164 19446 34192 21626
rect 33968 19440 34020 19446
rect 33968 19382 34020 19388
rect 34152 19440 34204 19446
rect 34152 19382 34204 19388
rect 34256 19378 34284 22986
rect 34060 19372 34112 19378
rect 34060 19314 34112 19320
rect 34244 19372 34296 19378
rect 34244 19314 34296 19320
rect 34072 19242 34100 19314
rect 34060 19236 34112 19242
rect 34060 19178 34112 19184
rect 33968 19168 34020 19174
rect 33968 19110 34020 19116
rect 33796 16204 33916 16232
rect 33796 15910 33824 16204
rect 33876 16108 33928 16114
rect 33876 16050 33928 16056
rect 33784 15904 33836 15910
rect 33784 15846 33836 15852
rect 33690 12880 33746 12889
rect 33690 12815 33746 12824
rect 33796 12442 33824 15846
rect 33888 15366 33916 16050
rect 33876 15360 33928 15366
rect 33876 15302 33928 15308
rect 33980 15162 34008 19110
rect 34060 18148 34112 18154
rect 34060 18090 34112 18096
rect 34072 17882 34100 18090
rect 34060 17876 34112 17882
rect 34060 17818 34112 17824
rect 34348 17762 34376 23666
rect 34440 22710 34468 25706
rect 34520 23860 34572 23866
rect 34520 23802 34572 23808
rect 34532 23254 34560 23802
rect 34520 23248 34572 23254
rect 34520 23190 34572 23196
rect 34428 22704 34480 22710
rect 34428 22646 34480 22652
rect 34440 22094 34468 22646
rect 34440 22066 34560 22094
rect 34428 21888 34480 21894
rect 34428 21830 34480 21836
rect 34440 21418 34468 21830
rect 34428 21412 34480 21418
rect 34428 21354 34480 21360
rect 34440 20942 34468 21354
rect 34428 20936 34480 20942
rect 34428 20878 34480 20884
rect 34440 20330 34468 20878
rect 34428 20324 34480 20330
rect 34428 20266 34480 20272
rect 34428 19984 34480 19990
rect 34428 19926 34480 19932
rect 34440 19242 34468 19926
rect 34428 19236 34480 19242
rect 34428 19178 34480 19184
rect 34440 18834 34468 19178
rect 34428 18828 34480 18834
rect 34428 18770 34480 18776
rect 34532 18748 34560 22066
rect 34624 21690 34652 29022
rect 34900 28948 34928 29718
rect 35072 29572 35124 29578
rect 35072 29514 35124 29520
rect 35084 29481 35112 29514
rect 35070 29472 35126 29481
rect 35070 29407 35126 29416
rect 34978 29336 35034 29345
rect 34978 29271 35034 29280
rect 35072 29300 35124 29306
rect 34992 29170 35020 29271
rect 35176 29288 35204 29718
rect 35124 29260 35204 29288
rect 35072 29242 35124 29248
rect 34980 29164 35032 29170
rect 34980 29106 35032 29112
rect 35268 29034 35296 29786
rect 35440 29640 35492 29646
rect 35440 29582 35492 29588
rect 35622 29608 35678 29617
rect 35452 29220 35480 29582
rect 35728 29594 35756 30246
rect 36096 30054 36124 30806
rect 36268 30796 36320 30802
rect 36268 30738 36320 30744
rect 36176 30728 36228 30734
rect 36176 30670 36228 30676
rect 36188 30598 36216 30670
rect 36176 30592 36228 30598
rect 36176 30534 36228 30540
rect 36188 30190 36216 30534
rect 36280 30258 36308 30738
rect 36372 30569 36400 30874
rect 36358 30560 36414 30569
rect 36358 30495 36414 30504
rect 36360 30388 36412 30394
rect 36360 30330 36412 30336
rect 36268 30252 36320 30258
rect 36268 30194 36320 30200
rect 36176 30184 36228 30190
rect 36176 30126 36228 30132
rect 36084 30048 36136 30054
rect 36084 29990 36136 29996
rect 36096 29782 36124 29990
rect 36084 29776 36136 29782
rect 36084 29718 36136 29724
rect 36188 29714 36216 30126
rect 36372 30054 36400 30330
rect 36360 30048 36412 30054
rect 36360 29990 36412 29996
rect 36464 29850 36492 31282
rect 36556 30394 36584 31690
rect 37188 31408 37240 31414
rect 37240 31356 37320 31362
rect 37188 31350 37320 31356
rect 37200 31334 37320 31350
rect 37384 31346 37412 32234
rect 37292 31142 37320 31334
rect 37372 31340 37424 31346
rect 37372 31282 37424 31288
rect 37476 31210 37504 32302
rect 37568 31754 37596 32302
rect 37568 31726 37688 31754
rect 37660 31362 37688 31726
rect 37844 31634 37872 32302
rect 38016 32224 38068 32230
rect 38016 32166 38068 32172
rect 38028 32026 38056 32166
rect 38016 32020 38068 32026
rect 38016 31962 38068 31968
rect 38212 31822 38240 32370
rect 38660 31952 38712 31958
rect 38660 31894 38712 31900
rect 38672 31822 38700 31894
rect 38200 31816 38252 31822
rect 38200 31758 38252 31764
rect 38292 31816 38344 31822
rect 38292 31758 38344 31764
rect 38568 31816 38620 31822
rect 38568 31758 38620 31764
rect 38660 31816 38712 31822
rect 38660 31758 38712 31764
rect 37752 31606 37872 31634
rect 37752 31482 37780 31606
rect 37740 31476 37792 31482
rect 37740 31418 37792 31424
rect 37832 31476 37884 31482
rect 37832 31418 37884 31424
rect 37844 31362 37872 31418
rect 37660 31334 37872 31362
rect 38212 31346 38240 31758
rect 37556 31272 37608 31278
rect 37608 31232 37688 31260
rect 37556 31214 37608 31220
rect 37464 31204 37516 31210
rect 37464 31146 37516 31152
rect 37280 31136 37332 31142
rect 37280 31078 37332 31084
rect 37476 30938 37504 31146
rect 37464 30932 37516 30938
rect 37464 30874 37516 30880
rect 36820 30864 36872 30870
rect 36820 30806 36872 30812
rect 37004 30864 37056 30870
rect 37004 30806 37056 30812
rect 36832 30734 36860 30806
rect 36820 30728 36872 30734
rect 36820 30670 36872 30676
rect 36728 30592 36780 30598
rect 36728 30534 36780 30540
rect 36544 30388 36596 30394
rect 36544 30330 36596 30336
rect 36542 30152 36598 30161
rect 36542 30087 36598 30096
rect 36452 29844 36504 29850
rect 36452 29786 36504 29792
rect 36176 29708 36228 29714
rect 36176 29650 36228 29656
rect 35728 29566 36124 29594
rect 35622 29543 35624 29552
rect 35676 29543 35678 29552
rect 35624 29514 35676 29520
rect 35992 29504 36044 29510
rect 36096 29492 36124 29566
rect 36176 29504 36228 29510
rect 36096 29464 36176 29492
rect 35992 29446 36044 29452
rect 36176 29446 36228 29452
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 36004 29288 36032 29446
rect 36084 29300 36136 29306
rect 36004 29260 36084 29288
rect 35532 29232 35584 29238
rect 35452 29192 35532 29220
rect 35532 29174 35584 29180
rect 35714 29200 35770 29209
rect 35256 29028 35308 29034
rect 35256 28970 35308 28976
rect 34702 28928 34758 28937
rect 34702 28863 34758 28872
rect 34808 28920 34928 28948
rect 34716 26217 34744 28863
rect 34702 26208 34758 26217
rect 34702 26143 34758 26152
rect 34704 25696 34756 25702
rect 34704 25638 34756 25644
rect 34612 21684 34664 21690
rect 34612 21626 34664 21632
rect 34612 21548 34664 21554
rect 34716 21536 34744 25638
rect 34808 25226 34836 28920
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35440 28620 35492 28626
rect 35440 28562 35492 28568
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35348 26784 35400 26790
rect 35348 26726 35400 26732
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35360 26518 35388 26726
rect 35348 26512 35400 26518
rect 35348 26454 35400 26460
rect 34888 26240 34940 26246
rect 34888 26182 34940 26188
rect 35072 26240 35124 26246
rect 35072 26182 35124 26188
rect 35162 26208 35218 26217
rect 34900 25906 34928 26182
rect 35084 25906 35112 26182
rect 35162 26143 35218 26152
rect 34888 25900 34940 25906
rect 34888 25842 34940 25848
rect 35072 25900 35124 25906
rect 35072 25842 35124 25848
rect 35176 25838 35204 26143
rect 35348 25968 35400 25974
rect 35348 25910 35400 25916
rect 35164 25832 35216 25838
rect 35164 25774 35216 25780
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35360 25514 35388 25910
rect 35268 25486 35388 25514
rect 34796 25220 34848 25226
rect 34796 25162 34848 25168
rect 35268 24818 35296 25486
rect 35348 25152 35400 25158
rect 35348 25094 35400 25100
rect 35360 24818 35388 25094
rect 35256 24812 35308 24818
rect 35256 24754 35308 24760
rect 35348 24812 35400 24818
rect 35348 24754 35400 24760
rect 35268 24721 35296 24754
rect 35254 24712 35310 24721
rect 35254 24647 35310 24656
rect 35348 24676 35400 24682
rect 35348 24618 35400 24624
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35360 24070 35388 24618
rect 35348 24064 35400 24070
rect 35348 24006 35400 24012
rect 34886 23760 34942 23769
rect 34886 23695 34888 23704
rect 34940 23695 34942 23704
rect 34888 23666 34940 23672
rect 34796 23656 34848 23662
rect 34794 23624 34796 23633
rect 34848 23624 34850 23633
rect 34794 23559 34850 23568
rect 34796 23520 34848 23526
rect 34796 23462 34848 23468
rect 34808 22574 34836 23462
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35254 22808 35310 22817
rect 35254 22743 35310 22752
rect 34796 22568 34848 22574
rect 34796 22510 34848 22516
rect 34808 22216 34836 22510
rect 35268 22386 35296 22743
rect 35268 22358 35301 22386
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35273 22250 35301 22358
rect 35268 22222 35301 22250
rect 34808 22188 34928 22216
rect 34796 21684 34848 21690
rect 34796 21626 34848 21632
rect 34664 21508 34744 21536
rect 34612 21490 34664 21496
rect 34808 21434 34836 21626
rect 34900 21554 34928 22188
rect 35268 21622 35296 22222
rect 35256 21616 35308 21622
rect 35256 21558 35308 21564
rect 34888 21548 34940 21554
rect 34888 21490 34940 21496
rect 34716 21406 34836 21434
rect 34610 20768 34666 20777
rect 34610 20703 34666 20712
rect 34624 19446 34652 20703
rect 34716 20466 34744 21406
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34796 21072 34848 21078
rect 34796 21014 34848 21020
rect 34704 20460 34756 20466
rect 34704 20402 34756 20408
rect 34808 19514 34836 21014
rect 35256 20800 35308 20806
rect 35256 20742 35308 20748
rect 35268 20262 35296 20742
rect 35256 20256 35308 20262
rect 35256 20198 35308 20204
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35360 20074 35388 24006
rect 35452 22642 35480 28562
rect 35544 28558 35572 29174
rect 35714 29135 35770 29144
rect 35728 28994 35756 29135
rect 35636 28966 35756 28994
rect 35808 29028 35860 29034
rect 35808 28970 35860 28976
rect 35532 28552 35584 28558
rect 35532 28494 35584 28500
rect 35636 28422 35664 28966
rect 35820 28626 35848 28970
rect 35808 28620 35860 28626
rect 35808 28562 35860 28568
rect 36004 28558 36032 29260
rect 36084 29242 36136 29248
rect 36082 29200 36138 29209
rect 36082 29135 36084 29144
rect 36136 29135 36138 29144
rect 36084 29106 36136 29112
rect 35992 28552 36044 28558
rect 35992 28494 36044 28500
rect 36188 28490 36216 29446
rect 36464 29238 36492 29786
rect 36556 29782 36584 30087
rect 36544 29776 36596 29782
rect 36544 29718 36596 29724
rect 36634 29744 36690 29753
rect 36634 29679 36636 29688
rect 36688 29679 36690 29688
rect 36636 29650 36688 29656
rect 36740 29238 36768 30534
rect 36832 30258 36860 30670
rect 36820 30252 36872 30258
rect 36820 30194 36872 30200
rect 36818 29880 36874 29889
rect 36818 29815 36874 29824
rect 36832 29646 36860 29815
rect 36820 29640 36872 29646
rect 36820 29582 36872 29588
rect 36910 29608 36966 29617
rect 36910 29543 36966 29552
rect 36924 29238 36952 29543
rect 36452 29232 36504 29238
rect 36452 29174 36504 29180
rect 36728 29232 36780 29238
rect 36728 29174 36780 29180
rect 36912 29232 36964 29238
rect 36912 29174 36964 29180
rect 36268 29164 36320 29170
rect 36268 29106 36320 29112
rect 36544 29164 36596 29170
rect 36544 29106 36596 29112
rect 36280 29034 36308 29106
rect 36556 29050 36584 29106
rect 36268 29028 36320 29034
rect 36556 29022 36676 29050
rect 36268 28970 36320 28976
rect 36176 28484 36228 28490
rect 36176 28426 36228 28432
rect 35624 28416 35676 28422
rect 35624 28358 35676 28364
rect 36084 28416 36136 28422
rect 36084 28358 36136 28364
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 36096 27674 36124 28358
rect 36084 27668 36136 27674
rect 36084 27610 36136 27616
rect 35992 27328 36044 27334
rect 35992 27270 36044 27276
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35594 27163 35902 27172
rect 35622 26888 35678 26897
rect 35532 26852 35584 26858
rect 35622 26823 35678 26832
rect 35532 26794 35584 26800
rect 35544 26382 35572 26794
rect 35532 26376 35584 26382
rect 35532 26318 35584 26324
rect 35636 26314 35664 26823
rect 36004 26314 36032 27270
rect 35624 26308 35676 26314
rect 35624 26250 35676 26256
rect 35992 26308 36044 26314
rect 35992 26250 36044 26256
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 36096 26042 36124 27610
rect 36084 26036 36136 26042
rect 36084 25978 36136 25984
rect 36176 25968 36228 25974
rect 36176 25910 36228 25916
rect 35992 25832 36044 25838
rect 35992 25774 36044 25780
rect 35808 25696 35860 25702
rect 35808 25638 35860 25644
rect 35820 25498 35848 25638
rect 35808 25492 35860 25498
rect 35808 25434 35860 25440
rect 35532 25288 35584 25294
rect 35530 25256 35532 25265
rect 35584 25256 35586 25265
rect 36004 25226 36032 25774
rect 36084 25288 36136 25294
rect 36084 25230 36136 25236
rect 35530 25191 35586 25200
rect 35992 25220 36044 25226
rect 35992 25162 36044 25168
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 35594 23964 35902 23973
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 36004 23848 36032 25162
rect 36096 24410 36124 25230
rect 36188 25158 36216 25910
rect 36176 25152 36228 25158
rect 36176 25094 36228 25100
rect 36084 24404 36136 24410
rect 36084 24346 36136 24352
rect 35912 23820 36032 23848
rect 35912 22982 35940 23820
rect 35992 23044 36044 23050
rect 35992 22986 36044 22992
rect 35900 22976 35952 22982
rect 35900 22918 35952 22924
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 35440 22636 35492 22642
rect 35440 22578 35492 22584
rect 35594 21788 35902 21797
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 36004 21554 36032 22986
rect 36280 22778 36308 28970
rect 36452 28756 36504 28762
rect 36452 28698 36504 28704
rect 36360 26920 36412 26926
rect 36360 26862 36412 26868
rect 36372 26586 36400 26862
rect 36360 26580 36412 26586
rect 36360 26522 36412 26528
rect 36360 25696 36412 25702
rect 36360 25638 36412 25644
rect 36372 25294 36400 25638
rect 36360 25288 36412 25294
rect 36360 25230 36412 25236
rect 36464 25158 36492 28698
rect 36544 27328 36596 27334
rect 36544 27270 36596 27276
rect 36556 27130 36584 27270
rect 36544 27124 36596 27130
rect 36544 27066 36596 27072
rect 36544 26240 36596 26246
rect 36544 26182 36596 26188
rect 36452 25152 36504 25158
rect 36452 25094 36504 25100
rect 36556 24206 36584 26182
rect 36648 24936 36676 29022
rect 36740 25974 36768 29174
rect 37016 27946 37044 30806
rect 37556 30796 37608 30802
rect 37556 30738 37608 30744
rect 37372 30728 37424 30734
rect 37372 30670 37424 30676
rect 37384 30258 37412 30670
rect 37464 30660 37516 30666
rect 37464 30602 37516 30608
rect 37372 30252 37424 30258
rect 37372 30194 37424 30200
rect 37280 30048 37332 30054
rect 37280 29990 37332 29996
rect 37372 30048 37424 30054
rect 37476 30036 37504 30602
rect 37568 30258 37596 30738
rect 37660 30734 37688 31232
rect 37648 30728 37700 30734
rect 37648 30670 37700 30676
rect 37648 30592 37700 30598
rect 37648 30534 37700 30540
rect 37556 30252 37608 30258
rect 37556 30194 37608 30200
rect 37424 30008 37504 30036
rect 37372 29990 37424 29996
rect 37292 29170 37320 29990
rect 37384 29578 37412 29990
rect 37660 29646 37688 30534
rect 37844 30410 37872 31334
rect 38200 31340 38252 31346
rect 38200 31282 38252 31288
rect 38108 30660 38160 30666
rect 38108 30602 38160 30608
rect 37752 30382 37872 30410
rect 37924 30388 37976 30394
rect 37464 29640 37516 29646
rect 37464 29582 37516 29588
rect 37648 29640 37700 29646
rect 37648 29582 37700 29588
rect 37372 29572 37424 29578
rect 37372 29514 37424 29520
rect 37280 29164 37332 29170
rect 37280 29106 37332 29112
rect 37004 27940 37056 27946
rect 37004 27882 37056 27888
rect 36820 27464 36872 27470
rect 36820 27406 36872 27412
rect 36832 26994 36860 27406
rect 36912 27328 36964 27334
rect 36912 27270 36964 27276
rect 36820 26988 36872 26994
rect 36820 26930 36872 26936
rect 36728 25968 36780 25974
rect 36728 25910 36780 25916
rect 36818 25392 36874 25401
rect 36818 25327 36820 25336
rect 36872 25327 36874 25336
rect 36820 25298 36872 25304
rect 36728 24948 36780 24954
rect 36648 24908 36728 24936
rect 36728 24890 36780 24896
rect 36636 24744 36688 24750
rect 36636 24686 36688 24692
rect 36544 24200 36596 24206
rect 36544 24142 36596 24148
rect 36360 23792 36412 23798
rect 36360 23734 36412 23740
rect 36268 22772 36320 22778
rect 36268 22714 36320 22720
rect 36174 22672 36230 22681
rect 36174 22607 36176 22616
rect 36228 22607 36230 22616
rect 36176 22578 36228 22584
rect 36280 21622 36308 22714
rect 36268 21616 36320 21622
rect 36268 21558 36320 21564
rect 35716 21548 35768 21554
rect 35716 21490 35768 21496
rect 35900 21548 35952 21554
rect 35900 21490 35952 21496
rect 35992 21548 36044 21554
rect 35992 21490 36044 21496
rect 35728 21078 35756 21490
rect 35716 21072 35768 21078
rect 35716 21014 35768 21020
rect 35912 20806 35940 21490
rect 35992 21344 36044 21350
rect 36176 21344 36228 21350
rect 36044 21304 36124 21332
rect 35992 21286 36044 21292
rect 36096 21078 36124 21304
rect 36176 21286 36228 21292
rect 36084 21072 36136 21078
rect 36084 21014 36136 21020
rect 35900 20800 35952 20806
rect 35900 20742 35952 20748
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 35992 20324 36044 20330
rect 35992 20266 36044 20272
rect 35360 20046 35480 20074
rect 35164 19916 35216 19922
rect 35164 19858 35216 19864
rect 35348 19916 35400 19922
rect 35348 19858 35400 19864
rect 34796 19508 34848 19514
rect 34796 19450 34848 19456
rect 34612 19440 34664 19446
rect 34612 19382 34664 19388
rect 34702 19408 34758 19417
rect 34624 18902 34652 19382
rect 34808 19394 34836 19450
rect 34808 19366 34928 19394
rect 35176 19378 35204 19858
rect 34702 19343 34758 19352
rect 34716 19156 34744 19343
rect 34900 19310 34928 19366
rect 34980 19372 35032 19378
rect 34980 19314 35032 19320
rect 35164 19372 35216 19378
rect 35164 19314 35216 19320
rect 34888 19304 34940 19310
rect 34888 19246 34940 19252
rect 34992 19156 35020 19314
rect 34716 19128 35020 19156
rect 34612 18896 34664 18902
rect 34612 18838 34664 18844
rect 34704 18760 34756 18766
rect 34532 18720 34704 18748
rect 34704 18702 34756 18708
rect 34612 18624 34664 18630
rect 34612 18566 34664 18572
rect 34428 18352 34480 18358
rect 34426 18320 34428 18329
rect 34480 18320 34482 18329
rect 34426 18255 34482 18264
rect 34520 18216 34572 18222
rect 34520 18158 34572 18164
rect 34072 17734 34376 17762
rect 34072 16522 34100 17734
rect 34152 17672 34204 17678
rect 34428 17672 34480 17678
rect 34152 17614 34204 17620
rect 34256 17632 34428 17660
rect 34164 17542 34192 17614
rect 34152 17536 34204 17542
rect 34152 17478 34204 17484
rect 34060 16516 34112 16522
rect 34060 16458 34112 16464
rect 34060 16176 34112 16182
rect 34060 16118 34112 16124
rect 33968 15156 34020 15162
rect 33968 15098 34020 15104
rect 33980 15026 34008 15098
rect 33968 15020 34020 15026
rect 33968 14962 34020 14968
rect 34072 14822 34100 16118
rect 34060 14816 34112 14822
rect 34060 14758 34112 14764
rect 34164 13530 34192 17478
rect 34256 16182 34284 17632
rect 34428 17614 34480 17620
rect 34428 17536 34480 17542
rect 34428 17478 34480 17484
rect 34440 17270 34468 17478
rect 34428 17264 34480 17270
rect 34428 17206 34480 17212
rect 34244 16176 34296 16182
rect 34428 16176 34480 16182
rect 34244 16118 34296 16124
rect 34426 16144 34428 16153
rect 34480 16144 34482 16153
rect 34532 16114 34560 18158
rect 34426 16079 34482 16088
rect 34520 16108 34572 16114
rect 34520 16050 34572 16056
rect 34244 16040 34296 16046
rect 34244 15982 34296 15988
rect 34152 13524 34204 13530
rect 34152 13466 34204 13472
rect 33968 13252 34020 13258
rect 33968 13194 34020 13200
rect 33784 12436 33836 12442
rect 33784 12378 33836 12384
rect 33876 12368 33928 12374
rect 33876 12310 33928 12316
rect 33600 11892 33652 11898
rect 33600 11834 33652 11840
rect 33508 11824 33560 11830
rect 33508 11766 33560 11772
rect 33598 11792 33654 11801
rect 33598 11727 33600 11736
rect 33652 11727 33654 11736
rect 33600 11698 33652 11704
rect 33508 11688 33560 11694
rect 33508 11630 33560 11636
rect 33416 11552 33468 11558
rect 33416 11494 33468 11500
rect 33324 11212 33376 11218
rect 33324 11154 33376 11160
rect 33416 11144 33468 11150
rect 33416 11086 33468 11092
rect 33324 11076 33376 11082
rect 33244 11036 33324 11064
rect 33324 11018 33376 11024
rect 33232 10600 33284 10606
rect 33232 10542 33284 10548
rect 33048 10056 33100 10062
rect 33048 9998 33100 10004
rect 32956 9988 33008 9994
rect 32956 9930 33008 9936
rect 32588 9580 32640 9586
rect 32588 9522 32640 9528
rect 32680 9580 32732 9586
rect 32680 9522 32732 9528
rect 32864 9580 32916 9586
rect 32864 9522 32916 9528
rect 32404 9036 32456 9042
rect 32404 8978 32456 8984
rect 32600 8974 32628 9522
rect 32588 8968 32640 8974
rect 32588 8910 32640 8916
rect 32600 8498 32628 8910
rect 32692 8838 32720 9522
rect 32876 8974 32904 9522
rect 32864 8968 32916 8974
rect 32864 8910 32916 8916
rect 32680 8832 32732 8838
rect 32680 8774 32732 8780
rect 31760 8492 31812 8498
rect 31760 8434 31812 8440
rect 32588 8492 32640 8498
rect 32588 8434 32640 8440
rect 33048 8424 33100 8430
rect 33244 8378 33272 10542
rect 33336 9586 33364 11018
rect 33428 10266 33456 11086
rect 33416 10260 33468 10266
rect 33416 10202 33468 10208
rect 33324 9580 33376 9586
rect 33324 9522 33376 9528
rect 33416 9036 33468 9042
rect 33416 8978 33468 8984
rect 33324 8900 33376 8906
rect 33324 8842 33376 8848
rect 33100 8372 33272 8378
rect 33048 8366 33272 8372
rect 33060 8350 33272 8366
rect 32312 8288 32364 8294
rect 32312 8230 32364 8236
rect 32324 7954 32352 8230
rect 33060 7954 33088 8350
rect 32312 7948 32364 7954
rect 33048 7948 33100 7954
rect 32364 7908 32444 7936
rect 32312 7890 32364 7896
rect 32312 7744 32364 7750
rect 32312 7686 32364 7692
rect 32324 7342 32352 7686
rect 32416 7410 32444 7908
rect 33048 7890 33100 7896
rect 33336 7818 33364 8842
rect 33428 7954 33456 8978
rect 33520 8072 33548 11630
rect 33600 11212 33652 11218
rect 33600 11154 33652 11160
rect 33612 11121 33640 11154
rect 33888 11150 33916 12310
rect 33980 12238 34008 13194
rect 33968 12232 34020 12238
rect 33968 12174 34020 12180
rect 34060 11756 34112 11762
rect 34060 11698 34112 11704
rect 33968 11280 34020 11286
rect 33968 11222 34020 11228
rect 33876 11144 33928 11150
rect 33598 11112 33654 11121
rect 33876 11086 33928 11092
rect 33980 11082 34008 11222
rect 33598 11047 33654 11056
rect 33968 11076 34020 11082
rect 33968 11018 34020 11024
rect 33980 10742 34008 11018
rect 33968 10736 34020 10742
rect 33968 10678 34020 10684
rect 34072 10538 34100 11698
rect 34060 10532 34112 10538
rect 34060 10474 34112 10480
rect 33784 9988 33836 9994
rect 33784 9930 33836 9936
rect 33600 9512 33652 9518
rect 33600 9454 33652 9460
rect 33612 8906 33640 9454
rect 33692 9172 33744 9178
rect 33692 9114 33744 9120
rect 33600 8900 33652 8906
rect 33600 8842 33652 8848
rect 33704 8362 33732 9114
rect 33796 8634 33824 9930
rect 34164 9586 34192 13466
rect 34256 12102 34284 15982
rect 34336 15700 34388 15706
rect 34336 15642 34388 15648
rect 34244 12096 34296 12102
rect 34244 12038 34296 12044
rect 34256 9636 34284 12038
rect 34348 11801 34376 15642
rect 34520 15564 34572 15570
rect 34520 15506 34572 15512
rect 34428 14816 34480 14822
rect 34428 14758 34480 14764
rect 34334 11792 34390 11801
rect 34334 11727 34390 11736
rect 34336 11144 34388 11150
rect 34336 11086 34388 11092
rect 34348 10742 34376 11086
rect 34336 10736 34388 10742
rect 34336 10678 34388 10684
rect 34440 9722 34468 14758
rect 34532 12170 34560 15506
rect 34624 14958 34652 18566
rect 34716 15706 34744 18702
rect 34808 17320 34836 19128
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35360 18766 35388 19858
rect 35452 19378 35480 20046
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 35532 19508 35584 19514
rect 35532 19450 35584 19456
rect 35808 19508 35860 19514
rect 35808 19450 35860 19456
rect 35544 19417 35572 19450
rect 35530 19408 35586 19417
rect 35440 19372 35492 19378
rect 35820 19378 35848 19450
rect 35530 19343 35586 19352
rect 35808 19372 35860 19378
rect 35440 19314 35492 19320
rect 35348 18760 35400 18766
rect 35348 18702 35400 18708
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35360 17898 35388 18702
rect 35452 18290 35480 19314
rect 35544 18970 35572 19343
rect 35808 19314 35860 19320
rect 35898 19272 35954 19281
rect 35898 19207 35954 19216
rect 35912 19174 35940 19207
rect 35808 19168 35860 19174
rect 35808 19110 35860 19116
rect 35900 19168 35952 19174
rect 35900 19110 35952 19116
rect 35820 18986 35848 19110
rect 36004 18986 36032 20266
rect 35532 18964 35584 18970
rect 35532 18906 35584 18912
rect 35820 18958 36032 18986
rect 35820 18766 35848 18958
rect 35992 18896 36044 18902
rect 35898 18864 35954 18873
rect 35992 18838 36044 18844
rect 35898 18799 35954 18808
rect 35912 18766 35940 18799
rect 35808 18760 35860 18766
rect 35808 18702 35860 18708
rect 35900 18760 35952 18766
rect 35900 18702 35952 18708
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 35440 18284 35492 18290
rect 35440 18226 35492 18232
rect 35268 17870 35388 17898
rect 34886 17640 34942 17649
rect 34886 17575 34942 17584
rect 34900 17542 34928 17575
rect 34888 17536 34940 17542
rect 34888 17478 34940 17484
rect 34808 17292 34928 17320
rect 34796 17196 34848 17202
rect 34796 17138 34848 17144
rect 34808 16046 34836 17138
rect 34900 16980 34928 17292
rect 35268 17202 35296 17870
rect 35346 17504 35402 17513
rect 35346 17439 35402 17448
rect 35360 17202 35388 17439
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35594 17371 35902 17380
rect 36004 17202 36032 18838
rect 36096 17678 36124 21014
rect 36188 21010 36216 21286
rect 36176 21004 36228 21010
rect 36176 20946 36228 20952
rect 36372 20942 36400 23734
rect 36556 23118 36584 24142
rect 36452 23112 36504 23118
rect 36450 23080 36452 23089
rect 36544 23112 36596 23118
rect 36504 23080 36506 23089
rect 36544 23054 36596 23060
rect 36450 23015 36506 23024
rect 36556 22642 36584 23054
rect 36544 22636 36596 22642
rect 36544 22578 36596 22584
rect 36556 21962 36584 22578
rect 36544 21956 36596 21962
rect 36544 21898 36596 21904
rect 36556 21554 36584 21898
rect 36452 21548 36504 21554
rect 36452 21490 36504 21496
rect 36544 21548 36596 21554
rect 36544 21490 36596 21496
rect 36464 21146 36492 21490
rect 36452 21140 36504 21146
rect 36452 21082 36504 21088
rect 36360 20936 36412 20942
rect 36360 20878 36412 20884
rect 36268 20868 36320 20874
rect 36268 20810 36320 20816
rect 36176 19780 36228 19786
rect 36176 19722 36228 19728
rect 36188 19378 36216 19722
rect 36176 19372 36228 19378
rect 36176 19314 36228 19320
rect 36176 19236 36228 19242
rect 36176 19178 36228 19184
rect 36188 18630 36216 19178
rect 36176 18624 36228 18630
rect 36176 18566 36228 18572
rect 36188 18222 36216 18566
rect 36176 18216 36228 18222
rect 36176 18158 36228 18164
rect 36084 17672 36136 17678
rect 36084 17614 36136 17620
rect 36176 17672 36228 17678
rect 36176 17614 36228 17620
rect 35256 17196 35308 17202
rect 35256 17138 35308 17144
rect 35348 17196 35400 17202
rect 35348 17138 35400 17144
rect 35992 17196 36044 17202
rect 35992 17138 36044 17144
rect 35348 17060 35400 17066
rect 35348 17002 35400 17008
rect 34900 16952 35296 16980
rect 35268 16946 35296 16952
rect 35268 16918 35301 16946
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35273 16810 35301 16918
rect 35268 16782 35301 16810
rect 35360 16794 35388 17002
rect 35440 16992 35492 16998
rect 35440 16934 35492 16940
rect 35348 16788 35400 16794
rect 34980 16448 35032 16454
rect 34980 16390 35032 16396
rect 34888 16108 34940 16114
rect 34888 16050 34940 16056
rect 34796 16040 34848 16046
rect 34796 15982 34848 15988
rect 34704 15700 34756 15706
rect 34704 15642 34756 15648
rect 34808 15502 34836 15982
rect 34900 15910 34928 16050
rect 34992 16046 35020 16390
rect 35164 16176 35216 16182
rect 35162 16144 35164 16153
rect 35216 16144 35218 16153
rect 35162 16079 35218 16088
rect 34980 16040 35032 16046
rect 34980 15982 35032 15988
rect 34888 15904 34940 15910
rect 34888 15846 34940 15852
rect 35268 15858 35296 16782
rect 35348 16730 35400 16736
rect 35268 15830 35301 15858
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35273 15722 35301 15830
rect 34980 15700 35032 15706
rect 34980 15642 35032 15648
rect 35268 15694 35301 15722
rect 34796 15496 34848 15502
rect 34796 15438 34848 15444
rect 34992 15162 35020 15642
rect 34980 15156 35032 15162
rect 34980 15098 35032 15104
rect 34612 14952 34664 14958
rect 34612 14894 34664 14900
rect 35268 14770 35296 15694
rect 35452 15094 35480 16934
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 36084 15360 36136 15366
rect 36084 15302 36136 15308
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 35440 15088 35492 15094
rect 35440 15030 35492 15036
rect 35348 15020 35400 15026
rect 35348 14962 35400 14968
rect 35268 14742 35301 14770
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35273 14634 35301 14742
rect 35268 14606 35301 14634
rect 34704 14000 34756 14006
rect 34704 13942 34756 13948
rect 34716 13326 34744 13942
rect 35268 13682 35296 14606
rect 35360 14278 35388 14962
rect 35348 14272 35400 14278
rect 35348 14214 35400 14220
rect 35268 13654 35301 13682
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35273 13546 35301 13654
rect 35268 13518 35301 13546
rect 34704 13320 34756 13326
rect 34704 13262 34756 13268
rect 34796 13252 34848 13258
rect 34796 13194 34848 13200
rect 34702 13152 34758 13161
rect 34702 13087 34758 13096
rect 34612 12776 34664 12782
rect 34612 12718 34664 12724
rect 34624 12306 34652 12718
rect 34716 12322 34744 13087
rect 34808 12850 34836 13194
rect 34796 12844 34848 12850
rect 34796 12786 34848 12792
rect 34808 12442 34836 12786
rect 35268 12594 35296 13518
rect 35360 13190 35388 14214
rect 35452 13394 35480 15030
rect 36096 14618 36124 15302
rect 35900 14612 35952 14618
rect 35900 14554 35952 14560
rect 36084 14612 36136 14618
rect 36084 14554 36136 14560
rect 35912 14414 35940 14554
rect 35900 14408 35952 14414
rect 35900 14350 35952 14356
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 36084 14000 36136 14006
rect 36084 13942 36136 13948
rect 35440 13388 35492 13394
rect 35440 13330 35492 13336
rect 35348 13184 35400 13190
rect 35348 13126 35400 13132
rect 35360 12918 35388 13126
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 35348 12912 35400 12918
rect 35348 12854 35400 12860
rect 35532 12912 35584 12918
rect 35532 12854 35584 12860
rect 35268 12566 35301 12594
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35273 12458 35301 12566
rect 34796 12436 34848 12442
rect 34796 12378 34848 12384
rect 35268 12430 35301 12458
rect 34612 12300 34664 12306
rect 34716 12294 34836 12322
rect 34612 12242 34664 12248
rect 34520 12164 34572 12170
rect 34520 12106 34572 12112
rect 34624 11558 34652 12242
rect 34704 12164 34756 12170
rect 34704 12106 34756 12112
rect 34612 11552 34664 11558
rect 34612 11494 34664 11500
rect 34612 11144 34664 11150
rect 34612 11086 34664 11092
rect 34624 11014 34652 11086
rect 34716 11014 34744 12106
rect 34808 11898 34836 12294
rect 35072 12164 35124 12170
rect 35072 12106 35124 12112
rect 34888 12096 34940 12102
rect 34888 12038 34940 12044
rect 34796 11892 34848 11898
rect 34796 11834 34848 11840
rect 34900 11830 34928 12038
rect 35084 11898 35112 12106
rect 35268 12102 35296 12430
rect 35544 12238 35572 12854
rect 36096 12782 36124 13942
rect 36084 12776 36136 12782
rect 36084 12718 36136 12724
rect 35348 12232 35400 12238
rect 35348 12174 35400 12180
rect 35532 12232 35584 12238
rect 35532 12174 35584 12180
rect 35256 12096 35308 12102
rect 35256 12038 35308 12044
rect 35072 11892 35124 11898
rect 35072 11834 35124 11840
rect 34888 11824 34940 11830
rect 34794 11792 34850 11801
rect 34888 11766 34940 11772
rect 34794 11727 34850 11736
rect 34612 11008 34664 11014
rect 34612 10950 34664 10956
rect 34704 11008 34756 11014
rect 34704 10950 34756 10956
rect 34520 10056 34572 10062
rect 34520 9998 34572 10004
rect 34428 9716 34480 9722
rect 34428 9658 34480 9664
rect 34256 9608 34376 9636
rect 34532 9625 34560 9998
rect 33876 9580 33928 9586
rect 33876 9522 33928 9528
rect 34152 9580 34204 9586
rect 34152 9522 34204 9528
rect 33784 8628 33836 8634
rect 33784 8570 33836 8576
rect 33888 8430 33916 9522
rect 34242 8936 34298 8945
rect 34242 8871 34298 8880
rect 34256 8634 34284 8871
rect 33968 8628 34020 8634
rect 33968 8570 34020 8576
rect 34244 8628 34296 8634
rect 34244 8570 34296 8576
rect 33980 8498 34008 8570
rect 34060 8560 34112 8566
rect 34060 8502 34112 8508
rect 33968 8492 34020 8498
rect 33968 8434 34020 8440
rect 33876 8424 33928 8430
rect 33876 8366 33928 8372
rect 33692 8356 33744 8362
rect 33692 8298 33744 8304
rect 33520 8044 33640 8072
rect 33506 7984 33562 7993
rect 33416 7948 33468 7954
rect 33506 7919 33508 7928
rect 33416 7890 33468 7896
rect 33560 7919 33562 7928
rect 33508 7890 33560 7896
rect 33324 7812 33376 7818
rect 33324 7754 33376 7760
rect 33428 7546 33456 7890
rect 33416 7540 33468 7546
rect 33416 7482 33468 7488
rect 32404 7404 32456 7410
rect 32404 7346 32456 7352
rect 31300 7336 31352 7342
rect 31300 7278 31352 7284
rect 31576 7336 31628 7342
rect 31576 7278 31628 7284
rect 31668 7336 31720 7342
rect 31668 7278 31720 7284
rect 32312 7336 32364 7342
rect 32312 7278 32364 7284
rect 31312 7206 31340 7278
rect 31208 7200 31260 7206
rect 31208 7142 31260 7148
rect 31300 7200 31352 7206
rect 31300 7142 31352 7148
rect 29920 6792 29972 6798
rect 29920 6734 29972 6740
rect 30196 6792 30248 6798
rect 30196 6734 30248 6740
rect 30104 6656 30156 6662
rect 30104 6598 30156 6604
rect 30196 6656 30248 6662
rect 30196 6598 30248 6604
rect 30116 6458 30144 6598
rect 29552 6452 29604 6458
rect 29552 6394 29604 6400
rect 30104 6452 30156 6458
rect 30104 6394 30156 6400
rect 30208 6390 30236 6598
rect 30196 6384 30248 6390
rect 29550 6352 29606 6361
rect 30196 6326 30248 6332
rect 29550 6287 29606 6296
rect 29460 6112 29512 6118
rect 29460 6054 29512 6060
rect 29184 5704 29236 5710
rect 29184 5646 29236 5652
rect 29472 5642 29500 6054
rect 29564 5914 29592 6287
rect 29552 5908 29604 5914
rect 29552 5850 29604 5856
rect 29460 5636 29512 5642
rect 29460 5578 29512 5584
rect 29092 5568 29144 5574
rect 29092 5510 29144 5516
rect 29104 5370 29132 5510
rect 29092 5364 29144 5370
rect 29092 5306 29144 5312
rect 29182 5264 29238 5273
rect 29000 5228 29052 5234
rect 30208 5234 30236 6326
rect 31680 6322 31708 7278
rect 33612 6866 33640 8044
rect 33600 6860 33652 6866
rect 33600 6802 33652 6808
rect 33704 6798 33732 8298
rect 33784 7880 33836 7886
rect 33784 7822 33836 7828
rect 33796 7410 33824 7822
rect 33784 7404 33836 7410
rect 33784 7346 33836 7352
rect 33888 7002 33916 8366
rect 33980 7750 34008 8434
rect 33968 7744 34020 7750
rect 33968 7686 34020 7692
rect 33980 7410 34008 7686
rect 33968 7404 34020 7410
rect 33968 7346 34020 7352
rect 34072 7342 34100 8502
rect 34348 8401 34376 9608
rect 34518 9616 34574 9625
rect 34518 9551 34520 9560
rect 34572 9551 34574 9560
rect 34624 9568 34652 10950
rect 34716 10674 34744 10950
rect 34704 10668 34756 10674
rect 34704 10610 34756 10616
rect 34704 10464 34756 10470
rect 34704 10406 34756 10412
rect 34716 10266 34744 10406
rect 34704 10260 34756 10266
rect 34704 10202 34756 10208
rect 34704 9580 34756 9586
rect 34520 9522 34572 9528
rect 34624 9540 34704 9568
rect 34624 9382 34652 9540
rect 34808 9568 34836 11727
rect 35084 11642 35112 11834
rect 35360 11762 35388 12174
rect 35440 12096 35492 12102
rect 35440 12038 35492 12044
rect 35348 11756 35400 11762
rect 35348 11698 35400 11704
rect 35084 11614 35296 11642
rect 35268 11506 35296 11614
rect 35268 11478 35301 11506
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35273 11370 35301 11478
rect 35268 11342 35301 11370
rect 34978 11248 35034 11257
rect 34978 11183 35034 11192
rect 34992 11150 35020 11183
rect 34980 11144 35032 11150
rect 34980 11086 35032 11092
rect 34888 11008 34940 11014
rect 34886 10976 34888 10985
rect 34940 10976 34942 10985
rect 34886 10911 34942 10920
rect 35268 10418 35296 11342
rect 35360 11218 35388 11698
rect 35348 11212 35400 11218
rect 35348 11154 35400 11160
rect 35348 10464 35400 10470
rect 35268 10390 35301 10418
rect 35348 10406 35400 10412
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35273 10282 35301 10390
rect 35268 10254 35301 10282
rect 35268 10146 35296 10254
rect 35176 10130 35296 10146
rect 35164 10124 35296 10130
rect 35216 10118 35296 10124
rect 35164 10066 35216 10072
rect 35072 10056 35124 10062
rect 35072 9998 35124 10004
rect 35084 9761 35112 9998
rect 35070 9752 35126 9761
rect 35070 9687 35126 9696
rect 34888 9580 34940 9586
rect 34808 9540 34888 9568
rect 34704 9522 34756 9528
rect 34888 9522 34940 9528
rect 35176 9466 35204 10066
rect 35256 9920 35308 9926
rect 35256 9862 35308 9868
rect 34808 9438 35204 9466
rect 34612 9376 34664 9382
rect 34612 9318 34664 9324
rect 34428 8900 34480 8906
rect 34428 8842 34480 8848
rect 34440 8412 34468 8842
rect 34520 8832 34572 8838
rect 34520 8774 34572 8780
rect 34532 8634 34560 8774
rect 34520 8628 34572 8634
rect 34520 8570 34572 8576
rect 34532 8514 34560 8570
rect 34532 8486 34652 8514
rect 34520 8424 34572 8430
rect 34334 8392 34390 8401
rect 34440 8384 34520 8412
rect 34520 8366 34572 8372
rect 34334 8327 34390 8336
rect 34348 7410 34376 8327
rect 34532 7818 34560 8366
rect 34520 7812 34572 7818
rect 34520 7754 34572 7760
rect 34624 7750 34652 8486
rect 34704 8356 34756 8362
rect 34704 8298 34756 8304
rect 34716 7886 34744 8298
rect 34808 7954 34836 9438
rect 35268 9330 35296 9862
rect 35360 9722 35388 10406
rect 35452 9926 35480 12038
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 35992 11144 36044 11150
rect 35992 11086 36044 11092
rect 36004 10962 36032 11086
rect 36096 11082 36124 12718
rect 36084 11076 36136 11082
rect 36084 11018 36136 11024
rect 36188 10962 36216 17614
rect 36280 11762 36308 20810
rect 36372 19786 36400 20878
rect 36544 20528 36596 20534
rect 36544 20470 36596 20476
rect 36452 19848 36504 19854
rect 36452 19790 36504 19796
rect 36360 19780 36412 19786
rect 36360 19722 36412 19728
rect 36360 19440 36412 19446
rect 36360 19382 36412 19388
rect 36372 16590 36400 19382
rect 36464 19378 36492 19790
rect 36452 19372 36504 19378
rect 36452 19314 36504 19320
rect 36556 19174 36584 20470
rect 36544 19168 36596 19174
rect 36544 19110 36596 19116
rect 36544 18964 36596 18970
rect 36544 18906 36596 18912
rect 36452 18284 36504 18290
rect 36452 18226 36504 18232
rect 36464 17660 36492 18226
rect 36556 17814 36584 18906
rect 36544 17808 36596 17814
rect 36544 17750 36596 17756
rect 36544 17672 36596 17678
rect 36464 17632 36544 17660
rect 36464 17134 36492 17632
rect 36544 17614 36596 17620
rect 36452 17128 36504 17134
rect 36452 17070 36504 17076
rect 36648 16946 36676 24686
rect 36556 16918 36676 16946
rect 36452 16788 36504 16794
rect 36452 16730 36504 16736
rect 36360 16584 36412 16590
rect 36360 16526 36412 16532
rect 36464 14770 36492 16730
rect 36556 16114 36584 16918
rect 36636 16584 36688 16590
rect 36636 16526 36688 16532
rect 36544 16108 36596 16114
rect 36544 16050 36596 16056
rect 36556 15638 36584 16050
rect 36648 15638 36676 16526
rect 36544 15632 36596 15638
rect 36544 15574 36596 15580
rect 36636 15632 36688 15638
rect 36636 15574 36688 15580
rect 36464 14742 36584 14770
rect 36452 14612 36504 14618
rect 36452 14554 36504 14560
rect 36464 12434 36492 14554
rect 36556 12594 36584 14742
rect 36648 14414 36676 15574
rect 36740 14498 36768 24890
rect 36832 24750 36860 25298
rect 36924 25294 36952 27270
rect 37016 25838 37044 27882
rect 37096 27668 37148 27674
rect 37096 27610 37148 27616
rect 37108 27169 37136 27610
rect 37476 27554 37504 29582
rect 37752 29073 37780 30382
rect 37924 30330 37976 30336
rect 37832 30048 37884 30054
rect 37832 29990 37884 29996
rect 37844 29646 37872 29990
rect 37832 29640 37884 29646
rect 37832 29582 37884 29588
rect 37844 29170 37872 29582
rect 37832 29164 37884 29170
rect 37832 29106 37884 29112
rect 37738 29064 37794 29073
rect 37556 29028 37608 29034
rect 37738 28999 37740 29008
rect 37556 28970 37608 28976
rect 37792 28999 37794 29008
rect 37740 28970 37792 28976
rect 37200 27538 37504 27554
rect 37188 27532 37504 27538
rect 37240 27526 37504 27532
rect 37188 27474 37240 27480
rect 37094 27160 37150 27169
rect 37094 27095 37150 27104
rect 37096 26988 37148 26994
rect 37096 26930 37148 26936
rect 37108 26450 37136 26930
rect 37292 26450 37320 27526
rect 37372 27464 37424 27470
rect 37370 27432 37372 27441
rect 37424 27432 37426 27441
rect 37370 27367 37426 27376
rect 37464 27328 37516 27334
rect 37464 27270 37516 27276
rect 37476 26994 37504 27270
rect 37568 27062 37596 28970
rect 37832 27124 37884 27130
rect 37832 27066 37884 27072
rect 37556 27056 37608 27062
rect 37556 26998 37608 27004
rect 37464 26988 37516 26994
rect 37464 26930 37516 26936
rect 37648 26988 37700 26994
rect 37648 26930 37700 26936
rect 37740 26988 37792 26994
rect 37740 26930 37792 26936
rect 37372 26784 37424 26790
rect 37372 26726 37424 26732
rect 37096 26444 37148 26450
rect 37096 26386 37148 26392
rect 37280 26444 37332 26450
rect 37280 26386 37332 26392
rect 37004 25832 37056 25838
rect 37004 25774 37056 25780
rect 37096 25424 37148 25430
rect 37096 25366 37148 25372
rect 36912 25288 36964 25294
rect 36912 25230 36964 25236
rect 36820 24744 36872 24750
rect 36820 24686 36872 24692
rect 36924 19854 36952 25230
rect 37004 24676 37056 24682
rect 37004 24618 37056 24624
rect 37016 21146 37044 24618
rect 37108 24070 37136 25366
rect 37280 24608 37332 24614
rect 37280 24550 37332 24556
rect 37096 24064 37148 24070
rect 37096 24006 37148 24012
rect 37292 23497 37320 24550
rect 37278 23488 37334 23497
rect 37278 23423 37334 23432
rect 37280 23316 37332 23322
rect 37280 23258 37332 23264
rect 37292 21894 37320 23258
rect 37384 23050 37412 26726
rect 37556 26512 37608 26518
rect 37556 26454 37608 26460
rect 37464 25356 37516 25362
rect 37464 25298 37516 25304
rect 37476 24818 37504 25298
rect 37464 24812 37516 24818
rect 37464 24754 37516 24760
rect 37568 23730 37596 26454
rect 37660 25906 37688 26930
rect 37752 26382 37780 26930
rect 37844 26382 37872 27066
rect 37740 26376 37792 26382
rect 37740 26318 37792 26324
rect 37832 26376 37884 26382
rect 37832 26318 37884 26324
rect 37648 25900 37700 25906
rect 37648 25842 37700 25848
rect 37740 25152 37792 25158
rect 37740 25094 37792 25100
rect 37752 24818 37780 25094
rect 37936 24834 37964 30330
rect 38016 30184 38068 30190
rect 38016 30126 38068 30132
rect 38028 29782 38056 30126
rect 38016 29776 38068 29782
rect 38016 29718 38068 29724
rect 38016 29504 38068 29510
rect 38016 29446 38068 29452
rect 38028 28558 38056 29446
rect 38120 28762 38148 30602
rect 38212 30258 38240 31282
rect 38304 30938 38332 31758
rect 38384 31748 38436 31754
rect 38384 31690 38436 31696
rect 38396 31482 38424 31690
rect 38580 31482 38608 31758
rect 38384 31476 38436 31482
rect 38384 31418 38436 31424
rect 38568 31476 38620 31482
rect 38568 31418 38620 31424
rect 38580 31385 38608 31418
rect 38566 31376 38622 31385
rect 38566 31311 38622 31320
rect 38568 31136 38620 31142
rect 38568 31078 38620 31084
rect 38292 30932 38344 30938
rect 38292 30874 38344 30880
rect 38304 30734 38332 30874
rect 38292 30728 38344 30734
rect 38292 30670 38344 30676
rect 38200 30252 38252 30258
rect 38200 30194 38252 30200
rect 38212 29170 38240 30194
rect 38476 30184 38528 30190
rect 38396 30132 38476 30138
rect 38396 30126 38528 30132
rect 38396 30110 38516 30126
rect 38292 30048 38344 30054
rect 38292 29990 38344 29996
rect 38200 29164 38252 29170
rect 38200 29106 38252 29112
rect 38200 29028 38252 29034
rect 38200 28970 38252 28976
rect 38108 28756 38160 28762
rect 38108 28698 38160 28704
rect 38016 28552 38068 28558
rect 38016 28494 38068 28500
rect 38120 28490 38148 28698
rect 38108 28484 38160 28490
rect 38108 28426 38160 28432
rect 38108 27532 38160 27538
rect 38108 27474 38160 27480
rect 38016 27464 38068 27470
rect 38016 27406 38068 27412
rect 38028 27130 38056 27406
rect 38016 27124 38068 27130
rect 38016 27066 38068 27072
rect 38120 27033 38148 27474
rect 38106 27024 38162 27033
rect 38106 26959 38162 26968
rect 38016 26852 38068 26858
rect 38016 26794 38068 26800
rect 38028 26042 38056 26794
rect 38120 26450 38148 26959
rect 38108 26444 38160 26450
rect 38108 26386 38160 26392
rect 38212 26330 38240 28970
rect 38304 28694 38332 29990
rect 38396 29850 38424 30110
rect 38384 29844 38436 29850
rect 38384 29786 38436 29792
rect 38396 29714 38516 29730
rect 38384 29708 38516 29714
rect 38436 29702 38516 29708
rect 38384 29650 38436 29656
rect 38384 29572 38436 29578
rect 38384 29514 38436 29520
rect 38396 28762 38424 29514
rect 38488 29238 38516 29702
rect 38476 29232 38528 29238
rect 38476 29174 38528 29180
rect 38384 28756 38436 28762
rect 38384 28698 38436 28704
rect 38292 28688 38344 28694
rect 38292 28630 38344 28636
rect 38384 26988 38436 26994
rect 38384 26930 38436 26936
rect 38292 26852 38344 26858
rect 38292 26794 38344 26800
rect 38120 26302 38240 26330
rect 38304 26330 38332 26794
rect 38396 26586 38424 26930
rect 38384 26580 38436 26586
rect 38384 26522 38436 26528
rect 38476 26512 38528 26518
rect 38476 26454 38528 26460
rect 38382 26344 38438 26353
rect 38304 26302 38382 26330
rect 38016 26036 38068 26042
rect 38016 25978 38068 25984
rect 38016 25696 38068 25702
rect 38016 25638 38068 25644
rect 38028 25294 38056 25638
rect 38016 25288 38068 25294
rect 38016 25230 38068 25236
rect 37936 24818 38056 24834
rect 37740 24812 37792 24818
rect 37936 24812 38068 24818
rect 37936 24806 38016 24812
rect 37740 24754 37792 24760
rect 38016 24754 38068 24760
rect 37924 24744 37976 24750
rect 38120 24698 38148 26302
rect 38382 26279 38384 26288
rect 38436 26279 38438 26288
rect 38384 26250 38436 26256
rect 38488 25906 38516 26454
rect 38476 25900 38528 25906
rect 38476 25842 38528 25848
rect 38476 25152 38528 25158
rect 38476 25094 38528 25100
rect 38198 24848 38254 24857
rect 38198 24783 38254 24792
rect 38292 24812 38344 24818
rect 38212 24750 38240 24783
rect 38292 24754 38344 24760
rect 37924 24686 37976 24692
rect 37936 24410 37964 24686
rect 38028 24670 38148 24698
rect 38200 24744 38252 24750
rect 38200 24686 38252 24692
rect 37924 24404 37976 24410
rect 37924 24346 37976 24352
rect 37832 24268 37884 24274
rect 37832 24210 37884 24216
rect 37556 23724 37608 23730
rect 37608 23684 37688 23712
rect 37556 23666 37608 23672
rect 37556 23248 37608 23254
rect 37556 23190 37608 23196
rect 37372 23044 37424 23050
rect 37372 22986 37424 22992
rect 37464 22500 37516 22506
rect 37464 22442 37516 22448
rect 37476 22166 37504 22442
rect 37464 22160 37516 22166
rect 37464 22102 37516 22108
rect 37280 21888 37332 21894
rect 37280 21830 37332 21836
rect 37280 21344 37332 21350
rect 37280 21286 37332 21292
rect 37004 21140 37056 21146
rect 37004 21082 37056 21088
rect 37004 21004 37056 21010
rect 37004 20946 37056 20952
rect 36912 19848 36964 19854
rect 36912 19790 36964 19796
rect 36820 19168 36872 19174
rect 36820 19110 36872 19116
rect 36832 16794 36860 19110
rect 36820 16788 36872 16794
rect 36820 16730 36872 16736
rect 36832 16658 36860 16730
rect 36912 16720 36964 16726
rect 36912 16662 36964 16668
rect 36820 16652 36872 16658
rect 36820 16594 36872 16600
rect 36818 16552 36874 16561
rect 36818 16487 36874 16496
rect 36832 16182 36860 16487
rect 36820 16176 36872 16182
rect 36820 16118 36872 16124
rect 36924 15502 36952 16662
rect 37016 16454 37044 20946
rect 37292 20942 37320 21286
rect 37280 20936 37332 20942
rect 37280 20878 37332 20884
rect 37280 20800 37332 20806
rect 37280 20742 37332 20748
rect 37096 20392 37148 20398
rect 37096 20334 37148 20340
rect 37108 17746 37136 20334
rect 37292 19854 37320 20742
rect 37280 19848 37332 19854
rect 37186 19816 37242 19825
rect 37280 19790 37332 19796
rect 37186 19751 37188 19760
rect 37240 19751 37242 19760
rect 37188 19722 37240 19728
rect 37372 19712 37424 19718
rect 37372 19654 37424 19660
rect 37464 19712 37516 19718
rect 37464 19654 37516 19660
rect 37188 19508 37240 19514
rect 37188 19450 37240 19456
rect 37096 17740 37148 17746
rect 37096 17682 37148 17688
rect 37096 17128 37148 17134
rect 37096 17070 37148 17076
rect 37004 16448 37056 16454
rect 37004 16390 37056 16396
rect 37108 15910 37136 17070
rect 37096 15904 37148 15910
rect 37096 15846 37148 15852
rect 36912 15496 36964 15502
rect 36912 15438 36964 15444
rect 36910 15328 36966 15337
rect 36910 15263 36966 15272
rect 36740 14470 36860 14498
rect 36832 14414 36860 14470
rect 36636 14408 36688 14414
rect 36636 14350 36688 14356
rect 36820 14408 36872 14414
rect 36820 14350 36872 14356
rect 36832 14006 36860 14350
rect 36820 14000 36872 14006
rect 36820 13942 36872 13948
rect 36924 13938 36952 15263
rect 37004 14068 37056 14074
rect 37004 14010 37056 14016
rect 36728 13932 36780 13938
rect 36728 13874 36780 13880
rect 36912 13932 36964 13938
rect 36912 13874 36964 13880
rect 36740 13530 36768 13874
rect 36820 13796 36872 13802
rect 36820 13738 36872 13744
rect 36832 13530 36860 13738
rect 36728 13524 36780 13530
rect 36728 13466 36780 13472
rect 36820 13524 36872 13530
rect 36820 13466 36872 13472
rect 36556 12566 36676 12594
rect 36464 12406 36584 12434
rect 36556 11762 36584 12406
rect 36648 12306 36676 12566
rect 36636 12300 36688 12306
rect 36636 12242 36688 12248
rect 36648 11762 36676 12242
rect 36268 11756 36320 11762
rect 36268 11698 36320 11704
rect 36544 11756 36596 11762
rect 36544 11698 36596 11704
rect 36636 11756 36688 11762
rect 36820 11756 36872 11762
rect 36688 11716 36768 11744
rect 36636 11698 36688 11704
rect 36004 10934 36216 10962
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 36084 10532 36136 10538
rect 36084 10474 36136 10480
rect 35440 9920 35492 9926
rect 35440 9862 35492 9868
rect 35348 9716 35400 9722
rect 35348 9658 35400 9664
rect 35348 9580 35400 9586
rect 35348 9522 35400 9528
rect 35268 9302 35301 9330
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 35273 9194 35301 9302
rect 35268 9166 35301 9194
rect 35360 9178 35388 9522
rect 35348 9172 35400 9178
rect 35164 8968 35216 8974
rect 35164 8910 35216 8916
rect 34980 8832 35032 8838
rect 34980 8774 35032 8780
rect 34992 8430 35020 8774
rect 34980 8424 35032 8430
rect 34980 8366 35032 8372
rect 35176 8294 35204 8910
rect 35268 8838 35296 9166
rect 35348 9114 35400 9120
rect 35360 9081 35388 9114
rect 35346 9072 35402 9081
rect 35346 9007 35402 9016
rect 35452 8974 35480 9862
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 36096 9654 36124 10474
rect 35624 9648 35676 9654
rect 36084 9648 36136 9654
rect 35624 9590 35676 9596
rect 35990 9616 36046 9625
rect 35532 9580 35584 9586
rect 35532 9522 35584 9528
rect 35544 9382 35572 9522
rect 35532 9376 35584 9382
rect 35532 9318 35584 9324
rect 35440 8968 35492 8974
rect 35440 8910 35492 8916
rect 35256 8832 35308 8838
rect 35636 8820 35664 9590
rect 36084 9590 36136 9596
rect 35990 9551 35992 9560
rect 36044 9551 36046 9560
rect 35992 9522 36044 9528
rect 36096 9330 36124 9590
rect 36188 9450 36216 10934
rect 36280 9722 36308 11698
rect 36740 11150 36768 11716
rect 36820 11698 36872 11704
rect 36832 11665 36860 11698
rect 36818 11656 36874 11665
rect 36818 11591 36874 11600
rect 36636 11144 36688 11150
rect 36634 11112 36636 11121
rect 36728 11144 36780 11150
rect 36688 11112 36690 11121
rect 36728 11086 36780 11092
rect 36634 11047 36690 11056
rect 36360 9988 36412 9994
rect 36360 9930 36412 9936
rect 36636 9988 36688 9994
rect 36636 9930 36688 9936
rect 36268 9716 36320 9722
rect 36268 9658 36320 9664
rect 36268 9580 36320 9586
rect 36268 9522 36320 9528
rect 36280 9450 36308 9522
rect 36372 9518 36400 9930
rect 36648 9722 36676 9930
rect 36636 9716 36688 9722
rect 36636 9658 36688 9664
rect 36452 9648 36504 9654
rect 36452 9590 36504 9596
rect 36360 9512 36412 9518
rect 36360 9454 36412 9460
rect 36176 9444 36228 9450
rect 36176 9386 36228 9392
rect 36268 9444 36320 9450
rect 36268 9386 36320 9392
rect 36464 9330 36492 9590
rect 36544 9580 36596 9586
rect 36544 9522 36596 9528
rect 36096 9302 36492 9330
rect 36084 8968 36136 8974
rect 36084 8910 36136 8916
rect 35256 8774 35308 8780
rect 35360 8792 35664 8820
rect 35164 8288 35216 8294
rect 35164 8230 35216 8236
rect 35268 8242 35296 8774
rect 35268 8214 35301 8242
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35273 8106 35301 8214
rect 35268 8078 35301 8106
rect 34796 7948 34848 7954
rect 34796 7890 34848 7896
rect 34704 7880 34756 7886
rect 34704 7822 34756 7828
rect 34612 7744 34664 7750
rect 34612 7686 34664 7692
rect 34624 7410 34652 7686
rect 34716 7546 34744 7822
rect 35072 7744 35124 7750
rect 35072 7686 35124 7692
rect 34704 7540 34756 7546
rect 34704 7482 34756 7488
rect 35084 7410 35112 7686
rect 34336 7404 34388 7410
rect 34336 7346 34388 7352
rect 34612 7404 34664 7410
rect 34612 7346 34664 7352
rect 35072 7404 35124 7410
rect 35072 7346 35124 7352
rect 34060 7336 34112 7342
rect 34060 7278 34112 7284
rect 35072 7268 35124 7274
rect 35268 7256 35296 8078
rect 35360 7342 35388 8792
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 36096 8634 36124 8910
rect 36176 8900 36228 8906
rect 36176 8842 36228 8848
rect 36188 8634 36216 8842
rect 36084 8628 36136 8634
rect 36084 8570 36136 8576
rect 36176 8628 36228 8634
rect 36176 8570 36228 8576
rect 35440 8560 35492 8566
rect 35440 8502 35492 8508
rect 35452 7954 35480 8502
rect 35992 8016 36044 8022
rect 35992 7958 36044 7964
rect 35440 7948 35492 7954
rect 35440 7890 35492 7896
rect 35452 7410 35480 7890
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 36004 7410 36032 7958
rect 36096 7886 36124 8570
rect 36188 8362 36216 8570
rect 36556 8498 36584 9522
rect 36820 9376 36872 9382
rect 36820 9318 36872 9324
rect 36544 8492 36596 8498
rect 36544 8434 36596 8440
rect 36176 8356 36228 8362
rect 36176 8298 36228 8304
rect 36188 8090 36216 8298
rect 36832 8090 36860 9318
rect 36176 8084 36228 8090
rect 36176 8026 36228 8032
rect 36820 8084 36872 8090
rect 36820 8026 36872 8032
rect 36084 7880 36136 7886
rect 36084 7822 36136 7828
rect 37016 7818 37044 14010
rect 37108 11218 37136 15846
rect 37200 14006 37228 19450
rect 37384 17898 37412 19654
rect 37476 18154 37504 19654
rect 37464 18148 37516 18154
rect 37464 18090 37516 18096
rect 37568 18034 37596 23190
rect 37660 20398 37688 23684
rect 37740 22228 37792 22234
rect 37740 22170 37792 22176
rect 37648 20392 37700 20398
rect 37648 20334 37700 20340
rect 37568 18006 37688 18034
rect 37384 17870 37596 17898
rect 37278 17776 37334 17785
rect 37278 17711 37334 17720
rect 37292 16425 37320 17711
rect 37372 17604 37424 17610
rect 37372 17546 37424 17552
rect 37384 16726 37412 17546
rect 37372 16720 37424 16726
rect 37372 16662 37424 16668
rect 37278 16416 37334 16425
rect 37278 16351 37334 16360
rect 37280 14272 37332 14278
rect 37280 14214 37332 14220
rect 37188 14000 37240 14006
rect 37188 13942 37240 13948
rect 37292 13734 37320 14214
rect 37280 13728 37332 13734
rect 37280 13670 37332 13676
rect 37188 12436 37240 12442
rect 37188 12378 37240 12384
rect 37096 11212 37148 11218
rect 37096 11154 37148 11160
rect 37200 10130 37228 12378
rect 37292 11354 37320 13670
rect 37384 11694 37412 16662
rect 37464 16584 37516 16590
rect 37464 16526 37516 16532
rect 37476 16114 37504 16526
rect 37464 16108 37516 16114
rect 37464 16050 37516 16056
rect 37464 15428 37516 15434
rect 37464 15370 37516 15376
rect 37476 14618 37504 15370
rect 37568 14890 37596 17870
rect 37556 14884 37608 14890
rect 37556 14826 37608 14832
rect 37464 14612 37516 14618
rect 37464 14554 37516 14560
rect 37476 13938 37504 14554
rect 37464 13932 37516 13938
rect 37464 13874 37516 13880
rect 37556 13932 37608 13938
rect 37556 13874 37608 13880
rect 37372 11688 37424 11694
rect 37372 11630 37424 11636
rect 37280 11348 37332 11354
rect 37280 11290 37332 11296
rect 37280 11144 37332 11150
rect 37280 11086 37332 11092
rect 37292 10266 37320 11086
rect 37568 10810 37596 13874
rect 37660 13870 37688 18006
rect 37648 13864 37700 13870
rect 37648 13806 37700 13812
rect 37556 10804 37608 10810
rect 37556 10746 37608 10752
rect 37556 10668 37608 10674
rect 37556 10610 37608 10616
rect 37280 10260 37332 10266
rect 37280 10202 37332 10208
rect 37188 10124 37240 10130
rect 37188 10066 37240 10072
rect 37200 9518 37228 10066
rect 37568 10062 37596 10610
rect 37752 10606 37780 22170
rect 37844 12374 37872 24210
rect 37924 23520 37976 23526
rect 37924 23462 37976 23468
rect 37936 22574 37964 23462
rect 38028 23089 38056 24670
rect 38200 24132 38252 24138
rect 38120 24092 38200 24120
rect 38014 23080 38070 23089
rect 38014 23015 38070 23024
rect 38016 22976 38068 22982
rect 38016 22918 38068 22924
rect 38028 22642 38056 22918
rect 38016 22636 38068 22642
rect 38016 22578 38068 22584
rect 37924 22568 37976 22574
rect 37924 22510 37976 22516
rect 38014 22536 38070 22545
rect 38014 22471 38070 22480
rect 37924 22432 37976 22438
rect 37924 22374 37976 22380
rect 37936 22234 37964 22374
rect 37924 22228 37976 22234
rect 37924 22170 37976 22176
rect 37924 22024 37976 22030
rect 37924 21966 37976 21972
rect 37936 19922 37964 21966
rect 38028 20534 38056 22471
rect 38120 21894 38148 24092
rect 38200 24074 38252 24080
rect 38200 23656 38252 23662
rect 38200 23598 38252 23604
rect 38108 21888 38160 21894
rect 38108 21830 38160 21836
rect 38120 21049 38148 21830
rect 38106 21040 38162 21049
rect 38106 20975 38162 20984
rect 38108 20936 38160 20942
rect 38108 20878 38160 20884
rect 38016 20528 38068 20534
rect 38016 20470 38068 20476
rect 38120 20466 38148 20878
rect 38108 20460 38160 20466
rect 38108 20402 38160 20408
rect 38016 20324 38068 20330
rect 38016 20266 38068 20272
rect 37924 19916 37976 19922
rect 37924 19858 37976 19864
rect 38028 19854 38056 20266
rect 38106 19952 38162 19961
rect 38106 19887 38162 19896
rect 38016 19848 38068 19854
rect 38016 19790 38068 19796
rect 38028 18290 38056 19790
rect 38120 19786 38148 19887
rect 38108 19780 38160 19786
rect 38108 19722 38160 19728
rect 38120 19514 38148 19722
rect 38108 19508 38160 19514
rect 38108 19450 38160 19456
rect 38016 18284 38068 18290
rect 38016 18226 38068 18232
rect 37924 16992 37976 16998
rect 37924 16934 37976 16940
rect 37936 15706 37964 16934
rect 38028 16590 38056 18226
rect 38108 17536 38160 17542
rect 38108 17478 38160 17484
rect 38120 17202 38148 17478
rect 38108 17196 38160 17202
rect 38108 17138 38160 17144
rect 38016 16584 38068 16590
rect 38016 16526 38068 16532
rect 37924 15700 37976 15706
rect 37924 15642 37976 15648
rect 38108 13796 38160 13802
rect 38108 13738 38160 13744
rect 38120 13326 38148 13738
rect 38108 13320 38160 13326
rect 38108 13262 38160 13268
rect 38108 13184 38160 13190
rect 38108 13126 38160 13132
rect 38120 12434 38148 13126
rect 37936 12406 38148 12434
rect 37832 12368 37884 12374
rect 37832 12310 37884 12316
rect 37740 10600 37792 10606
rect 37740 10542 37792 10548
rect 37936 10062 37964 12406
rect 38212 12209 38240 23598
rect 38304 23100 38332 24754
rect 38384 23792 38436 23798
rect 38384 23734 38436 23740
rect 38396 23322 38424 23734
rect 38384 23316 38436 23322
rect 38384 23258 38436 23264
rect 38488 23254 38516 25094
rect 38580 24342 38608 31078
rect 38672 29646 38700 31758
rect 38764 30666 38792 33390
rect 39672 32768 39724 32774
rect 39672 32710 39724 32716
rect 39488 31748 39540 31754
rect 39488 31690 39540 31696
rect 38844 31680 38896 31686
rect 38844 31622 38896 31628
rect 38856 31414 38884 31622
rect 39500 31414 39528 31690
rect 38844 31408 38896 31414
rect 38844 31350 38896 31356
rect 39488 31408 39540 31414
rect 39488 31350 39540 31356
rect 38752 30660 38804 30666
rect 38752 30602 38804 30608
rect 39028 30660 39080 30666
rect 39028 30602 39080 30608
rect 38660 29640 38712 29646
rect 38660 29582 38712 29588
rect 38936 29640 38988 29646
rect 38936 29582 38988 29588
rect 38844 29572 38896 29578
rect 38844 29514 38896 29520
rect 38660 29504 38712 29510
rect 38712 29464 38792 29492
rect 38660 29446 38712 29452
rect 38660 27600 38712 27606
rect 38660 27542 38712 27548
rect 38672 26994 38700 27542
rect 38764 27130 38792 29464
rect 38856 28626 38884 29514
rect 38948 29102 38976 29582
rect 38936 29096 38988 29102
rect 38936 29038 38988 29044
rect 38844 28620 38896 28626
rect 38844 28562 38896 28568
rect 38844 27396 38896 27402
rect 38844 27338 38896 27344
rect 38752 27124 38804 27130
rect 38752 27066 38804 27072
rect 38660 26988 38712 26994
rect 38660 26930 38712 26936
rect 38856 26926 38884 27338
rect 38948 26994 38976 29038
rect 38936 26988 38988 26994
rect 38936 26930 38988 26936
rect 38752 26920 38804 26926
rect 38752 26862 38804 26868
rect 38844 26920 38896 26926
rect 38896 26868 38976 26874
rect 38844 26862 38976 26868
rect 38764 26738 38792 26862
rect 38856 26846 38976 26862
rect 38844 26784 38896 26790
rect 38764 26732 38844 26738
rect 38764 26726 38896 26732
rect 38764 26710 38884 26726
rect 38752 25832 38804 25838
rect 38752 25774 38804 25780
rect 38568 24336 38620 24342
rect 38568 24278 38620 24284
rect 38476 23248 38528 23254
rect 38764 23225 38792 25774
rect 38856 24886 38884 26710
rect 38948 26518 38976 26846
rect 38936 26512 38988 26518
rect 38936 26454 38988 26460
rect 38844 24880 38896 24886
rect 38844 24822 38896 24828
rect 38856 23866 38884 24822
rect 38936 24812 38988 24818
rect 38936 24754 38988 24760
rect 38844 23860 38896 23866
rect 38844 23802 38896 23808
rect 38476 23190 38528 23196
rect 38750 23216 38806 23225
rect 38750 23151 38806 23160
rect 38568 23112 38620 23118
rect 38304 23072 38516 23100
rect 38384 22568 38436 22574
rect 38384 22510 38436 22516
rect 38396 22250 38424 22510
rect 38304 22222 38424 22250
rect 38304 20874 38332 22222
rect 38488 20942 38516 23072
rect 38568 23054 38620 23060
rect 38476 20936 38528 20942
rect 38476 20878 38528 20884
rect 38292 20868 38344 20874
rect 38292 20810 38344 20816
rect 38384 20800 38436 20806
rect 38384 20742 38436 20748
rect 38396 20534 38424 20742
rect 38384 20528 38436 20534
rect 38384 20470 38436 20476
rect 38292 20460 38344 20466
rect 38292 20402 38344 20408
rect 38304 18737 38332 20402
rect 38580 19530 38608 23054
rect 38660 23044 38712 23050
rect 38660 22986 38712 22992
rect 38672 22234 38700 22986
rect 38660 22228 38712 22234
rect 38660 22170 38712 22176
rect 38396 19502 38608 19530
rect 38290 18728 38346 18737
rect 38290 18663 38346 18672
rect 38292 18284 38344 18290
rect 38292 18226 38344 18232
rect 38304 18057 38332 18226
rect 38290 18048 38346 18057
rect 38290 17983 38346 17992
rect 38292 17808 38344 17814
rect 38292 17750 38344 17756
rect 38304 17218 38332 17750
rect 38396 17338 38424 19502
rect 38764 19174 38792 23151
rect 38948 21486 38976 24754
rect 38936 21480 38988 21486
rect 38936 21422 38988 21428
rect 38844 20868 38896 20874
rect 38844 20810 38896 20816
rect 38752 19168 38804 19174
rect 38752 19110 38804 19116
rect 38568 18624 38620 18630
rect 38568 18566 38620 18572
rect 38580 18290 38608 18566
rect 38568 18284 38620 18290
rect 38568 18226 38620 18232
rect 38568 18148 38620 18154
rect 38568 18090 38620 18096
rect 38580 17746 38608 18090
rect 38752 18080 38804 18086
rect 38752 18022 38804 18028
rect 38568 17740 38620 17746
rect 38568 17682 38620 17688
rect 38476 17672 38528 17678
rect 38476 17614 38528 17620
rect 38384 17332 38436 17338
rect 38384 17274 38436 17280
rect 38304 17190 38424 17218
rect 38292 16788 38344 16794
rect 38292 16730 38344 16736
rect 38304 15978 38332 16730
rect 38292 15972 38344 15978
rect 38292 15914 38344 15920
rect 38304 15706 38332 15914
rect 38292 15700 38344 15706
rect 38292 15642 38344 15648
rect 38396 15552 38424 17190
rect 38488 16658 38516 17614
rect 38476 16652 38528 16658
rect 38476 16594 38528 16600
rect 38304 15524 38424 15552
rect 38198 12200 38254 12209
rect 38108 12164 38160 12170
rect 38198 12135 38254 12144
rect 38108 12106 38160 12112
rect 38120 11898 38148 12106
rect 38108 11892 38160 11898
rect 38108 11834 38160 11840
rect 38016 11756 38068 11762
rect 38016 11698 38068 11704
rect 37556 10056 37608 10062
rect 37556 9998 37608 10004
rect 37832 10056 37884 10062
rect 37832 9998 37884 10004
rect 37924 10056 37976 10062
rect 37924 9998 37976 10004
rect 37372 9920 37424 9926
rect 37372 9862 37424 9868
rect 37464 9920 37516 9926
rect 37464 9862 37516 9868
rect 37188 9512 37240 9518
rect 37188 9454 37240 9460
rect 37004 7812 37056 7818
rect 37004 7754 37056 7760
rect 36360 7744 36412 7750
rect 36360 7686 36412 7692
rect 37280 7744 37332 7750
rect 37280 7686 37332 7692
rect 35440 7404 35492 7410
rect 35440 7346 35492 7352
rect 35992 7404 36044 7410
rect 35992 7346 36044 7352
rect 35348 7336 35400 7342
rect 35348 7278 35400 7284
rect 35532 7336 35584 7342
rect 35532 7278 35584 7284
rect 35124 7228 35296 7256
rect 35072 7210 35124 7216
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35544 7002 35572 7278
rect 36372 7002 36400 7686
rect 37292 7410 37320 7686
rect 37280 7404 37332 7410
rect 37280 7346 37332 7352
rect 37292 7002 37320 7346
rect 37384 7002 37412 9862
rect 37476 9450 37504 9862
rect 37740 9648 37792 9654
rect 37740 9590 37792 9596
rect 37648 9580 37700 9586
rect 37648 9522 37700 9528
rect 37464 9444 37516 9450
rect 37464 9386 37516 9392
rect 37556 9444 37608 9450
rect 37556 9386 37608 9392
rect 37476 8566 37504 9386
rect 37568 8974 37596 9386
rect 37660 9178 37688 9522
rect 37648 9172 37700 9178
rect 37648 9114 37700 9120
rect 37752 8974 37780 9590
rect 37556 8968 37608 8974
rect 37556 8910 37608 8916
rect 37740 8968 37792 8974
rect 37740 8910 37792 8916
rect 37464 8560 37516 8566
rect 37464 8502 37516 8508
rect 37568 8362 37596 8910
rect 37752 8634 37780 8910
rect 37740 8628 37792 8634
rect 37740 8570 37792 8576
rect 37738 8528 37794 8537
rect 37738 8463 37740 8472
rect 37792 8463 37794 8472
rect 37740 8434 37792 8440
rect 37556 8356 37608 8362
rect 37556 8298 37608 8304
rect 37464 7812 37516 7818
rect 37464 7754 37516 7760
rect 37476 7206 37504 7754
rect 37752 7546 37780 8434
rect 37844 8294 37872 9998
rect 37924 9920 37976 9926
rect 37924 9862 37976 9868
rect 37936 8974 37964 9862
rect 38028 9654 38056 11698
rect 38212 10130 38240 12135
rect 38304 11762 38332 15524
rect 38568 15496 38620 15502
rect 38568 15438 38620 15444
rect 38476 15156 38528 15162
rect 38476 15098 38528 15104
rect 38384 13932 38436 13938
rect 38384 13874 38436 13880
rect 38396 12986 38424 13874
rect 38384 12980 38436 12986
rect 38384 12922 38436 12928
rect 38384 12232 38436 12238
rect 38384 12174 38436 12180
rect 38292 11756 38344 11762
rect 38292 11698 38344 11704
rect 38396 11558 38424 12174
rect 38384 11552 38436 11558
rect 38384 11494 38436 11500
rect 38488 11286 38516 15098
rect 38580 13734 38608 15438
rect 38660 15360 38712 15366
rect 38660 15302 38712 15308
rect 38672 15026 38700 15302
rect 38660 15020 38712 15026
rect 38660 14962 38712 14968
rect 38660 14816 38712 14822
rect 38660 14758 38712 14764
rect 38568 13728 38620 13734
rect 38568 13670 38620 13676
rect 38568 13388 38620 13394
rect 38568 13330 38620 13336
rect 38580 12782 38608 13330
rect 38672 12986 38700 14758
rect 38764 13190 38792 18022
rect 38856 15026 38884 20810
rect 38948 18834 38976 21422
rect 39040 19666 39068 30602
rect 39500 30326 39528 31350
rect 39488 30320 39540 30326
rect 39488 30262 39540 30268
rect 39120 29640 39172 29646
rect 39120 29582 39172 29588
rect 39132 24750 39160 29582
rect 39212 29504 39264 29510
rect 39212 29446 39264 29452
rect 39304 29504 39356 29510
rect 39304 29446 39356 29452
rect 39224 29306 39252 29446
rect 39212 29300 39264 29306
rect 39212 29242 39264 29248
rect 39316 29186 39344 29446
rect 39500 29238 39528 30262
rect 39224 29158 39344 29186
rect 39488 29232 39540 29238
rect 39488 29174 39540 29180
rect 39224 28558 39252 29158
rect 39212 28552 39264 28558
rect 39212 28494 39264 28500
rect 39224 26790 39252 28494
rect 39500 27146 39528 29174
rect 39580 27396 39632 27402
rect 39580 27338 39632 27344
rect 39592 27305 39620 27338
rect 39578 27296 39634 27305
rect 39578 27231 39634 27240
rect 39500 27118 39620 27146
rect 39304 27056 39356 27062
rect 39304 26998 39356 27004
rect 39212 26784 39264 26790
rect 39212 26726 39264 26732
rect 39316 26518 39344 26998
rect 39304 26512 39356 26518
rect 39304 26454 39356 26460
rect 39120 24744 39172 24750
rect 39120 24686 39172 24692
rect 39120 23656 39172 23662
rect 39120 23598 39172 23604
rect 39132 22030 39160 23598
rect 39316 23186 39344 26454
rect 39396 24608 39448 24614
rect 39396 24550 39448 24556
rect 39408 24206 39436 24550
rect 39488 24404 39540 24410
rect 39488 24346 39540 24352
rect 39396 24200 39448 24206
rect 39396 24142 39448 24148
rect 39304 23180 39356 23186
rect 39304 23122 39356 23128
rect 39408 22030 39436 24142
rect 39500 23662 39528 24346
rect 39592 23730 39620 27118
rect 39684 24410 39712 32710
rect 40040 30320 40092 30326
rect 40040 30262 40092 30268
rect 39764 28620 39816 28626
rect 39764 28562 39816 28568
rect 39776 26994 39804 28562
rect 39764 26988 39816 26994
rect 39764 26930 39816 26936
rect 39776 26382 39804 26930
rect 39856 26852 39908 26858
rect 39856 26794 39908 26800
rect 39764 26376 39816 26382
rect 39764 26318 39816 26324
rect 39672 24404 39724 24410
rect 39672 24346 39724 24352
rect 39684 24290 39712 24346
rect 39684 24262 39804 24290
rect 39672 24200 39724 24206
rect 39672 24142 39724 24148
rect 39684 23905 39712 24142
rect 39670 23896 39726 23905
rect 39670 23831 39726 23840
rect 39580 23724 39632 23730
rect 39580 23666 39632 23672
rect 39488 23656 39540 23662
rect 39488 23598 39540 23604
rect 39592 23322 39620 23666
rect 39580 23316 39632 23322
rect 39580 23258 39632 23264
rect 39488 23180 39540 23186
rect 39488 23122 39540 23128
rect 39120 22024 39172 22030
rect 39120 21966 39172 21972
rect 39304 22024 39356 22030
rect 39304 21966 39356 21972
rect 39396 22024 39448 22030
rect 39396 21966 39448 21972
rect 39316 20262 39344 21966
rect 39304 20256 39356 20262
rect 39304 20198 39356 20204
rect 39212 19848 39264 19854
rect 39212 19790 39264 19796
rect 39040 19638 39160 19666
rect 39028 19508 39080 19514
rect 39028 19450 39080 19456
rect 38936 18828 38988 18834
rect 38936 18770 38988 18776
rect 39040 15162 39068 19450
rect 39132 18766 39160 19638
rect 39224 19310 39252 19790
rect 39500 19514 39528 23122
rect 39776 23118 39804 24262
rect 39764 23112 39816 23118
rect 39764 23054 39816 23060
rect 39764 22432 39816 22438
rect 39764 22374 39816 22380
rect 39580 20256 39632 20262
rect 39580 20198 39632 20204
rect 39488 19508 39540 19514
rect 39488 19450 39540 19456
rect 39212 19304 39264 19310
rect 39212 19246 39264 19252
rect 39224 18766 39252 19246
rect 39120 18760 39172 18766
rect 39120 18702 39172 18708
rect 39212 18760 39264 18766
rect 39212 18702 39264 18708
rect 39132 15502 39160 18702
rect 39224 15638 39252 18702
rect 39396 18216 39448 18222
rect 39396 18158 39448 18164
rect 39408 17785 39436 18158
rect 39394 17776 39450 17785
rect 39394 17711 39450 17720
rect 39488 16448 39540 16454
rect 39488 16390 39540 16396
rect 39212 15632 39264 15638
rect 39212 15574 39264 15580
rect 39120 15496 39172 15502
rect 39120 15438 39172 15444
rect 39396 15496 39448 15502
rect 39396 15438 39448 15444
rect 39028 15156 39080 15162
rect 39028 15098 39080 15104
rect 38844 15020 38896 15026
rect 38844 14962 38896 14968
rect 39028 14816 39080 14822
rect 39028 14758 39080 14764
rect 38844 13796 38896 13802
rect 38844 13738 38896 13744
rect 38856 13512 38884 13738
rect 38936 13524 38988 13530
rect 38856 13484 38936 13512
rect 38936 13466 38988 13472
rect 38752 13184 38804 13190
rect 38752 13126 38804 13132
rect 38660 12980 38712 12986
rect 38660 12922 38712 12928
rect 38660 12844 38712 12850
rect 38660 12786 38712 12792
rect 38568 12776 38620 12782
rect 38568 12718 38620 12724
rect 38672 12442 38700 12786
rect 38660 12436 38712 12442
rect 38660 12378 38712 12384
rect 39040 12050 39068 14758
rect 39212 14068 39264 14074
rect 39212 14010 39264 14016
rect 39120 12640 39172 12646
rect 39120 12582 39172 12588
rect 38948 12022 39068 12050
rect 38752 11756 38804 11762
rect 38752 11698 38804 11704
rect 38568 11552 38620 11558
rect 38568 11494 38620 11500
rect 38476 11280 38528 11286
rect 38476 11222 38528 11228
rect 38292 11008 38344 11014
rect 38292 10950 38344 10956
rect 38304 10674 38332 10950
rect 38292 10668 38344 10674
rect 38292 10610 38344 10616
rect 38200 10124 38252 10130
rect 38200 10066 38252 10072
rect 38016 9648 38068 9654
rect 38016 9590 38068 9596
rect 38014 9208 38070 9217
rect 38014 9143 38016 9152
rect 38068 9143 38070 9152
rect 38016 9114 38068 9120
rect 37924 8968 37976 8974
rect 37924 8910 37976 8916
rect 37832 8288 37884 8294
rect 37832 8230 37884 8236
rect 38212 7954 38240 10066
rect 38580 8634 38608 11494
rect 38764 10538 38792 11698
rect 38948 11694 38976 12022
rect 38936 11688 38988 11694
rect 38936 11630 38988 11636
rect 39132 10742 39160 12582
rect 39120 10736 39172 10742
rect 39120 10678 39172 10684
rect 39224 10674 39252 14010
rect 39408 14006 39436 15438
rect 39396 14000 39448 14006
rect 39396 13942 39448 13948
rect 39500 13802 39528 16390
rect 39488 13796 39540 13802
rect 39488 13738 39540 13744
rect 39304 13184 39356 13190
rect 39304 13126 39356 13132
rect 39316 11558 39344 13126
rect 39500 12714 39528 13738
rect 39488 12708 39540 12714
rect 39488 12650 39540 12656
rect 39592 12306 39620 20198
rect 39672 19780 39724 19786
rect 39672 19722 39724 19728
rect 39684 18222 39712 19722
rect 39672 18216 39724 18222
rect 39672 18158 39724 18164
rect 39580 12300 39632 12306
rect 39580 12242 39632 12248
rect 39304 11552 39356 11558
rect 39304 11494 39356 11500
rect 39684 11218 39712 18158
rect 39776 13938 39804 22374
rect 39868 17882 39896 26794
rect 39948 26376 40000 26382
rect 39948 26318 40000 26324
rect 39960 25945 39988 26318
rect 39946 25936 40002 25945
rect 39946 25871 40002 25880
rect 40052 24954 40080 30262
rect 40224 26988 40276 26994
rect 40224 26930 40276 26936
rect 40236 26625 40264 26930
rect 40222 26616 40278 26625
rect 40222 26551 40278 26560
rect 40040 24948 40092 24954
rect 40040 24890 40092 24896
rect 40224 24812 40276 24818
rect 40224 24754 40276 24760
rect 40236 24585 40264 24754
rect 40222 24576 40278 24585
rect 40222 24511 40278 24520
rect 40132 24200 40184 24206
rect 40132 24142 40184 24148
rect 39856 17876 39908 17882
rect 39856 17818 39908 17824
rect 39764 13932 39816 13938
rect 39764 13874 39816 13880
rect 39868 13326 39896 17818
rect 39856 13320 39908 13326
rect 39856 13262 39908 13268
rect 40144 12434 40172 24142
rect 40052 12406 40172 12434
rect 39672 11212 39724 11218
rect 39672 11154 39724 11160
rect 39212 10668 39264 10674
rect 39212 10610 39264 10616
rect 38752 10532 38804 10538
rect 38752 10474 38804 10480
rect 38660 10464 38712 10470
rect 38660 10406 38712 10412
rect 39396 10464 39448 10470
rect 39396 10406 39448 10412
rect 38568 8628 38620 8634
rect 38568 8570 38620 8576
rect 38476 8424 38528 8430
rect 38476 8366 38528 8372
rect 38200 7948 38252 7954
rect 38200 7890 38252 7896
rect 37740 7540 37792 7546
rect 37740 7482 37792 7488
rect 37464 7200 37516 7206
rect 37464 7142 37516 7148
rect 33876 6996 33928 7002
rect 33876 6938 33928 6944
rect 35532 6996 35584 7002
rect 35532 6938 35584 6944
rect 36360 6996 36412 7002
rect 36360 6938 36412 6944
rect 37280 6996 37332 7002
rect 37280 6938 37332 6944
rect 37372 6996 37424 7002
rect 37372 6938 37424 6944
rect 37476 6866 37504 7142
rect 38212 6866 38240 7890
rect 38488 7478 38516 8366
rect 38672 7478 38700 10406
rect 39408 9994 39436 10406
rect 39396 9988 39448 9994
rect 39396 9930 39448 9936
rect 39028 9920 39080 9926
rect 39028 9862 39080 9868
rect 39040 8566 39068 9862
rect 39948 9648 40000 9654
rect 39948 9590 40000 9596
rect 39028 8560 39080 8566
rect 39028 8502 39080 8508
rect 39040 7750 39068 8502
rect 39028 7744 39080 7750
rect 39028 7686 39080 7692
rect 39040 7478 39068 7686
rect 39960 7546 39988 9590
rect 40052 7886 40080 12406
rect 40040 7880 40092 7886
rect 40040 7822 40092 7828
rect 39948 7540 40000 7546
rect 39948 7482 40000 7488
rect 38476 7472 38528 7478
rect 38476 7414 38528 7420
rect 38660 7472 38712 7478
rect 38660 7414 38712 7420
rect 39028 7472 39080 7478
rect 39028 7414 39080 7420
rect 39040 7206 39068 7414
rect 39028 7200 39080 7206
rect 39028 7142 39080 7148
rect 37464 6860 37516 6866
rect 37464 6802 37516 6808
rect 38200 6860 38252 6866
rect 38200 6802 38252 6808
rect 33692 6792 33744 6798
rect 33692 6734 33744 6740
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 31300 6316 31352 6322
rect 31300 6258 31352 6264
rect 31668 6316 31720 6322
rect 31668 6258 31720 6264
rect 31312 5778 31340 6258
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 31300 5772 31352 5778
rect 31300 5714 31352 5720
rect 30288 5636 30340 5642
rect 30288 5578 30340 5584
rect 30300 5370 30328 5578
rect 30288 5364 30340 5370
rect 30288 5306 30340 5312
rect 31312 5302 31340 5714
rect 40052 5522 40080 7822
rect 39960 5494 40080 5522
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 31300 5296 31352 5302
rect 31300 5238 31352 5244
rect 29182 5199 29184 5208
rect 29000 5170 29052 5176
rect 29236 5199 29238 5208
rect 30196 5228 30248 5234
rect 29184 5170 29236 5176
rect 30196 5170 30248 5176
rect 28632 5024 28684 5030
rect 28632 4966 28684 4972
rect 28644 4146 28672 4966
rect 29196 4282 29224 5170
rect 29184 4276 29236 4282
rect 29184 4218 29236 4224
rect 28172 4140 28224 4146
rect 28172 4082 28224 4088
rect 28632 4140 28684 4146
rect 28632 4082 28684 4088
rect 29196 4026 29224 4218
rect 30208 4214 30236 5170
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 39960 4690 39988 5494
rect 39948 4684 40000 4690
rect 39948 4626 40000 4632
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 30196 4208 30248 4214
rect 30196 4150 30248 4156
rect 29196 4010 29316 4026
rect 29196 4004 29328 4010
rect 29196 3998 29276 4004
rect 29276 3946 29328 3952
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 39960 3670 39988 4626
rect 39948 3664 40000 3670
rect 39948 3606 40000 3612
rect 24860 3596 24912 3602
rect 24860 3538 24912 3544
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 26792 3528 26844 3534
rect 26792 3470 26844 3476
rect 40130 3496 40186 3505
rect 24216 3392 24268 3398
rect 24216 3334 24268 3340
rect 24308 3392 24360 3398
rect 24308 3334 24360 3340
rect 24228 3126 24256 3334
rect 23480 3120 23532 3126
rect 23480 3062 23532 3068
rect 23940 3120 23992 3126
rect 23940 3062 23992 3068
rect 24216 3120 24268 3126
rect 24216 3062 24268 3068
rect 24320 3058 24348 3334
rect 26804 3194 26832 3470
rect 40130 3431 40132 3440
rect 40184 3431 40186 3440
rect 40132 3402 40184 3408
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 26792 3188 26844 3194
rect 26792 3130 26844 3136
rect 24308 3052 24360 3058
rect 24308 2994 24360 3000
rect 23388 2984 23440 2990
rect 23388 2926 23440 2932
rect 22940 2746 23060 2774
rect 23124 2746 23244 2774
rect 22744 2508 22796 2514
rect 22744 2450 22796 2456
rect 23032 2446 23060 2746
rect 23020 2440 23072 2446
rect 23020 2382 23072 2388
rect 22468 2372 22520 2378
rect 22468 2314 22520 2320
rect 23216 800 23244 2746
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 23860 800 23888 2246
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 18 0 74 800
rect 662 0 718 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 18050 0 18106 800
rect 19338 0 19394 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 23202 0 23258 800
rect 23846 0 23902 800
<< via2 >>
rect 4880 41370 4936 41372
rect 4960 41370 5016 41372
rect 5040 41370 5096 41372
rect 5120 41370 5176 41372
rect 4880 41318 4926 41370
rect 4926 41318 4936 41370
rect 4960 41318 4990 41370
rect 4990 41318 5002 41370
rect 5002 41318 5016 41370
rect 5040 41318 5054 41370
rect 5054 41318 5066 41370
rect 5066 41318 5096 41370
rect 5120 41318 5130 41370
rect 5130 41318 5176 41370
rect 4880 41316 4936 41318
rect 4960 41316 5016 41318
rect 5040 41316 5096 41318
rect 5120 41316 5176 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4880 40282 4936 40284
rect 4960 40282 5016 40284
rect 5040 40282 5096 40284
rect 5120 40282 5176 40284
rect 4880 40230 4926 40282
rect 4926 40230 4936 40282
rect 4960 40230 4990 40282
rect 4990 40230 5002 40282
rect 5002 40230 5016 40282
rect 5040 40230 5054 40282
rect 5054 40230 5066 40282
rect 5066 40230 5096 40282
rect 5120 40230 5130 40282
rect 5130 40230 5176 40282
rect 4880 40228 4936 40230
rect 4960 40228 5016 40230
rect 5040 40228 5096 40230
rect 5120 40228 5176 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4880 39194 4936 39196
rect 4960 39194 5016 39196
rect 5040 39194 5096 39196
rect 5120 39194 5176 39196
rect 4880 39142 4926 39194
rect 4926 39142 4936 39194
rect 4960 39142 4990 39194
rect 4990 39142 5002 39194
rect 5002 39142 5016 39194
rect 5040 39142 5054 39194
rect 5054 39142 5066 39194
rect 5066 39142 5096 39194
rect 5120 39142 5130 39194
rect 5130 39142 5176 39194
rect 4880 39140 4936 39142
rect 4960 39140 5016 39142
rect 5040 39140 5096 39142
rect 5120 39140 5176 39142
rect 3422 38800 3478 38856
rect 2962 36080 3018 36136
rect 1306 34720 1362 34776
rect 1674 34040 1730 34096
rect 1674 33396 1676 33416
rect 1676 33396 1728 33416
rect 1728 33396 1730 33416
rect 1674 33360 1730 33396
rect 1490 32680 1546 32736
rect 1582 30660 1638 30696
rect 1582 30640 1584 30660
rect 1584 30640 1636 30660
rect 1636 30640 1638 30660
rect 3238 31320 3294 31376
rect 846 30096 902 30152
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 8022 38292 8024 38312
rect 8024 38292 8076 38312
rect 8076 38292 8078 38312
rect 8022 38256 8078 38292
rect 6274 35264 6330 35320
rect 8850 38256 8906 38312
rect 9034 38292 9036 38312
rect 9036 38292 9088 38312
rect 9088 38292 9090 38312
rect 9034 38256 9090 38292
rect 7286 36116 7288 36136
rect 7288 36116 7340 36136
rect 7340 36116 7342 36136
rect 7286 36080 7342 36116
rect 6458 35148 6514 35184
rect 6458 35128 6460 35148
rect 6460 35128 6512 35148
rect 6512 35128 6514 35148
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4802 30796 4858 30832
rect 4802 30776 4804 30796
rect 4804 30776 4856 30796
rect 4856 30776 4858 30796
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4802 25356 4858 25392
rect 4802 25336 4804 25356
rect 4804 25336 4856 25356
rect 4856 25336 4858 25356
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 3514 21528 3570 21584
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 5078 23704 5134 23760
rect 5998 28092 6000 28112
rect 6000 28092 6052 28112
rect 6052 28092 6054 28112
rect 5998 28056 6054 28092
rect 7378 35128 7434 35184
rect 7562 35264 7618 35320
rect 4618 21972 4620 21992
rect 4620 21972 4672 21992
rect 4672 21972 4674 21992
rect 4618 21936 4674 21972
rect 5446 23432 5502 23488
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 3422 20848 3478 20904
rect 3606 21392 3662 21448
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 5170 21528 5226 21584
rect 4894 20984 4950 21040
rect 5078 21004 5134 21040
rect 5078 20984 5080 21004
rect 5080 20984 5132 21004
rect 5132 20984 5134 21004
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 7102 28092 7104 28112
rect 7104 28092 7156 28112
rect 7156 28092 7158 28112
rect 7102 28056 7158 28092
rect 6734 26696 6790 26752
rect 6090 25064 6146 25120
rect 6366 24384 6422 24440
rect 6090 23840 6146 23896
rect 6182 23568 6238 23624
rect 5538 20576 5594 20632
rect 5722 21120 5778 21176
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 3698 18128 3754 18184
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4710 18128 4766 18184
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4894 12844 4950 12880
rect 4894 12824 4896 12844
rect 4896 12824 4948 12844
rect 4948 12824 4950 12844
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 1858 10956 1860 10976
rect 1860 10956 1912 10976
rect 1912 10956 1914 10976
rect 1858 10920 1914 10956
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 6550 24520 6606 24576
rect 6550 23840 6606 23896
rect 6366 20440 6422 20496
rect 5998 20304 6054 20360
rect 6734 21140 6790 21176
rect 6734 21120 6736 21140
rect 6736 21120 6788 21140
rect 6788 21120 6790 21140
rect 6182 19896 6238 19952
rect 7102 25220 7158 25256
rect 7102 25200 7104 25220
rect 7104 25200 7156 25220
rect 7156 25200 7158 25220
rect 7102 21392 7158 21448
rect 7010 20440 7066 20496
rect 5906 12688 5962 12744
rect 7470 23704 7526 23760
rect 7470 21004 7526 21040
rect 7470 20984 7472 21004
rect 7472 20984 7524 21004
rect 7524 20984 7526 21004
rect 7930 24384 7986 24440
rect 9126 36116 9128 36136
rect 9128 36116 9180 36136
rect 9180 36116 9182 36136
rect 9126 36080 9182 36116
rect 8482 32544 8538 32600
rect 8390 26968 8446 27024
rect 8206 25200 8262 25256
rect 8114 24248 8170 24304
rect 8390 25100 8392 25120
rect 8392 25100 8444 25120
rect 8444 25100 8446 25120
rect 8390 25064 8446 25100
rect 6826 12688 6882 12744
rect 5722 10240 5778 10296
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 7562 14476 7618 14512
rect 7562 14456 7564 14476
rect 7564 14456 7616 14476
rect 7616 14456 7618 14476
rect 7470 12860 7472 12880
rect 7472 12860 7524 12880
rect 7524 12860 7526 12880
rect 7470 12824 7526 12860
rect 8206 22344 8262 22400
rect 8666 24012 8668 24032
rect 8668 24012 8720 24032
rect 8720 24012 8722 24032
rect 8666 23976 8722 24012
rect 8666 23840 8722 23896
rect 8574 23704 8630 23760
rect 8206 20984 8262 21040
rect 8942 26560 8998 26616
rect 10138 35944 10194 36000
rect 10506 35692 10562 35728
rect 10506 35672 10508 35692
rect 10508 35672 10560 35692
rect 10560 35672 10562 35692
rect 10138 34992 10194 35048
rect 9862 27920 9918 27976
rect 9034 24520 9090 24576
rect 8942 23976 8998 24032
rect 9310 24384 9366 24440
rect 9218 24248 9274 24304
rect 9126 23704 9182 23760
rect 8758 22208 8814 22264
rect 8114 20304 8170 20360
rect 8574 20576 8630 20632
rect 9034 22380 9036 22400
rect 9036 22380 9088 22400
rect 9088 22380 9090 22400
rect 9034 22344 9090 22380
rect 9678 24248 9734 24304
rect 9586 22208 9642 22264
rect 8758 17856 8814 17912
rect 9770 23044 9826 23080
rect 9770 23024 9772 23044
rect 9772 23024 9824 23044
rect 9824 23024 9826 23044
rect 11058 35944 11114 36000
rect 10966 35692 11022 35728
rect 10966 35672 10968 35692
rect 10968 35672 11020 35692
rect 11020 35672 11022 35692
rect 10966 31728 11022 31784
rect 11150 31592 11206 31648
rect 10782 29708 10838 29744
rect 10782 29688 10784 29708
rect 10784 29688 10836 29708
rect 10836 29688 10838 29708
rect 10690 29588 10692 29608
rect 10692 29588 10744 29608
rect 10744 29588 10746 29608
rect 10690 29552 10746 29588
rect 10690 27240 10746 27296
rect 10690 27104 10746 27160
rect 10230 23296 10286 23352
rect 10414 24812 10470 24848
rect 10414 24792 10416 24812
rect 10416 24792 10468 24812
rect 10468 24792 10470 24812
rect 12254 31728 12310 31784
rect 12254 31592 12310 31648
rect 10966 26444 11022 26480
rect 10966 26424 10968 26444
rect 10968 26424 11020 26444
rect 11020 26424 11022 26444
rect 10230 23024 10286 23080
rect 10414 23044 10470 23080
rect 10414 23024 10416 23044
rect 10416 23024 10468 23044
rect 10468 23024 10470 23044
rect 10690 23024 10746 23080
rect 10506 22072 10562 22128
rect 10506 21548 10562 21584
rect 10506 21528 10508 21548
rect 10508 21528 10560 21548
rect 10560 21528 10562 21548
rect 8022 14456 8078 14512
rect 7010 8900 7066 8936
rect 7010 8880 7012 8900
rect 7012 8880 7064 8900
rect 7064 8880 7066 8900
rect 8758 14476 8814 14512
rect 8758 14456 8760 14476
rect 8760 14456 8812 14476
rect 8812 14456 8814 14476
rect 8942 12708 8998 12744
rect 8942 12688 8944 12708
rect 8944 12688 8996 12708
rect 8996 12688 8998 12708
rect 10506 16652 10562 16688
rect 10506 16632 10508 16652
rect 10508 16632 10560 16652
rect 10560 16632 10562 16652
rect 7010 8372 7012 8392
rect 7012 8372 7064 8392
rect 7064 8372 7066 8392
rect 7010 8336 7066 8372
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 7930 8372 7932 8392
rect 7932 8372 7984 8392
rect 7984 8372 7986 8392
rect 7930 8336 7986 8372
rect 8206 8880 8262 8936
rect 10874 17060 10930 17096
rect 10874 17040 10876 17060
rect 10876 17040 10928 17060
rect 10928 17040 10930 17060
rect 11518 29416 11574 29472
rect 11702 29552 11758 29608
rect 12530 27820 12532 27840
rect 12532 27820 12584 27840
rect 12584 27820 12586 27840
rect 12530 27784 12586 27820
rect 11794 24520 11850 24576
rect 11978 24812 12034 24848
rect 11978 24792 11980 24812
rect 11980 24792 12032 24812
rect 12032 24792 12034 24812
rect 11978 23024 12034 23080
rect 10874 15816 10930 15872
rect 11978 22636 12034 22672
rect 11978 22616 11980 22636
rect 11980 22616 12032 22636
rect 12032 22616 12034 22636
rect 12622 26152 12678 26208
rect 12898 35028 12900 35048
rect 12900 35028 12952 35048
rect 12952 35028 12954 35048
rect 12898 34992 12954 35028
rect 11702 16652 11758 16688
rect 11702 16632 11704 16652
rect 11704 16632 11756 16652
rect 11756 16632 11758 16652
rect 12806 22072 12862 22128
rect 14186 36216 14242 36272
rect 13082 29552 13138 29608
rect 13358 29552 13414 29608
rect 13542 29416 13598 29472
rect 13726 27376 13782 27432
rect 13634 25900 13690 25936
rect 13634 25880 13636 25900
rect 13636 25880 13688 25900
rect 13688 25880 13690 25900
rect 14370 27820 14372 27840
rect 14372 27820 14424 27840
rect 14424 27820 14426 27840
rect 14094 26460 14096 26480
rect 14096 26460 14148 26480
rect 14148 26460 14150 26480
rect 14094 26424 14150 26460
rect 14370 27784 14426 27820
rect 14186 25880 14242 25936
rect 15842 36236 15898 36272
rect 15842 36216 15844 36236
rect 15844 36216 15896 36236
rect 15896 36216 15898 36236
rect 15566 32952 15622 33008
rect 14830 30640 14886 30696
rect 14646 29960 14702 30016
rect 14738 29724 14740 29744
rect 14740 29724 14792 29744
rect 14792 29724 14794 29744
rect 14738 29688 14794 29724
rect 14830 27240 14886 27296
rect 14646 26560 14702 26616
rect 14554 26424 14610 26480
rect 14186 25608 14242 25664
rect 13910 24928 13966 24984
rect 13818 22888 13874 22944
rect 13450 21528 13506 21584
rect 12990 19796 12992 19816
rect 12992 19796 13044 19816
rect 13044 19796 13046 19816
rect 12990 19760 13046 19796
rect 11886 8880 11942 8936
rect 11610 8200 11666 8256
rect 13634 19896 13690 19952
rect 12806 15952 12862 16008
rect 14738 24520 14794 24576
rect 14370 22072 14426 22128
rect 14186 19760 14242 19816
rect 14370 19780 14426 19816
rect 14370 19760 14372 19780
rect 14372 19760 14424 19780
rect 14424 19760 14426 19780
rect 13818 17040 13874 17096
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 11518 6840 11574 6896
rect 12898 12008 12954 12064
rect 14738 22344 14794 22400
rect 15566 30676 15568 30696
rect 15568 30676 15620 30696
rect 15620 30676 15622 30696
rect 15566 30640 15622 30676
rect 15658 30096 15714 30152
rect 15474 29708 15530 29744
rect 15474 29688 15476 29708
rect 15476 29688 15528 29708
rect 15528 29688 15530 29708
rect 15566 27376 15622 27432
rect 16486 32952 16542 33008
rect 16118 31728 16174 31784
rect 16026 30096 16082 30152
rect 16302 29688 16358 29744
rect 15658 26424 15714 26480
rect 17498 35536 17554 35592
rect 18050 35572 18052 35592
rect 18052 35572 18104 35592
rect 18104 35572 18106 35592
rect 18050 35536 18106 35572
rect 18694 35012 18750 35048
rect 18694 34992 18696 35012
rect 18696 34992 18748 35012
rect 18748 34992 18750 35012
rect 16486 27124 16542 27160
rect 16486 27104 16488 27124
rect 16488 27104 16540 27124
rect 16540 27104 16542 27124
rect 16854 26424 16910 26480
rect 15658 26308 15714 26344
rect 15658 26288 15660 26308
rect 15660 26288 15712 26308
rect 15712 26288 15714 26308
rect 15382 23296 15438 23352
rect 14922 19896 14978 19952
rect 15566 19896 15622 19952
rect 15290 19796 15292 19816
rect 15292 19796 15344 19816
rect 15344 19796 15346 19816
rect 15290 19760 15346 19796
rect 15566 18284 15622 18320
rect 15566 18264 15568 18284
rect 15568 18264 15620 18284
rect 15620 18264 15622 18284
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 12530 7384 12586 7440
rect 15198 17040 15254 17096
rect 17774 29144 17830 29200
rect 17222 26988 17278 27024
rect 17222 26968 17224 26988
rect 17224 26968 17276 26988
rect 17276 26968 17278 26988
rect 16946 26288 17002 26344
rect 16302 20460 16358 20496
rect 16302 20440 16304 20460
rect 16304 20440 16356 20460
rect 16356 20440 16358 20460
rect 14094 7928 14150 7984
rect 17314 26188 17316 26208
rect 17316 26188 17368 26208
rect 17368 26188 17370 26208
rect 17314 26152 17370 26188
rect 17130 25200 17186 25256
rect 16946 17720 17002 17776
rect 13910 4120 13966 4176
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 15658 8492 15714 8528
rect 15658 8472 15660 8492
rect 15660 8472 15712 8492
rect 15712 8472 15714 8492
rect 15566 8064 15622 8120
rect 16486 9560 16542 9616
rect 17498 20712 17554 20768
rect 18326 29960 18382 30016
rect 18326 25472 18382 25528
rect 18050 23024 18106 23080
rect 17958 21528 18014 21584
rect 18602 29552 18658 29608
rect 18510 27512 18566 27568
rect 18418 23604 18420 23624
rect 18420 23604 18472 23624
rect 18472 23604 18474 23624
rect 18418 23568 18474 23604
rect 18970 27512 19026 27568
rect 20534 35028 20536 35048
rect 20536 35028 20588 35048
rect 20588 35028 20590 35048
rect 20534 34992 20590 35028
rect 22006 35692 22062 35728
rect 22006 35672 22008 35692
rect 22008 35672 22060 35692
rect 22060 35672 22062 35692
rect 21362 35400 21418 35456
rect 21454 34992 21510 35048
rect 19430 26832 19486 26888
rect 18694 23180 18750 23216
rect 18694 23160 18696 23180
rect 18696 23160 18748 23180
rect 18748 23160 18750 23180
rect 17130 12824 17186 12880
rect 17590 12824 17646 12880
rect 16854 10260 16910 10296
rect 16854 10240 16856 10260
rect 16856 10240 16908 10260
rect 16908 10240 16910 10260
rect 16394 6452 16450 6488
rect 16394 6432 16396 6452
rect 16396 6432 16448 6452
rect 16448 6432 16450 6452
rect 17222 10104 17278 10160
rect 18786 22616 18842 22672
rect 18694 12724 18696 12744
rect 18696 12724 18748 12744
rect 18748 12724 18750 12744
rect 18694 12688 18750 12724
rect 18510 11192 18566 11248
rect 19154 23604 19156 23624
rect 19156 23604 19208 23624
rect 19208 23604 19210 23624
rect 19154 23568 19210 23604
rect 19338 23704 19394 23760
rect 19522 23840 19578 23896
rect 20718 29028 20774 29064
rect 20718 29008 20720 29028
rect 20720 29008 20772 29028
rect 20772 29008 20774 29028
rect 20166 24928 20222 24984
rect 19890 23976 19946 24032
rect 20442 23976 20498 24032
rect 19890 22208 19946 22264
rect 19798 21664 19854 21720
rect 19522 11600 19578 11656
rect 19798 14612 19854 14648
rect 19798 14592 19800 14612
rect 19800 14592 19852 14612
rect 19852 14592 19854 14612
rect 20442 22344 20498 22400
rect 20718 26732 20720 26752
rect 20720 26732 20772 26752
rect 20772 26732 20774 26752
rect 20718 26696 20774 26732
rect 21822 32000 21878 32056
rect 21178 28500 21180 28520
rect 21180 28500 21232 28520
rect 21232 28500 21234 28520
rect 21178 28464 21234 28500
rect 21178 28192 21234 28248
rect 21086 24792 21142 24848
rect 20534 22072 20590 22128
rect 20442 20204 20444 20224
rect 20444 20204 20496 20224
rect 20496 20204 20498 20224
rect 20442 20168 20498 20204
rect 20626 20340 20628 20360
rect 20628 20340 20680 20360
rect 20680 20340 20682 20360
rect 20626 20304 20682 20340
rect 20074 19796 20076 19816
rect 20076 19796 20128 19816
rect 20128 19796 20130 19816
rect 20074 19760 20130 19796
rect 20534 19624 20590 19680
rect 20166 14492 20168 14512
rect 20168 14492 20220 14512
rect 20220 14492 20222 14512
rect 20166 14456 20222 14492
rect 19706 13096 19762 13152
rect 20442 16652 20498 16688
rect 20442 16632 20444 16652
rect 20444 16632 20496 16652
rect 20496 16632 20498 16652
rect 20810 20868 20866 20904
rect 20810 20848 20812 20868
rect 20812 20848 20864 20868
rect 20864 20848 20866 20868
rect 20810 20712 20866 20768
rect 19798 9988 19854 10024
rect 19798 9968 19800 9988
rect 19800 9968 19852 9988
rect 19852 9968 19854 9988
rect 19430 8336 19486 8392
rect 20810 16516 20866 16552
rect 20810 16496 20812 16516
rect 20812 16496 20864 16516
rect 20864 16496 20866 16516
rect 20718 13388 20774 13424
rect 20718 13368 20720 13388
rect 20720 13368 20772 13388
rect 20772 13368 20774 13388
rect 21546 29008 21602 29064
rect 21454 28328 21510 28384
rect 21362 26832 21418 26888
rect 21362 21800 21418 21856
rect 21362 21684 21418 21720
rect 21362 21664 21364 21684
rect 21364 21664 21416 21684
rect 21416 21664 21418 21684
rect 21270 19624 21326 19680
rect 21270 19372 21326 19408
rect 21270 19352 21272 19372
rect 21272 19352 21324 19372
rect 21324 19352 21326 19372
rect 21178 18672 21234 18728
rect 20074 8336 20130 8392
rect 20810 10668 20866 10704
rect 20810 10648 20812 10668
rect 20812 10648 20864 10668
rect 20864 10648 20866 10668
rect 20810 9580 20866 9616
rect 20810 9560 20812 9580
rect 20812 9560 20864 9580
rect 20864 9560 20866 9580
rect 20902 9424 20958 9480
rect 20902 9016 20958 9072
rect 20442 7656 20498 7712
rect 21822 27648 21878 27704
rect 21822 26288 21878 26344
rect 21822 23296 21878 23352
rect 21822 22344 21878 22400
rect 21914 22208 21970 22264
rect 23754 35672 23810 35728
rect 22466 35400 22522 35456
rect 22190 32428 22246 32464
rect 22190 32408 22192 32428
rect 22192 32408 22244 32428
rect 22244 32408 22246 32428
rect 22190 31764 22192 31784
rect 22192 31764 22244 31784
rect 22244 31764 22246 31784
rect 22190 31728 22246 31764
rect 22742 32272 22798 32328
rect 22374 31220 22376 31240
rect 22376 31220 22428 31240
rect 22428 31220 22430 31240
rect 22374 31184 22430 31220
rect 22374 30368 22430 30424
rect 22282 29824 22338 29880
rect 35600 41370 35656 41372
rect 35680 41370 35736 41372
rect 35760 41370 35816 41372
rect 35840 41370 35896 41372
rect 35600 41318 35646 41370
rect 35646 41318 35656 41370
rect 35680 41318 35710 41370
rect 35710 41318 35722 41370
rect 35722 41318 35736 41370
rect 35760 41318 35774 41370
rect 35774 41318 35786 41370
rect 35786 41318 35816 41370
rect 35840 41318 35850 41370
rect 35850 41318 35896 41370
rect 35600 41316 35656 41318
rect 35680 41316 35736 41318
rect 35760 41316 35816 41318
rect 35840 41316 35896 41318
rect 23846 32816 23902 32872
rect 23018 31320 23074 31376
rect 22834 29824 22890 29880
rect 22742 29588 22744 29608
rect 22744 29588 22796 29608
rect 22796 29588 22798 29608
rect 22190 26832 22246 26888
rect 22190 26560 22246 26616
rect 22190 26324 22192 26344
rect 22192 26324 22244 26344
rect 22244 26324 22246 26344
rect 22190 26288 22246 26324
rect 22742 29552 22798 29588
rect 22466 26580 22522 26616
rect 22466 26560 22468 26580
rect 22468 26560 22520 26580
rect 22520 26560 22522 26580
rect 22374 26324 22376 26344
rect 22376 26324 22428 26344
rect 22428 26324 22430 26344
rect 22374 26288 22430 26324
rect 22098 23976 22154 24032
rect 22006 21936 22062 21992
rect 21822 20576 21878 20632
rect 22650 26696 22706 26752
rect 23018 29416 23074 29472
rect 23570 29824 23626 29880
rect 23662 29280 23718 29336
rect 23202 28872 23258 28928
rect 22006 20748 22008 20768
rect 22008 20748 22060 20768
rect 22060 20748 22062 20768
rect 22006 20712 22062 20748
rect 21730 19896 21786 19952
rect 21730 19216 21786 19272
rect 21914 19352 21970 19408
rect 21822 18536 21878 18592
rect 21362 10648 21418 10704
rect 21178 9152 21234 9208
rect 21086 7404 21142 7440
rect 21086 7384 21088 7404
rect 21088 7384 21140 7404
rect 21140 7384 21142 7404
rect 19982 5908 20038 5944
rect 19982 5888 19984 5908
rect 19984 5888 20036 5908
rect 20036 5888 20038 5908
rect 22558 23840 22614 23896
rect 22742 23724 22798 23760
rect 22742 23704 22744 23724
rect 22744 23704 22796 23724
rect 22796 23704 22798 23724
rect 23846 28872 23902 28928
rect 23018 26288 23074 26344
rect 23294 25608 23350 25664
rect 23018 23840 23074 23896
rect 22466 21972 22468 21992
rect 22468 21972 22520 21992
rect 22520 21972 22522 21992
rect 22466 21936 22522 21972
rect 22006 15816 22062 15872
rect 22098 15564 22154 15600
rect 22098 15544 22100 15564
rect 22100 15544 22152 15564
rect 22152 15544 22154 15564
rect 22926 18808 22982 18864
rect 22926 17312 22982 17368
rect 22650 16768 22706 16824
rect 22926 16788 22982 16824
rect 22926 16768 22928 16788
rect 22928 16768 22980 16788
rect 22980 16768 22982 16788
rect 22190 14612 22246 14648
rect 22190 14592 22192 14612
rect 22192 14592 22244 14612
rect 22244 14592 22246 14612
rect 22374 14184 22430 14240
rect 22098 13232 22154 13288
rect 22006 13096 22062 13152
rect 22006 11872 22062 11928
rect 22282 11736 22338 11792
rect 21822 10668 21878 10704
rect 21822 10648 21824 10668
rect 21824 10648 21876 10668
rect 21876 10648 21878 10668
rect 22190 8356 22246 8392
rect 22190 8336 22192 8356
rect 22192 8336 22244 8356
rect 22244 8336 22246 8356
rect 24306 30776 24362 30832
rect 24030 29416 24086 29472
rect 24306 29416 24362 29472
rect 24490 32000 24546 32056
rect 24950 32272 25006 32328
rect 24490 29008 24546 29064
rect 24214 28484 24270 28520
rect 24214 28464 24216 28484
rect 24216 28464 24268 28484
rect 24268 28464 24270 28484
rect 23662 24792 23718 24848
rect 23478 23840 23534 23896
rect 23386 23432 23442 23488
rect 23110 20168 23166 20224
rect 23202 19932 23204 19952
rect 23204 19932 23256 19952
rect 23256 19932 23258 19952
rect 23202 19896 23258 19932
rect 23110 19488 23166 19544
rect 23386 21564 23388 21584
rect 23388 21564 23440 21584
rect 23440 21564 23442 21584
rect 23386 21528 23442 21564
rect 24674 29452 24676 29472
rect 24676 29452 24728 29472
rect 24728 29452 24730 29472
rect 24674 29416 24730 29452
rect 24858 25492 24914 25528
rect 24858 25472 24860 25492
rect 24860 25472 24912 25492
rect 24912 25472 24914 25492
rect 24030 23976 24086 24032
rect 24214 23976 24270 24032
rect 24030 22480 24086 22536
rect 23938 22208 23994 22264
rect 23754 20712 23810 20768
rect 23570 19488 23626 19544
rect 22742 13404 22744 13424
rect 22744 13404 22796 13424
rect 22796 13404 22798 13424
rect 22742 13368 22798 13404
rect 22742 12844 22798 12880
rect 22742 12824 22744 12844
rect 22744 12824 22796 12844
rect 22796 12824 22798 12844
rect 23110 11464 23166 11520
rect 22926 10512 22982 10568
rect 22834 9696 22890 9752
rect 22374 6160 22430 6216
rect 21362 5364 21418 5400
rect 21362 5344 21364 5364
rect 21364 5344 21416 5364
rect 21416 5344 21418 5364
rect 21362 3984 21418 4040
rect 23386 16496 23442 16552
rect 24030 20712 24086 20768
rect 23294 8628 23350 8664
rect 23294 8608 23296 8628
rect 23296 8608 23348 8628
rect 23348 8608 23350 8628
rect 24306 19352 24362 19408
rect 24766 24812 24822 24848
rect 25410 32272 25466 32328
rect 25042 29552 25098 29608
rect 26146 32852 26148 32872
rect 26148 32852 26200 32872
rect 26200 32852 26202 32872
rect 26146 32816 26202 32852
rect 25594 32428 25650 32464
rect 25594 32408 25596 32428
rect 25596 32408 25648 32428
rect 25648 32408 25650 32428
rect 25410 31048 25466 31104
rect 25962 30776 26018 30832
rect 25318 29588 25320 29608
rect 25320 29588 25372 29608
rect 25372 29588 25374 29608
rect 25318 29552 25374 29588
rect 25778 29824 25834 29880
rect 25594 28464 25650 28520
rect 24766 24792 24768 24812
rect 24768 24792 24820 24812
rect 24820 24792 24822 24812
rect 24398 18944 24454 19000
rect 23938 14456 23994 14512
rect 23938 14068 23994 14104
rect 24766 22072 24822 22128
rect 25134 24148 25136 24168
rect 25136 24148 25188 24168
rect 25188 24148 25190 24168
rect 25134 24112 25190 24148
rect 24858 19760 24914 19816
rect 24674 17312 24730 17368
rect 24674 15020 24730 15056
rect 24674 15000 24676 15020
rect 24676 15000 24728 15020
rect 24728 15000 24730 15020
rect 23938 14048 23940 14068
rect 23940 14048 23992 14068
rect 23992 14048 23994 14068
rect 23662 12416 23718 12472
rect 23846 12416 23902 12472
rect 24490 14068 24546 14104
rect 24490 14048 24492 14068
rect 24492 14048 24544 14068
rect 24544 14048 24546 14068
rect 24674 13948 24676 13968
rect 24676 13948 24728 13968
rect 24728 13948 24730 13968
rect 24674 13912 24730 13948
rect 24490 11872 24546 11928
rect 25410 24792 25466 24848
rect 25318 23704 25374 23760
rect 25318 20304 25374 20360
rect 26146 28500 26148 28520
rect 26148 28500 26200 28520
rect 26200 28500 26202 28520
rect 26146 28464 26202 28500
rect 25870 24148 25872 24168
rect 25872 24148 25924 24168
rect 25924 24148 25926 24168
rect 25870 24112 25926 24148
rect 25594 20576 25650 20632
rect 25042 14456 25098 14512
rect 25318 14320 25374 14376
rect 23846 8336 23902 8392
rect 24214 8916 24216 8936
rect 24216 8916 24268 8936
rect 24268 8916 24270 8936
rect 24214 8880 24270 8916
rect 24214 8608 24270 8664
rect 24122 7828 24124 7848
rect 24124 7828 24176 7848
rect 24176 7828 24178 7848
rect 24122 7792 24178 7828
rect 23846 7656 23902 7712
rect 24858 11056 24914 11112
rect 25318 11464 25374 11520
rect 25042 10648 25098 10704
rect 24766 9288 24822 9344
rect 24674 8084 24730 8120
rect 24674 8064 24676 8084
rect 24676 8064 24728 8084
rect 24728 8064 24730 8084
rect 24214 6996 24270 7032
rect 24214 6976 24216 6996
rect 24216 6976 24268 6996
rect 24268 6976 24270 6996
rect 24490 5752 24546 5808
rect 21822 3984 21878 4040
rect 22834 3848 22890 3904
rect 25410 11056 25466 11112
rect 25318 10668 25374 10704
rect 25318 10648 25320 10668
rect 25320 10648 25372 10668
rect 25372 10648 25374 10668
rect 25594 11736 25650 11792
rect 26238 24792 26294 24848
rect 27250 31764 27252 31784
rect 27252 31764 27304 31784
rect 27304 31764 27306 31784
rect 27250 31728 27306 31764
rect 26790 31592 26846 31648
rect 26422 29280 26478 29336
rect 26514 28500 26516 28520
rect 26516 28500 26568 28520
rect 26568 28500 26570 28520
rect 26514 28464 26570 28500
rect 26514 28364 26516 28384
rect 26516 28364 26568 28384
rect 26568 28364 26570 28384
rect 26514 28328 26570 28364
rect 27250 31340 27306 31376
rect 27250 31320 27252 31340
rect 27252 31320 27304 31340
rect 27304 31320 27306 31340
rect 26974 31204 27030 31240
rect 26974 31184 26976 31204
rect 26976 31184 27028 31204
rect 27028 31184 27030 31204
rect 27158 30912 27214 30968
rect 27894 31048 27950 31104
rect 27802 30912 27858 30968
rect 27342 30776 27398 30832
rect 27618 30776 27674 30832
rect 27894 29824 27950 29880
rect 26422 24248 26478 24304
rect 25962 18708 25964 18728
rect 25964 18708 26016 18728
rect 26016 18708 26018 18728
rect 25962 18672 26018 18708
rect 26054 18284 26110 18320
rect 26054 18264 26056 18284
rect 26056 18264 26108 18284
rect 26108 18264 26110 18284
rect 26698 25336 26754 25392
rect 26974 25356 27030 25392
rect 26974 25336 26976 25356
rect 26976 25336 27028 25356
rect 27028 25336 27030 25356
rect 29550 32952 29606 33008
rect 28906 32816 28962 32872
rect 29090 32272 29146 32328
rect 29366 32000 29422 32056
rect 28538 31592 28594 31648
rect 28446 31340 28502 31376
rect 28446 31320 28448 31340
rect 28448 31320 28500 31340
rect 28500 31320 28502 31340
rect 28998 30368 29054 30424
rect 27802 26324 27804 26344
rect 27804 26324 27856 26344
rect 27856 26324 27858 26344
rect 27802 26288 27858 26324
rect 27618 25064 27674 25120
rect 26146 17856 26202 17912
rect 26146 17720 26202 17776
rect 27894 26152 27950 26208
rect 28630 26152 28686 26208
rect 28170 24248 28226 24304
rect 27986 23840 28042 23896
rect 28262 23976 28318 24032
rect 28538 24248 28594 24304
rect 28814 26324 28816 26344
rect 28816 26324 28868 26344
rect 28868 26324 28870 26344
rect 28814 26288 28870 26324
rect 28446 23704 28502 23760
rect 27802 22072 27858 22128
rect 27618 20576 27674 20632
rect 27250 20304 27306 20360
rect 27066 19352 27122 19408
rect 27526 20168 27582 20224
rect 27986 21548 28042 21584
rect 27986 21528 27988 21548
rect 27988 21528 28040 21548
rect 28040 21528 28042 21548
rect 27250 18672 27306 18728
rect 27434 18572 27436 18592
rect 27436 18572 27488 18592
rect 27488 18572 27490 18592
rect 27434 18536 27490 18572
rect 27342 16632 27398 16688
rect 27710 19236 27766 19272
rect 27710 19216 27712 19236
rect 27712 19216 27764 19236
rect 27764 19216 27766 19236
rect 27618 18264 27674 18320
rect 27618 17856 27674 17912
rect 27526 16496 27582 16552
rect 26514 14184 26570 14240
rect 26238 13268 26240 13288
rect 26240 13268 26292 13288
rect 26292 13268 26294 13288
rect 26238 13232 26294 13268
rect 25594 10004 25596 10024
rect 25596 10004 25648 10024
rect 25648 10004 25650 10024
rect 25594 9968 25650 10004
rect 25502 9560 25558 9616
rect 25042 9016 25098 9072
rect 24950 8744 25006 8800
rect 26054 10804 26110 10840
rect 26054 10784 26056 10804
rect 26056 10784 26108 10804
rect 26108 10784 26110 10804
rect 27434 15000 27490 15056
rect 27066 14068 27122 14104
rect 27066 14048 27068 14068
rect 27068 14048 27120 14068
rect 27120 14048 27122 14068
rect 26882 11620 26938 11656
rect 26882 11600 26884 11620
rect 26884 11600 26936 11620
rect 26936 11600 26938 11620
rect 26514 9696 26570 9752
rect 26790 9152 26846 9208
rect 27894 17312 27950 17368
rect 28354 18536 28410 18592
rect 28998 23024 29054 23080
rect 28998 21564 29000 21584
rect 29000 21564 29052 21584
rect 29052 21564 29054 21584
rect 28998 21528 29054 21564
rect 30562 32816 30618 32872
rect 30654 31748 30710 31784
rect 30930 32680 30986 32736
rect 30654 31728 30656 31748
rect 30656 31728 30708 31748
rect 30708 31728 30710 31748
rect 30746 30912 30802 30968
rect 30746 30676 30748 30696
rect 30748 30676 30800 30696
rect 30800 30676 30802 30696
rect 30746 30640 30802 30676
rect 30470 30096 30526 30152
rect 30470 29824 30526 29880
rect 30286 29008 30342 29064
rect 29734 26696 29790 26752
rect 29366 25744 29422 25800
rect 28906 20884 28908 20904
rect 28908 20884 28960 20904
rect 28960 20884 28962 20904
rect 28906 20848 28962 20884
rect 28722 20476 28724 20496
rect 28724 20476 28776 20496
rect 28776 20476 28778 20496
rect 28722 20440 28778 20476
rect 28722 19896 28778 19952
rect 28906 18944 28962 19000
rect 28722 18708 28724 18728
rect 28724 18708 28776 18728
rect 28776 18708 28778 18728
rect 28722 18672 28778 18708
rect 28354 17312 28410 17368
rect 27802 14456 27858 14512
rect 27710 14048 27766 14104
rect 27986 14592 28042 14648
rect 28078 14356 28080 14376
rect 28080 14356 28132 14376
rect 28132 14356 28134 14376
rect 28078 14320 28134 14356
rect 27710 11464 27766 11520
rect 28078 11328 28134 11384
rect 27618 10512 27674 10568
rect 27250 9152 27306 9208
rect 27710 9172 27766 9208
rect 27710 9152 27712 9172
rect 27712 9152 27764 9172
rect 27764 9152 27766 9172
rect 27250 8336 27306 8392
rect 27158 7792 27214 7848
rect 28998 17720 29054 17776
rect 28722 17176 28778 17232
rect 28906 17176 28962 17232
rect 28630 16532 28632 16552
rect 28632 16532 28684 16552
rect 28684 16532 28686 16552
rect 28630 16496 28686 16532
rect 28814 16632 28870 16688
rect 28538 14612 28594 14648
rect 28538 14592 28540 14612
rect 28540 14592 28592 14612
rect 28592 14592 28594 14612
rect 28354 11872 28410 11928
rect 29090 15272 29146 15328
rect 28906 14492 28908 14512
rect 28908 14492 28960 14512
rect 28960 14492 28962 14512
rect 28906 14456 28962 14492
rect 28906 14356 28908 14376
rect 28908 14356 28960 14376
rect 28960 14356 28962 14376
rect 28906 14320 28962 14356
rect 28906 14048 28962 14104
rect 29274 22480 29330 22536
rect 29458 20304 29514 20360
rect 29090 13640 29146 13696
rect 28262 9424 28318 9480
rect 28906 10512 28962 10568
rect 29090 9596 29092 9616
rect 29092 9596 29144 9616
rect 29144 9596 29146 9616
rect 29090 9560 29146 9596
rect 28906 9424 28962 9480
rect 28814 8628 28870 8664
rect 28814 8608 28816 8628
rect 28816 8608 28868 8628
rect 28868 8608 28870 8628
rect 28998 8356 29054 8392
rect 28998 8336 29000 8356
rect 29000 8336 29052 8356
rect 29052 8336 29054 8356
rect 29182 7404 29238 7440
rect 29182 7384 29184 7404
rect 29184 7384 29236 7404
rect 29236 7384 29238 7404
rect 28722 5908 28778 5944
rect 28722 5888 28724 5908
rect 28724 5888 28776 5908
rect 28776 5888 28778 5908
rect 29642 23024 29698 23080
rect 30010 22480 30066 22536
rect 29918 22344 29974 22400
rect 29826 22072 29882 22128
rect 29826 20712 29882 20768
rect 29734 20476 29736 20496
rect 29736 20476 29788 20496
rect 29788 20476 29790 20496
rect 29734 20440 29790 20476
rect 29550 17720 29606 17776
rect 29550 11192 29606 11248
rect 29458 10956 29460 10976
rect 29460 10956 29512 10976
rect 29512 10956 29514 10976
rect 29458 10920 29514 10956
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 35600 40282 35656 40284
rect 35680 40282 35736 40284
rect 35760 40282 35816 40284
rect 35840 40282 35896 40284
rect 35600 40230 35646 40282
rect 35646 40230 35656 40282
rect 35680 40230 35710 40282
rect 35710 40230 35722 40282
rect 35722 40230 35736 40282
rect 35760 40230 35774 40282
rect 35774 40230 35786 40282
rect 35786 40230 35816 40282
rect 35840 40230 35850 40282
rect 35850 40230 35896 40282
rect 35600 40228 35656 40230
rect 35680 40228 35736 40230
rect 35760 40228 35816 40230
rect 35840 40228 35896 40230
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 35600 39194 35656 39196
rect 35680 39194 35736 39196
rect 35760 39194 35816 39196
rect 35840 39194 35896 39196
rect 35600 39142 35646 39194
rect 35646 39142 35656 39194
rect 35680 39142 35710 39194
rect 35710 39142 35722 39194
rect 35722 39142 35736 39194
rect 35760 39142 35774 39194
rect 35774 39142 35786 39194
rect 35786 39142 35816 39194
rect 35840 39142 35850 39194
rect 35850 39142 35896 39194
rect 35600 39140 35656 39142
rect 35680 39140 35736 39142
rect 35760 39140 35816 39142
rect 35840 39140 35896 39142
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 35600 38106 35656 38108
rect 35680 38106 35736 38108
rect 35760 38106 35816 38108
rect 35840 38106 35896 38108
rect 35600 38054 35646 38106
rect 35646 38054 35656 38106
rect 35680 38054 35710 38106
rect 35710 38054 35722 38106
rect 35722 38054 35736 38106
rect 35760 38054 35774 38106
rect 35774 38054 35786 38106
rect 35786 38054 35816 38106
rect 35840 38054 35850 38106
rect 35850 38054 35896 38106
rect 35600 38052 35656 38054
rect 35680 38052 35736 38054
rect 35760 38052 35816 38054
rect 35840 38052 35896 38054
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 31206 32952 31262 33008
rect 31022 30096 31078 30152
rect 31022 29960 31078 30016
rect 30470 26968 30526 27024
rect 30746 26988 30802 27024
rect 30746 26968 30748 26988
rect 30748 26968 30800 26988
rect 30800 26968 30802 26988
rect 31114 27376 31170 27432
rect 31022 26832 31078 26888
rect 30930 26288 30986 26344
rect 30102 19760 30158 19816
rect 29918 18708 29920 18728
rect 29920 18708 29972 18728
rect 29972 18708 29974 18728
rect 29918 18672 29974 18708
rect 30470 20884 30472 20904
rect 30472 20884 30524 20904
rect 30524 20884 30526 20904
rect 30470 20848 30526 20884
rect 32126 32020 32182 32056
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 32126 32000 32128 32020
rect 32128 32000 32180 32020
rect 32180 32000 32182 32020
rect 31390 29960 31446 30016
rect 31574 30368 31630 30424
rect 31758 30268 31760 30288
rect 31760 30268 31812 30288
rect 31812 30268 31814 30288
rect 31758 30232 31814 30268
rect 32494 32680 32550 32736
rect 32218 29960 32274 30016
rect 31022 22208 31078 22264
rect 30470 18128 30526 18184
rect 30378 16360 30434 16416
rect 30378 16224 30434 16280
rect 30286 16088 30342 16144
rect 30930 19352 30986 19408
rect 30654 16224 30710 16280
rect 30470 14356 30472 14376
rect 30472 14356 30524 14376
rect 30524 14356 30526 14376
rect 30470 14320 30526 14356
rect 30194 12960 30250 13016
rect 29734 12724 29736 12744
rect 29736 12724 29788 12744
rect 29788 12724 29790 12744
rect 29734 12688 29790 12724
rect 29734 12280 29790 12336
rect 30470 12688 30526 12744
rect 30470 12416 30526 12472
rect 29550 10124 29606 10160
rect 29550 10104 29552 10124
rect 29552 10104 29604 10124
rect 29604 10104 29606 10124
rect 29734 9016 29790 9072
rect 29734 8608 29790 8664
rect 29550 7520 29606 7576
rect 32494 30096 32550 30152
rect 31666 26288 31722 26344
rect 31850 26324 31852 26344
rect 31852 26324 31904 26344
rect 31904 26324 31906 26344
rect 31850 26288 31906 26324
rect 31942 25336 31998 25392
rect 31850 22772 31906 22808
rect 31850 22752 31852 22772
rect 31852 22752 31904 22772
rect 31904 22752 31906 22772
rect 31850 22344 31906 22400
rect 31758 20476 31760 20496
rect 31760 20476 31812 20496
rect 31812 20476 31814 20496
rect 31758 20440 31814 20476
rect 31298 17448 31354 17504
rect 30838 12960 30894 13016
rect 30930 11192 30986 11248
rect 30378 8472 30434 8528
rect 31574 16632 31630 16688
rect 31206 15444 31208 15464
rect 31208 15444 31260 15464
rect 31260 15444 31262 15464
rect 31206 15408 31262 15444
rect 31482 15408 31538 15464
rect 31206 10512 31262 10568
rect 30838 9696 30894 9752
rect 31114 9016 31170 9072
rect 31850 17856 31906 17912
rect 32310 26968 32366 27024
rect 32494 26832 32550 26888
rect 32310 26560 32366 26616
rect 32494 26560 32550 26616
rect 32494 26324 32496 26344
rect 32496 26324 32548 26344
rect 32548 26324 32550 26344
rect 32494 26288 32550 26324
rect 32494 24928 32550 24984
rect 32402 24792 32458 24848
rect 32310 23604 32312 23624
rect 32312 23604 32364 23624
rect 32364 23604 32366 23624
rect 32310 23568 32366 23604
rect 31850 13504 31906 13560
rect 31574 10512 31630 10568
rect 31574 9288 31630 9344
rect 32218 13640 32274 13696
rect 32770 27512 32826 27568
rect 32770 27276 32772 27296
rect 32772 27276 32824 27296
rect 32824 27276 32826 27296
rect 32770 27240 32826 27276
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 35806 32816 35862 32872
rect 33506 30232 33562 30288
rect 33414 30116 33470 30152
rect 33414 30096 33416 30116
rect 33416 30096 33468 30116
rect 33468 30096 33470 30116
rect 33414 29688 33470 29744
rect 33690 30368 33746 30424
rect 33874 30676 33876 30696
rect 33876 30676 33928 30696
rect 33928 30676 33930 30696
rect 33874 30640 33930 30676
rect 33874 29688 33930 29744
rect 34610 32680 34666 32736
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 34794 32272 34850 32328
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 34610 30912 34666 30968
rect 34058 29824 34114 29880
rect 33966 29416 34022 29472
rect 33506 29280 33562 29336
rect 33690 29164 33746 29200
rect 33690 29144 33692 29164
rect 33692 29144 33744 29164
rect 33744 29144 33746 29164
rect 33874 29144 33930 29200
rect 33506 29008 33562 29064
rect 33230 26696 33286 26752
rect 33138 23724 33194 23760
rect 33138 23704 33140 23724
rect 33140 23704 33192 23724
rect 33192 23704 33194 23724
rect 33230 23180 33286 23216
rect 33230 23160 33232 23180
rect 33232 23160 33284 23180
rect 33284 23160 33286 23180
rect 33598 26460 33600 26480
rect 33600 26460 33652 26480
rect 33652 26460 33654 26480
rect 33598 26424 33654 26460
rect 33690 25236 33692 25256
rect 33692 25236 33744 25256
rect 33744 25236 33746 25256
rect 33690 25200 33746 25236
rect 34150 29452 34152 29472
rect 34152 29452 34204 29472
rect 34204 29452 34206 29472
rect 34150 29416 34206 29452
rect 32770 17584 32826 17640
rect 32586 16632 32642 16688
rect 32402 13368 32458 13424
rect 32126 9580 32182 9616
rect 32126 9560 32128 9580
rect 32128 9560 32180 9580
rect 32180 9560 32182 9580
rect 33506 22344 33562 22400
rect 32862 11092 32864 11112
rect 32864 11092 32916 11112
rect 32916 11092 32918 11112
rect 32862 11056 32918 11092
rect 34610 29164 34666 29200
rect 34610 29144 34612 29164
rect 34612 29144 34664 29164
rect 34664 29144 34666 29164
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 33598 17060 33654 17096
rect 33598 17040 33600 17060
rect 33600 17040 33652 17060
rect 33652 17040 33654 17060
rect 33506 12144 33562 12200
rect 33690 12824 33746 12880
rect 35070 29416 35126 29472
rect 34978 29280 35034 29336
rect 35622 29572 35678 29608
rect 35622 29552 35624 29572
rect 35624 29552 35676 29572
rect 35676 29552 35678 29572
rect 36358 30504 36414 30560
rect 36542 30096 36598 30152
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 34702 28872 34758 28928
rect 34702 26152 34758 26208
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35162 26152 35218 26208
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 35254 24656 35310 24712
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34886 23724 34942 23760
rect 34886 23704 34888 23724
rect 34888 23704 34940 23724
rect 34940 23704 34942 23724
rect 34794 23604 34796 23624
rect 34796 23604 34848 23624
rect 34848 23604 34850 23624
rect 34794 23568 34850 23604
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 35254 22752 35310 22808
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34610 20712 34666 20768
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 35714 29144 35770 29200
rect 36082 29164 36138 29200
rect 36082 29144 36084 29164
rect 36084 29144 36136 29164
rect 36136 29144 36138 29164
rect 36634 29708 36690 29744
rect 36634 29688 36636 29708
rect 36636 29688 36688 29708
rect 36688 29688 36690 29708
rect 36818 29824 36874 29880
rect 36910 29552 36966 29608
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 35622 26832 35678 26888
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 35530 25236 35532 25256
rect 35532 25236 35584 25256
rect 35584 25236 35586 25256
rect 35530 25200 35586 25236
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 36818 25356 36874 25392
rect 36818 25336 36820 25356
rect 36820 25336 36872 25356
rect 36872 25336 36874 25356
rect 36174 22636 36230 22672
rect 36174 22616 36176 22636
rect 36176 22616 36228 22636
rect 36228 22616 36230 22636
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 34702 19352 34758 19408
rect 34426 18300 34428 18320
rect 34428 18300 34480 18320
rect 34480 18300 34482 18320
rect 34426 18264 34482 18300
rect 34426 16124 34428 16144
rect 34428 16124 34480 16144
rect 34480 16124 34482 16144
rect 34426 16088 34482 16124
rect 33598 11756 33654 11792
rect 33598 11736 33600 11756
rect 33600 11736 33652 11756
rect 33652 11736 33654 11756
rect 33598 11056 33654 11112
rect 34334 11736 34390 11792
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 35530 19352 35586 19408
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 35898 19216 35954 19272
rect 35898 18808 35954 18864
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 34886 17584 34942 17640
rect 35346 17448 35402 17504
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 36450 23060 36452 23080
rect 36452 23060 36504 23080
rect 36504 23060 36506 23080
rect 36450 23024 36506 23060
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35162 16124 35164 16144
rect 35164 16124 35216 16144
rect 35216 16124 35218 16144
rect 35162 16088 35218 16124
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34702 13096 34758 13152
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34794 11736 34850 11792
rect 34242 8880 34298 8936
rect 33506 7948 33562 7984
rect 33506 7928 33508 7948
rect 33508 7928 33560 7948
rect 33560 7928 33562 7948
rect 29550 6296 29606 6352
rect 29182 5228 29238 5264
rect 34518 9580 34574 9616
rect 34518 9560 34520 9580
rect 34520 9560 34572 9580
rect 34572 9560 34574 9580
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34978 11192 35034 11248
rect 34886 10956 34888 10976
rect 34888 10956 34940 10976
rect 34940 10956 34942 10976
rect 34886 10920 34942 10956
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 35070 9696 35126 9752
rect 34334 8336 34390 8392
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 37738 29028 37794 29064
rect 37738 29008 37740 29028
rect 37740 29008 37792 29028
rect 37792 29008 37794 29028
rect 37094 27104 37150 27160
rect 37370 27412 37372 27432
rect 37372 27412 37424 27432
rect 37424 27412 37426 27432
rect 37370 27376 37426 27412
rect 37278 23432 37334 23488
rect 38566 31320 38622 31376
rect 38106 26968 38162 27024
rect 38382 26308 38438 26344
rect 38382 26288 38384 26308
rect 38384 26288 38436 26308
rect 38436 26288 38438 26308
rect 38198 24792 38254 24848
rect 36818 16496 36874 16552
rect 37186 19780 37242 19816
rect 37186 19760 37188 19780
rect 37188 19760 37240 19780
rect 37240 19760 37242 19780
rect 36910 15272 36966 15328
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 35346 9016 35402 9072
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 35990 9580 36046 9616
rect 35990 9560 35992 9580
rect 35992 9560 36044 9580
rect 36044 9560 36046 9580
rect 36818 11600 36874 11656
rect 36634 11092 36636 11112
rect 36636 11092 36688 11112
rect 36688 11092 36690 11112
rect 36634 11056 36690 11092
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 37278 17720 37334 17776
rect 37278 16360 37334 16416
rect 38014 23024 38070 23080
rect 38014 22480 38070 22536
rect 38106 20984 38162 21040
rect 38106 19896 38162 19952
rect 38750 23160 38806 23216
rect 38290 18672 38346 18728
rect 38290 17992 38346 18048
rect 38198 12144 38254 12200
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 37738 8492 37794 8528
rect 37738 8472 37740 8492
rect 37740 8472 37792 8492
rect 37792 8472 37794 8492
rect 39578 27240 39634 27296
rect 39670 23840 39726 23896
rect 39394 17720 39450 17776
rect 38014 9172 38070 9208
rect 38014 9152 38016 9172
rect 38016 9152 38068 9172
rect 38068 9152 38070 9172
rect 39946 25880 40002 25936
rect 40222 26560 40278 26616
rect 40222 24520 40278 24576
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 29182 5208 29184 5228
rect 29184 5208 29236 5228
rect 29236 5208 29238 5228
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 40130 3460 40186 3496
rect 40130 3440 40132 3460
rect 40132 3440 40184 3460
rect 40184 3440 40186 3460
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
<< metal3 >>
rect 4870 41376 5186 41377
rect 4870 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5186 41376
rect 4870 41311 5186 41312
rect 35590 41376 35906 41377
rect 35590 41312 35596 41376
rect 35660 41312 35676 41376
rect 35740 41312 35756 41376
rect 35820 41312 35836 41376
rect 35900 41312 35906 41376
rect 35590 41311 35906 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 4870 40288 5186 40289
rect 4870 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5186 40288
rect 4870 40223 5186 40224
rect 35590 40288 35906 40289
rect 35590 40224 35596 40288
rect 35660 40224 35676 40288
rect 35740 40224 35756 40288
rect 35820 40224 35836 40288
rect 35900 40224 35906 40288
rect 35590 40223 35906 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 4870 39200 5186 39201
rect 4870 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5186 39200
rect 4870 39135 5186 39136
rect 35590 39200 35906 39201
rect 35590 39136 35596 39200
rect 35660 39136 35676 39200
rect 35740 39136 35756 39200
rect 35820 39136 35836 39200
rect 35900 39136 35906 39200
rect 35590 39135 35906 39136
rect 0 38858 800 38888
rect 3417 38858 3483 38861
rect 0 38856 3483 38858
rect 0 38800 3422 38856
rect 3478 38800 3483 38856
rect 0 38798 3483 38800
rect 0 38768 800 38798
rect 3417 38795 3483 38798
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 8017 38314 8083 38317
rect 8845 38314 8911 38317
rect 9029 38314 9095 38317
rect 8017 38312 9095 38314
rect 8017 38256 8022 38312
rect 8078 38256 8850 38312
rect 8906 38256 9034 38312
rect 9090 38256 9095 38312
rect 8017 38254 9095 38256
rect 8017 38251 8083 38254
rect 8845 38251 8911 38254
rect 9029 38251 9095 38254
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 35590 38112 35906 38113
rect 35590 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35906 38112
rect 35590 38047 35906 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 14181 36274 14247 36277
rect 15837 36274 15903 36277
rect 14181 36272 15903 36274
rect 14181 36216 14186 36272
rect 14242 36216 15842 36272
rect 15898 36216 15903 36272
rect 14181 36214 15903 36216
rect 14181 36211 14247 36214
rect 15837 36211 15903 36214
rect 0 36138 800 36168
rect 2957 36138 3023 36141
rect 0 36136 3023 36138
rect 0 36080 2962 36136
rect 3018 36080 3023 36136
rect 0 36078 3023 36080
rect 0 36048 800 36078
rect 2957 36075 3023 36078
rect 7281 36138 7347 36141
rect 9121 36138 9187 36141
rect 7281 36136 9187 36138
rect 7281 36080 7286 36136
rect 7342 36080 9126 36136
rect 9182 36080 9187 36136
rect 7281 36078 9187 36080
rect 7281 36075 7347 36078
rect 9121 36075 9187 36078
rect 10133 36002 10199 36005
rect 11053 36002 11119 36005
rect 10133 36000 11119 36002
rect 10133 35944 10138 36000
rect 10194 35944 11058 36000
rect 11114 35944 11119 36000
rect 10133 35942 11119 35944
rect 10133 35939 10199 35942
rect 11053 35939 11119 35942
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 10501 35730 10567 35733
rect 10961 35730 11027 35733
rect 10501 35728 11027 35730
rect 10501 35672 10506 35728
rect 10562 35672 10966 35728
rect 11022 35672 11027 35728
rect 10501 35670 11027 35672
rect 10501 35667 10567 35670
rect 10961 35667 11027 35670
rect 22001 35730 22067 35733
rect 23749 35730 23815 35733
rect 22001 35728 23815 35730
rect 22001 35672 22006 35728
rect 22062 35672 23754 35728
rect 23810 35672 23815 35728
rect 22001 35670 23815 35672
rect 22001 35667 22067 35670
rect 23749 35667 23815 35670
rect 17493 35594 17559 35597
rect 18045 35594 18111 35597
rect 17493 35592 18111 35594
rect 17493 35536 17498 35592
rect 17554 35536 18050 35592
rect 18106 35536 18111 35592
rect 17493 35534 18111 35536
rect 17493 35531 17559 35534
rect 18045 35531 18111 35534
rect 21357 35458 21423 35461
rect 22461 35458 22527 35461
rect 21357 35456 22527 35458
rect 21357 35400 21362 35456
rect 21418 35400 22466 35456
rect 22522 35400 22527 35456
rect 21357 35398 22527 35400
rect 21357 35395 21423 35398
rect 22461 35395 22527 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 6269 35322 6335 35325
rect 7557 35322 7623 35325
rect 8150 35322 8156 35324
rect 6269 35320 8156 35322
rect 6269 35264 6274 35320
rect 6330 35264 7562 35320
rect 7618 35264 8156 35320
rect 6269 35262 8156 35264
rect 6269 35259 6335 35262
rect 7557 35259 7623 35262
rect 8150 35260 8156 35262
rect 8220 35260 8226 35324
rect 6453 35186 6519 35189
rect 7373 35186 7439 35189
rect 6453 35184 7439 35186
rect 6453 35128 6458 35184
rect 6514 35128 7378 35184
rect 7434 35128 7439 35184
rect 6453 35126 7439 35128
rect 6453 35123 6519 35126
rect 7373 35123 7439 35126
rect 10133 35050 10199 35053
rect 12893 35050 12959 35053
rect 18689 35050 18755 35053
rect 10133 35048 18755 35050
rect 10133 34992 10138 35048
rect 10194 34992 12898 35048
rect 12954 34992 18694 35048
rect 18750 34992 18755 35048
rect 10133 34990 18755 34992
rect 10133 34987 10199 34990
rect 12893 34987 12959 34990
rect 18689 34987 18755 34990
rect 20529 35050 20595 35053
rect 21449 35050 21515 35053
rect 20529 35048 21515 35050
rect 20529 34992 20534 35048
rect 20590 34992 21454 35048
rect 21510 34992 21515 35048
rect 20529 34990 21515 34992
rect 20529 34987 20595 34990
rect 21449 34987 21515 34990
rect 4870 34848 5186 34849
rect 0 34778 800 34808
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 1301 34778 1367 34781
rect 0 34776 1367 34778
rect 0 34720 1306 34776
rect 1362 34720 1367 34776
rect 0 34718 1367 34720
rect 0 34688 800 34718
rect 1301 34715 1367 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 0 34098 800 34128
rect 1669 34098 1735 34101
rect 0 34096 1735 34098
rect 0 34040 1674 34096
rect 1730 34040 1735 34096
rect 0 34038 1735 34040
rect 0 34008 800 34038
rect 1669 34035 1735 34038
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 0 33418 800 33448
rect 1669 33418 1735 33421
rect 0 33416 1735 33418
rect 0 33360 1674 33416
rect 1730 33360 1735 33416
rect 0 33358 1735 33360
rect 0 33328 800 33358
rect 1669 33355 1735 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 15561 33010 15627 33013
rect 16481 33010 16547 33013
rect 22502 33010 22508 33012
rect 15561 33008 22508 33010
rect 15561 32952 15566 33008
rect 15622 32952 16486 33008
rect 16542 32952 22508 33008
rect 15561 32950 22508 32952
rect 15561 32947 15627 32950
rect 16481 32947 16547 32950
rect 22502 32948 22508 32950
rect 22572 32948 22578 33012
rect 29545 33010 29611 33013
rect 30414 33010 30420 33012
rect 29545 33008 30420 33010
rect 29545 32952 29550 33008
rect 29606 32952 30420 33008
rect 29545 32950 30420 32952
rect 29545 32947 29611 32950
rect 30414 32948 30420 32950
rect 30484 33010 30490 33012
rect 31201 33010 31267 33013
rect 30484 33008 31267 33010
rect 30484 32952 31206 33008
rect 31262 32952 31267 33008
rect 30484 32950 31267 32952
rect 30484 32948 30490 32950
rect 31201 32947 31267 32950
rect 23841 32874 23907 32877
rect 26141 32874 26207 32877
rect 28901 32874 28967 32877
rect 23841 32872 28967 32874
rect 23841 32816 23846 32872
rect 23902 32816 26146 32872
rect 26202 32816 28906 32872
rect 28962 32816 28967 32872
rect 23841 32814 28967 32816
rect 23841 32811 23907 32814
rect 26141 32811 26207 32814
rect 28901 32811 28967 32814
rect 30557 32874 30623 32877
rect 35801 32874 35867 32877
rect 30557 32872 35867 32874
rect 30557 32816 30562 32872
rect 30618 32816 35806 32872
rect 35862 32816 35867 32872
rect 30557 32814 35867 32816
rect 30557 32811 30623 32814
rect 35801 32811 35867 32814
rect 0 32738 800 32768
rect 1485 32738 1551 32741
rect 0 32736 1551 32738
rect 0 32680 1490 32736
rect 1546 32680 1551 32736
rect 0 32678 1551 32680
rect 0 32648 800 32678
rect 1485 32675 1551 32678
rect 30925 32738 30991 32741
rect 32489 32738 32555 32741
rect 34605 32738 34671 32741
rect 30925 32736 34671 32738
rect 30925 32680 30930 32736
rect 30986 32680 32494 32736
rect 32550 32680 34610 32736
rect 34666 32680 34671 32736
rect 30925 32678 34671 32680
rect 30925 32675 30991 32678
rect 32489 32675 32555 32678
rect 34605 32675 34671 32678
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 35590 32607 35906 32608
rect 8477 32602 8543 32605
rect 9806 32602 9812 32604
rect 8477 32600 9812 32602
rect 8477 32544 8482 32600
rect 8538 32544 9812 32600
rect 8477 32542 9812 32544
rect 8477 32539 8543 32542
rect 9806 32540 9812 32542
rect 9876 32540 9882 32604
rect 22185 32466 22251 32469
rect 25589 32466 25655 32469
rect 22185 32464 25655 32466
rect 22185 32408 22190 32464
rect 22246 32408 25594 32464
rect 25650 32408 25655 32464
rect 22185 32406 25655 32408
rect 22185 32403 22251 32406
rect 25589 32403 25655 32406
rect 22737 32330 22803 32333
rect 24945 32330 25011 32333
rect 25405 32330 25471 32333
rect 22737 32328 25471 32330
rect 22737 32272 22742 32328
rect 22798 32272 24950 32328
rect 25006 32272 25410 32328
rect 25466 32272 25471 32328
rect 22737 32270 25471 32272
rect 22737 32267 22803 32270
rect 24945 32267 25011 32270
rect 25405 32267 25471 32270
rect 29085 32330 29151 32333
rect 34789 32330 34855 32333
rect 29085 32328 34855 32330
rect 29085 32272 29090 32328
rect 29146 32272 34794 32328
rect 34850 32272 34855 32328
rect 29085 32270 34855 32272
rect 29085 32267 29151 32270
rect 34789 32267 34855 32270
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 18454 31996 18460 32060
rect 18524 32058 18530 32060
rect 21817 32058 21883 32061
rect 18524 32056 21883 32058
rect 18524 32000 21822 32056
rect 21878 32000 21883 32056
rect 18524 31998 21883 32000
rect 18524 31996 18530 31998
rect 21817 31995 21883 31998
rect 24485 32060 24551 32061
rect 24485 32056 24532 32060
rect 24596 32058 24602 32060
rect 29361 32058 29427 32061
rect 32121 32058 32187 32061
rect 24485 32000 24490 32056
rect 24485 31996 24532 32000
rect 24596 31998 24642 32058
rect 29361 32056 32187 32058
rect 29361 32000 29366 32056
rect 29422 32000 32126 32056
rect 32182 32000 32187 32056
rect 29361 31998 32187 32000
rect 24596 31996 24602 31998
rect 24485 31995 24551 31996
rect 29361 31995 29427 31998
rect 32121 31995 32187 31998
rect 10961 31786 11027 31789
rect 12249 31786 12315 31789
rect 10961 31784 12315 31786
rect 10961 31728 10966 31784
rect 11022 31728 12254 31784
rect 12310 31728 12315 31784
rect 10961 31726 12315 31728
rect 10961 31723 11027 31726
rect 12249 31723 12315 31726
rect 13670 31724 13676 31788
rect 13740 31786 13746 31788
rect 16113 31786 16179 31789
rect 13740 31784 16179 31786
rect 13740 31728 16118 31784
rect 16174 31728 16179 31784
rect 13740 31726 16179 31728
rect 13740 31724 13746 31726
rect 16113 31723 16179 31726
rect 22185 31786 22251 31789
rect 27245 31786 27311 31789
rect 30649 31788 30715 31789
rect 27470 31786 27476 31788
rect 22185 31784 27476 31786
rect 22185 31728 22190 31784
rect 22246 31728 27250 31784
rect 27306 31728 27476 31784
rect 22185 31726 27476 31728
rect 22185 31723 22251 31726
rect 27245 31723 27311 31726
rect 27470 31724 27476 31726
rect 27540 31724 27546 31788
rect 30598 31786 30604 31788
rect 30558 31726 30604 31786
rect 30668 31784 30715 31788
rect 30710 31728 30715 31784
rect 30598 31724 30604 31726
rect 30668 31724 30715 31728
rect 30649 31723 30715 31724
rect 11145 31650 11211 31653
rect 12014 31650 12020 31652
rect 11145 31648 12020 31650
rect 11145 31592 11150 31648
rect 11206 31592 12020 31648
rect 11145 31590 12020 31592
rect 11145 31587 11211 31590
rect 12014 31588 12020 31590
rect 12084 31650 12090 31652
rect 12249 31650 12315 31653
rect 12084 31648 12315 31650
rect 12084 31592 12254 31648
rect 12310 31592 12315 31648
rect 12084 31590 12315 31592
rect 12084 31588 12090 31590
rect 12249 31587 12315 31590
rect 26785 31650 26851 31653
rect 28533 31650 28599 31653
rect 26785 31648 28599 31650
rect 26785 31592 26790 31648
rect 26846 31592 28538 31648
rect 28594 31592 28599 31648
rect 26785 31590 28599 31592
rect 26785 31587 26851 31590
rect 28533 31587 28599 31590
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 0 31378 800 31408
rect 3233 31378 3299 31381
rect 0 31376 3299 31378
rect 0 31320 3238 31376
rect 3294 31320 3299 31376
rect 0 31318 3299 31320
rect 0 31288 800 31318
rect 3233 31315 3299 31318
rect 23013 31378 23079 31381
rect 24894 31378 24900 31380
rect 23013 31376 24900 31378
rect 23013 31320 23018 31376
rect 23074 31320 24900 31376
rect 23013 31318 24900 31320
rect 23013 31315 23079 31318
rect 24894 31316 24900 31318
rect 24964 31316 24970 31380
rect 27245 31378 27311 31381
rect 28441 31378 28507 31381
rect 38561 31378 38627 31381
rect 27245 31376 38627 31378
rect 27245 31320 27250 31376
rect 27306 31320 28446 31376
rect 28502 31320 38566 31376
rect 38622 31320 38627 31376
rect 27245 31318 38627 31320
rect 27245 31315 27311 31318
rect 28441 31315 28507 31318
rect 38561 31315 38627 31318
rect 22369 31242 22435 31245
rect 26969 31242 27035 31245
rect 22369 31240 27035 31242
rect 22369 31184 22374 31240
rect 22430 31184 26974 31240
rect 27030 31184 27035 31240
rect 22369 31182 27035 31184
rect 22369 31179 22435 31182
rect 26969 31179 27035 31182
rect 25405 31106 25471 31109
rect 27889 31106 27955 31109
rect 25405 31104 27955 31106
rect 25405 31048 25410 31104
rect 25466 31048 27894 31104
rect 27950 31048 27955 31104
rect 25405 31046 27955 31048
rect 25405 31043 25471 31046
rect 27889 31043 27955 31046
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 27153 30970 27219 30973
rect 27797 30970 27863 30973
rect 27153 30968 27863 30970
rect 27153 30912 27158 30968
rect 27214 30912 27802 30968
rect 27858 30912 27863 30968
rect 27153 30910 27863 30912
rect 27153 30907 27219 30910
rect 27797 30907 27863 30910
rect 30741 30970 30807 30973
rect 34605 30972 34671 30973
rect 34605 30970 34652 30972
rect 30741 30968 34652 30970
rect 34716 30970 34722 30972
rect 30741 30912 30746 30968
rect 30802 30912 34610 30968
rect 30741 30910 34652 30912
rect 30741 30907 30807 30910
rect 34605 30908 34652 30910
rect 34716 30910 34798 30970
rect 34716 30908 34722 30910
rect 34605 30907 34671 30908
rect 4797 30834 4863 30837
rect 24301 30834 24367 30837
rect 4797 30832 24367 30834
rect 4797 30776 4802 30832
rect 4858 30776 24306 30832
rect 24362 30776 24367 30832
rect 4797 30774 24367 30776
rect 4797 30771 4863 30774
rect 24301 30771 24367 30774
rect 25957 30834 26023 30837
rect 27337 30834 27403 30837
rect 27613 30834 27679 30837
rect 25957 30832 27679 30834
rect 25957 30776 25962 30832
rect 26018 30776 27342 30832
rect 27398 30776 27618 30832
rect 27674 30776 27679 30832
rect 25957 30774 27679 30776
rect 25957 30771 26023 30774
rect 27337 30771 27403 30774
rect 27613 30771 27679 30774
rect 0 30698 800 30728
rect 1577 30698 1643 30701
rect 0 30696 1643 30698
rect 0 30640 1582 30696
rect 1638 30640 1643 30696
rect 0 30638 1643 30640
rect 0 30608 800 30638
rect 1577 30635 1643 30638
rect 14825 30698 14891 30701
rect 15561 30698 15627 30701
rect 14825 30696 15627 30698
rect 14825 30640 14830 30696
rect 14886 30640 15566 30696
rect 15622 30640 15627 30696
rect 14825 30638 15627 30640
rect 14825 30635 14891 30638
rect 15561 30635 15627 30638
rect 30741 30698 30807 30701
rect 33869 30698 33935 30701
rect 30741 30696 33935 30698
rect 30741 30640 30746 30696
rect 30802 30640 33874 30696
rect 33930 30640 33935 30696
rect 30741 30638 33935 30640
rect 30741 30635 30807 30638
rect 33869 30635 33935 30638
rect 36118 30500 36124 30564
rect 36188 30562 36194 30564
rect 36353 30562 36419 30565
rect 36188 30560 36419 30562
rect 36188 30504 36358 30560
rect 36414 30504 36419 30560
rect 36188 30502 36419 30504
rect 36188 30500 36194 30502
rect 36353 30499 36419 30502
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 22134 30364 22140 30428
rect 22204 30426 22210 30428
rect 22369 30426 22435 30429
rect 22204 30424 22435 30426
rect 22204 30368 22374 30424
rect 22430 30368 22435 30424
rect 22204 30366 22435 30368
rect 22204 30364 22210 30366
rect 22369 30363 22435 30366
rect 28993 30426 29059 30429
rect 29678 30426 29684 30428
rect 28993 30424 29684 30426
rect 28993 30368 28998 30424
rect 29054 30368 29684 30424
rect 28993 30366 29684 30368
rect 28993 30363 29059 30366
rect 29678 30364 29684 30366
rect 29748 30364 29754 30428
rect 31569 30426 31635 30429
rect 33685 30426 33751 30429
rect 31569 30424 33751 30426
rect 31569 30368 31574 30424
rect 31630 30368 33690 30424
rect 33746 30368 33751 30424
rect 31569 30366 33751 30368
rect 31569 30363 31635 30366
rect 33685 30363 33751 30366
rect 31753 30290 31819 30293
rect 33501 30290 33567 30293
rect 31753 30288 33567 30290
rect 31753 30232 31758 30288
rect 31814 30232 33506 30288
rect 33562 30232 33567 30288
rect 31753 30230 33567 30232
rect 31753 30227 31819 30230
rect 33501 30227 33567 30230
rect 841 30154 907 30157
rect 798 30152 907 30154
rect 798 30096 846 30152
rect 902 30096 907 30152
rect 798 30091 907 30096
rect 15653 30154 15719 30157
rect 16021 30154 16087 30157
rect 15653 30152 16087 30154
rect 15653 30096 15658 30152
rect 15714 30096 16026 30152
rect 16082 30096 16087 30152
rect 15653 30094 16087 30096
rect 15653 30091 15719 30094
rect 16021 30091 16087 30094
rect 30465 30154 30531 30157
rect 31017 30154 31083 30157
rect 32489 30154 32555 30157
rect 30465 30152 32555 30154
rect 30465 30096 30470 30152
rect 30526 30096 31022 30152
rect 31078 30096 32494 30152
rect 32550 30096 32555 30152
rect 30465 30094 32555 30096
rect 30465 30091 30531 30094
rect 31017 30091 31083 30094
rect 32489 30091 32555 30094
rect 33409 30154 33475 30157
rect 36537 30154 36603 30157
rect 33409 30152 36603 30154
rect 33409 30096 33414 30152
rect 33470 30096 36542 30152
rect 36598 30096 36603 30152
rect 33409 30094 36603 30096
rect 33409 30091 33475 30094
rect 36537 30091 36603 30094
rect 798 30048 858 30091
rect 0 29958 858 30048
rect 14641 30018 14707 30021
rect 18321 30018 18387 30021
rect 14641 30016 18387 30018
rect 14641 29960 14646 30016
rect 14702 29960 18326 30016
rect 18382 29960 18387 30016
rect 14641 29958 18387 29960
rect 0 29928 800 29958
rect 14641 29955 14707 29958
rect 18321 29955 18387 29958
rect 31017 30018 31083 30021
rect 31385 30018 31451 30021
rect 32213 30018 32279 30021
rect 31017 30016 32279 30018
rect 31017 29960 31022 30016
rect 31078 29960 31390 30016
rect 31446 29960 32218 30016
rect 32274 29960 32279 30016
rect 31017 29958 32279 29960
rect 31017 29955 31083 29958
rect 31385 29955 31451 29958
rect 32213 29955 32279 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 22277 29882 22343 29885
rect 22829 29882 22895 29885
rect 23565 29882 23631 29885
rect 22277 29880 23631 29882
rect 22277 29824 22282 29880
rect 22338 29824 22834 29880
rect 22890 29824 23570 29880
rect 23626 29824 23631 29880
rect 22277 29822 23631 29824
rect 22277 29819 22343 29822
rect 22829 29819 22895 29822
rect 23565 29819 23631 29822
rect 25773 29882 25839 29885
rect 27889 29882 27955 29885
rect 30465 29884 30531 29885
rect 30414 29882 30420 29884
rect 25773 29880 27955 29882
rect 25773 29824 25778 29880
rect 25834 29824 27894 29880
rect 27950 29824 27955 29880
rect 25773 29822 27955 29824
rect 30374 29822 30420 29882
rect 30484 29882 30531 29884
rect 34053 29882 34119 29885
rect 30484 29880 34119 29882
rect 30526 29824 34058 29880
rect 34114 29824 34119 29880
rect 25773 29819 25839 29822
rect 27889 29819 27955 29822
rect 30414 29820 30420 29822
rect 30484 29822 34119 29824
rect 30484 29820 30531 29822
rect 30465 29819 30531 29820
rect 34053 29819 34119 29822
rect 35382 29820 35388 29884
rect 35452 29882 35458 29884
rect 36813 29882 36879 29885
rect 35452 29880 36879 29882
rect 35452 29824 36818 29880
rect 36874 29824 36879 29880
rect 35452 29822 36879 29824
rect 35452 29820 35458 29822
rect 36813 29819 36879 29822
rect 10777 29746 10843 29749
rect 14733 29746 14799 29749
rect 10777 29744 14799 29746
rect 10777 29688 10782 29744
rect 10838 29688 14738 29744
rect 14794 29688 14799 29744
rect 10777 29686 14799 29688
rect 10777 29683 10843 29686
rect 14733 29683 14799 29686
rect 15469 29746 15535 29749
rect 16297 29746 16363 29749
rect 33409 29746 33475 29749
rect 15469 29744 33475 29746
rect 15469 29688 15474 29744
rect 15530 29688 16302 29744
rect 16358 29688 33414 29744
rect 33470 29688 33475 29744
rect 15469 29686 33475 29688
rect 15469 29683 15535 29686
rect 16297 29683 16363 29686
rect 33409 29683 33475 29686
rect 33869 29746 33935 29749
rect 36629 29746 36695 29749
rect 33869 29744 36695 29746
rect 33869 29688 33874 29744
rect 33930 29688 36634 29744
rect 36690 29688 36695 29744
rect 33869 29686 36695 29688
rect 33869 29683 33935 29686
rect 36629 29683 36695 29686
rect 10685 29610 10751 29613
rect 11697 29610 11763 29613
rect 10685 29608 11763 29610
rect 10685 29552 10690 29608
rect 10746 29552 11702 29608
rect 11758 29552 11763 29608
rect 10685 29550 11763 29552
rect 10685 29547 10751 29550
rect 11697 29547 11763 29550
rect 13077 29610 13143 29613
rect 13353 29610 13419 29613
rect 18597 29610 18663 29613
rect 13077 29608 18663 29610
rect 13077 29552 13082 29608
rect 13138 29552 13358 29608
rect 13414 29552 18602 29608
rect 18658 29552 18663 29608
rect 13077 29550 18663 29552
rect 13077 29547 13143 29550
rect 13353 29547 13419 29550
rect 18597 29547 18663 29550
rect 22737 29610 22803 29613
rect 25037 29610 25103 29613
rect 25313 29610 25379 29613
rect 22737 29608 25379 29610
rect 22737 29552 22742 29608
rect 22798 29552 25042 29608
rect 25098 29552 25318 29608
rect 25374 29552 25379 29608
rect 22737 29550 25379 29552
rect 22737 29547 22803 29550
rect 25037 29547 25103 29550
rect 25313 29547 25379 29550
rect 35617 29610 35683 29613
rect 36905 29610 36971 29613
rect 35617 29608 36971 29610
rect 35617 29552 35622 29608
rect 35678 29552 36910 29608
rect 36966 29552 36971 29608
rect 35617 29550 36971 29552
rect 35617 29547 35683 29550
rect 36905 29547 36971 29550
rect 11513 29474 11579 29477
rect 13537 29474 13603 29477
rect 11513 29472 13603 29474
rect 11513 29416 11518 29472
rect 11574 29416 13542 29472
rect 13598 29416 13603 29472
rect 11513 29414 13603 29416
rect 11513 29411 11579 29414
rect 13537 29411 13603 29414
rect 23013 29474 23079 29477
rect 24025 29474 24091 29477
rect 23013 29472 24091 29474
rect 23013 29416 23018 29472
rect 23074 29416 24030 29472
rect 24086 29416 24091 29472
rect 23013 29414 24091 29416
rect 23013 29411 23079 29414
rect 24025 29411 24091 29414
rect 24301 29474 24367 29477
rect 24669 29474 24735 29477
rect 24301 29472 24735 29474
rect 24301 29416 24306 29472
rect 24362 29416 24674 29472
rect 24730 29416 24735 29472
rect 24301 29414 24735 29416
rect 24301 29411 24367 29414
rect 24669 29411 24735 29414
rect 33961 29474 34027 29477
rect 34145 29474 34211 29477
rect 35065 29474 35131 29477
rect 33961 29472 35131 29474
rect 33961 29416 33966 29472
rect 34022 29416 34150 29472
rect 34206 29416 35070 29472
rect 35126 29416 35131 29472
rect 33961 29414 35131 29416
rect 33961 29411 34027 29414
rect 34145 29411 34211 29414
rect 35065 29411 35131 29414
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 23657 29338 23723 29341
rect 26417 29338 26483 29341
rect 23657 29336 26483 29338
rect 23657 29280 23662 29336
rect 23718 29280 26422 29336
rect 26478 29280 26483 29336
rect 23657 29278 26483 29280
rect 23657 29275 23723 29278
rect 26417 29275 26483 29278
rect 33501 29338 33567 29341
rect 34973 29338 35039 29341
rect 35382 29338 35388 29340
rect 33501 29336 34898 29338
rect 33501 29280 33506 29336
rect 33562 29280 34898 29336
rect 33501 29278 34898 29280
rect 33501 29275 33567 29278
rect 17769 29202 17835 29205
rect 33685 29202 33751 29205
rect 17769 29200 33751 29202
rect 17769 29144 17774 29200
rect 17830 29144 33690 29200
rect 33746 29144 33751 29200
rect 17769 29142 33751 29144
rect 17769 29139 17835 29142
rect 33685 29139 33751 29142
rect 33869 29202 33935 29205
rect 34605 29202 34671 29205
rect 33869 29200 34671 29202
rect 33869 29144 33874 29200
rect 33930 29144 34610 29200
rect 34666 29144 34671 29200
rect 33869 29142 34671 29144
rect 34838 29202 34898 29278
rect 34973 29336 35388 29338
rect 34973 29280 34978 29336
rect 35034 29280 35388 29336
rect 34973 29278 35388 29280
rect 34973 29275 35039 29278
rect 35382 29276 35388 29278
rect 35452 29276 35458 29340
rect 35709 29202 35775 29205
rect 36077 29204 36143 29205
rect 36077 29202 36124 29204
rect 34838 29200 35775 29202
rect 34838 29144 35714 29200
rect 35770 29144 35775 29200
rect 34838 29142 35775 29144
rect 36032 29200 36124 29202
rect 36032 29144 36082 29200
rect 36032 29142 36124 29144
rect 33869 29139 33935 29142
rect 34605 29139 34671 29142
rect 35709 29139 35775 29142
rect 36077 29140 36124 29142
rect 36188 29140 36194 29204
rect 36077 29139 36143 29140
rect 20110 29004 20116 29068
rect 20180 29066 20186 29068
rect 20713 29066 20779 29069
rect 20180 29064 20779 29066
rect 20180 29008 20718 29064
rect 20774 29008 20779 29064
rect 20180 29006 20779 29008
rect 20180 29004 20186 29006
rect 20713 29003 20779 29006
rect 21541 29066 21607 29069
rect 24485 29066 24551 29069
rect 30281 29066 30347 29069
rect 21541 29064 30347 29066
rect 21541 29008 21546 29064
rect 21602 29008 24490 29064
rect 24546 29008 30286 29064
rect 30342 29008 30347 29064
rect 21541 29006 30347 29008
rect 21541 29003 21607 29006
rect 24485 29003 24551 29006
rect 30281 29003 30347 29006
rect 33501 29066 33567 29069
rect 37733 29066 37799 29069
rect 33501 29064 37799 29066
rect 33501 29008 33506 29064
rect 33562 29008 37738 29064
rect 37794 29008 37799 29064
rect 33501 29006 37799 29008
rect 33501 29003 33567 29006
rect 37733 29003 37799 29006
rect 23197 28930 23263 28933
rect 23841 28930 23907 28933
rect 34697 28932 34763 28933
rect 23197 28928 23907 28930
rect 23197 28872 23202 28928
rect 23258 28872 23846 28928
rect 23902 28872 23907 28928
rect 23197 28870 23907 28872
rect 23197 28867 23263 28870
rect 23841 28867 23907 28870
rect 34646 28868 34652 28932
rect 34716 28930 34763 28932
rect 34716 28928 34808 28930
rect 34758 28872 34808 28928
rect 34716 28870 34808 28872
rect 34716 28868 34763 28870
rect 34697 28867 34763 28868
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 21173 28522 21239 28525
rect 24209 28522 24275 28525
rect 21173 28520 24275 28522
rect 21173 28464 21178 28520
rect 21234 28464 24214 28520
rect 24270 28464 24275 28520
rect 21173 28462 24275 28464
rect 21173 28459 21239 28462
rect 24209 28459 24275 28462
rect 25589 28522 25655 28525
rect 26141 28522 26207 28525
rect 25589 28520 26207 28522
rect 25589 28464 25594 28520
rect 25650 28464 26146 28520
rect 26202 28464 26207 28520
rect 25589 28462 26207 28464
rect 25589 28459 25655 28462
rect 26141 28459 26207 28462
rect 26509 28522 26575 28525
rect 27102 28522 27108 28524
rect 26509 28520 27108 28522
rect 26509 28464 26514 28520
rect 26570 28464 27108 28520
rect 26509 28462 27108 28464
rect 26509 28459 26575 28462
rect 27102 28460 27108 28462
rect 27172 28460 27178 28524
rect 21449 28386 21515 28389
rect 26509 28386 26575 28389
rect 21449 28384 26575 28386
rect 21449 28328 21454 28384
rect 21510 28328 26514 28384
rect 26570 28328 26575 28384
rect 21449 28326 26575 28328
rect 21449 28323 21515 28326
rect 26509 28323 26575 28326
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 21173 28250 21239 28253
rect 30598 28250 30604 28252
rect 21173 28248 30604 28250
rect 21173 28192 21178 28248
rect 21234 28192 30604 28248
rect 21173 28190 30604 28192
rect 21173 28187 21239 28190
rect 30598 28188 30604 28190
rect 30668 28188 30674 28252
rect 5993 28116 6059 28117
rect 5942 28114 5948 28116
rect 5866 28054 5948 28114
rect 6012 28114 6059 28116
rect 7097 28114 7163 28117
rect 6012 28112 7163 28114
rect 6054 28056 7102 28112
rect 7158 28056 7163 28112
rect 5942 28052 5948 28054
rect 6012 28054 7163 28056
rect 6012 28052 6059 28054
rect 5993 28051 6059 28052
rect 7097 28051 7163 28054
rect 9857 27978 9923 27981
rect 9990 27978 9996 27980
rect 9857 27976 9996 27978
rect 9857 27920 9862 27976
rect 9918 27920 9996 27976
rect 9857 27918 9996 27920
rect 9857 27915 9923 27918
rect 9990 27916 9996 27918
rect 10060 27916 10066 27980
rect 12525 27842 12591 27845
rect 14365 27842 14431 27845
rect 12525 27840 14431 27842
rect 12525 27784 12530 27840
rect 12586 27784 14370 27840
rect 14426 27784 14431 27840
rect 12525 27782 14431 27784
rect 12525 27779 12591 27782
rect 14365 27779 14431 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19926 27644 19932 27708
rect 19996 27706 20002 27708
rect 21817 27706 21883 27709
rect 19996 27704 21883 27706
rect 19996 27648 21822 27704
rect 21878 27648 21883 27704
rect 19996 27646 21883 27648
rect 19996 27644 20002 27646
rect 21817 27643 21883 27646
rect 18505 27570 18571 27573
rect 18965 27570 19031 27573
rect 18505 27568 19031 27570
rect 18505 27512 18510 27568
rect 18566 27512 18970 27568
rect 19026 27512 19031 27568
rect 18505 27510 19031 27512
rect 18505 27507 18571 27510
rect 18965 27507 19031 27510
rect 32765 27570 32831 27573
rect 32765 27568 37290 27570
rect 32765 27512 32770 27568
rect 32826 27512 37290 27568
rect 32765 27510 37290 27512
rect 32765 27507 32831 27510
rect 13721 27434 13787 27437
rect 15561 27434 15627 27437
rect 31109 27434 31175 27437
rect 13721 27432 31175 27434
rect 13721 27376 13726 27432
rect 13782 27376 15566 27432
rect 15622 27376 31114 27432
rect 31170 27376 31175 27432
rect 13721 27374 31175 27376
rect 37230 27434 37290 27510
rect 37365 27434 37431 27437
rect 37230 27432 37431 27434
rect 37230 27376 37370 27432
rect 37426 27376 37431 27432
rect 37230 27374 37431 27376
rect 13721 27371 13787 27374
rect 15561 27371 15627 27374
rect 31109 27371 31175 27374
rect 37365 27371 37431 27374
rect 10685 27298 10751 27301
rect 14825 27298 14891 27301
rect 32765 27300 32831 27301
rect 32765 27298 32812 27300
rect 10685 27296 14891 27298
rect 10685 27240 10690 27296
rect 10746 27240 14830 27296
rect 14886 27240 14891 27296
rect 10685 27238 14891 27240
rect 32720 27296 32812 27298
rect 32720 27240 32770 27296
rect 32720 27238 32812 27240
rect 10685 27235 10751 27238
rect 14825 27235 14891 27238
rect 32765 27236 32812 27238
rect 32876 27236 32882 27300
rect 39573 27298 39639 27301
rect 40957 27298 41757 27328
rect 39573 27296 41757 27298
rect 39573 27240 39578 27296
rect 39634 27240 41757 27296
rect 39573 27238 41757 27240
rect 32765 27235 32831 27236
rect 39573 27235 39639 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 40957 27208 41757 27238
rect 35590 27167 35906 27168
rect 10685 27162 10751 27165
rect 16481 27162 16547 27165
rect 37089 27162 37155 27165
rect 10685 27160 16547 27162
rect 10685 27104 10690 27160
rect 10746 27104 16486 27160
rect 16542 27104 16547 27160
rect 10685 27102 16547 27104
rect 10685 27099 10751 27102
rect 16481 27099 16547 27102
rect 37046 27160 37155 27162
rect 37046 27104 37094 27160
rect 37150 27104 37155 27160
rect 37046 27099 37155 27104
rect 8385 27026 8451 27029
rect 17217 27026 17283 27029
rect 30465 27026 30531 27029
rect 30741 27026 30807 27029
rect 32305 27026 32371 27029
rect 37046 27026 37106 27099
rect 38101 27026 38167 27029
rect 8385 27024 38167 27026
rect 8385 26968 8390 27024
rect 8446 26968 17222 27024
rect 17278 26968 30470 27024
rect 30526 26968 30746 27024
rect 30802 26968 32310 27024
rect 32366 26968 38106 27024
rect 38162 26968 38167 27024
rect 8385 26966 38167 26968
rect 8385 26963 8451 26966
rect 17217 26963 17283 26966
rect 30465 26963 30531 26966
rect 30741 26963 30807 26966
rect 32305 26963 32371 26966
rect 38101 26963 38167 26966
rect 19425 26890 19491 26893
rect 21357 26890 21423 26893
rect 19425 26888 21423 26890
rect 19425 26832 19430 26888
rect 19486 26832 21362 26888
rect 21418 26832 21423 26888
rect 19425 26830 21423 26832
rect 19425 26827 19491 26830
rect 21357 26827 21423 26830
rect 22185 26890 22251 26893
rect 22318 26890 22324 26892
rect 22185 26888 22324 26890
rect 22185 26832 22190 26888
rect 22246 26832 22324 26888
rect 22185 26830 22324 26832
rect 22185 26827 22251 26830
rect 22318 26828 22324 26830
rect 22388 26828 22394 26892
rect 31017 26890 31083 26893
rect 32489 26890 32555 26893
rect 35617 26890 35683 26893
rect 31017 26888 35683 26890
rect 31017 26832 31022 26888
rect 31078 26832 32494 26888
rect 32550 26832 35622 26888
rect 35678 26832 35683 26888
rect 31017 26830 35683 26832
rect 31017 26827 31083 26830
rect 32489 26827 32555 26830
rect 35617 26827 35683 26830
rect 6729 26754 6795 26757
rect 20713 26754 20779 26757
rect 22645 26754 22711 26757
rect 6729 26752 12450 26754
rect 6729 26696 6734 26752
rect 6790 26696 12450 26752
rect 6729 26694 12450 26696
rect 6729 26691 6795 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 8937 26620 9003 26621
rect 8334 26556 8340 26620
rect 8404 26618 8410 26620
rect 8886 26618 8892 26620
rect 8404 26558 8892 26618
rect 8956 26616 9003 26620
rect 8998 26560 9003 26616
rect 8404 26556 8410 26558
rect 8886 26556 8892 26558
rect 8956 26556 9003 26560
rect 12390 26618 12450 26694
rect 20713 26752 22711 26754
rect 20713 26696 20718 26752
rect 20774 26696 22650 26752
rect 22706 26696 22711 26752
rect 20713 26694 22711 26696
rect 20713 26691 20779 26694
rect 22645 26691 22711 26694
rect 29729 26754 29795 26757
rect 33225 26754 33291 26757
rect 29729 26752 33291 26754
rect 29729 26696 29734 26752
rect 29790 26696 33230 26752
rect 33286 26696 33291 26752
rect 29729 26694 33291 26696
rect 29729 26691 29795 26694
rect 33225 26691 33291 26694
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 14641 26618 14707 26621
rect 22185 26620 22251 26621
rect 12390 26616 14707 26618
rect 12390 26560 14646 26616
rect 14702 26560 14707 26616
rect 12390 26558 14707 26560
rect 8937 26555 9003 26556
rect 14641 26555 14707 26558
rect 22134 26556 22140 26620
rect 22204 26618 22251 26620
rect 22461 26620 22527 26621
rect 22461 26618 22508 26620
rect 22204 26616 22296 26618
rect 22246 26560 22296 26616
rect 22204 26558 22296 26560
rect 22416 26616 22508 26618
rect 22416 26560 22466 26616
rect 22416 26558 22508 26560
rect 22204 26556 22251 26558
rect 22185 26555 22251 26556
rect 22461 26556 22508 26558
rect 22572 26556 22578 26620
rect 32305 26618 32371 26621
rect 32489 26618 32555 26621
rect 32305 26616 32555 26618
rect 32305 26560 32310 26616
rect 32366 26560 32494 26616
rect 32550 26560 32555 26616
rect 32305 26558 32555 26560
rect 22461 26555 22527 26556
rect 32305 26555 32371 26558
rect 32489 26555 32555 26558
rect 40217 26618 40283 26621
rect 40957 26618 41757 26648
rect 40217 26616 41757 26618
rect 40217 26560 40222 26616
rect 40278 26560 41757 26616
rect 40217 26558 41757 26560
rect 40217 26555 40283 26558
rect 40957 26528 41757 26558
rect 10961 26482 11027 26485
rect 14089 26482 14155 26485
rect 10961 26480 14155 26482
rect 10961 26424 10966 26480
rect 11022 26424 14094 26480
rect 14150 26424 14155 26480
rect 10961 26422 14155 26424
rect 10961 26419 11027 26422
rect 14089 26419 14155 26422
rect 14549 26482 14615 26485
rect 15653 26482 15719 26485
rect 16849 26482 16915 26485
rect 33593 26482 33659 26485
rect 14549 26480 33659 26482
rect 14549 26424 14554 26480
rect 14610 26424 15658 26480
rect 15714 26424 16854 26480
rect 16910 26424 33598 26480
rect 33654 26424 33659 26480
rect 14549 26422 33659 26424
rect 14549 26419 14615 26422
rect 15653 26419 15719 26422
rect 16849 26419 16915 26422
rect 33593 26419 33659 26422
rect 15653 26346 15719 26349
rect 16941 26348 17007 26349
rect 21817 26348 21883 26349
rect 16430 26346 16436 26348
rect 15653 26344 16436 26346
rect 15653 26288 15658 26344
rect 15714 26288 16436 26344
rect 15653 26286 16436 26288
rect 15653 26283 15719 26286
rect 16430 26284 16436 26286
rect 16500 26284 16506 26348
rect 16941 26344 16988 26348
rect 17052 26346 17058 26348
rect 16941 26288 16946 26344
rect 16941 26284 16988 26288
rect 17052 26286 17098 26346
rect 17052 26284 17058 26286
rect 19190 26284 19196 26348
rect 19260 26346 19266 26348
rect 21766 26346 21772 26348
rect 19260 26286 21650 26346
rect 21726 26286 21772 26346
rect 21836 26344 21883 26348
rect 22185 26346 22251 26349
rect 21878 26288 21883 26344
rect 19260 26284 19266 26286
rect 16941 26283 17007 26284
rect 12617 26210 12683 26213
rect 17309 26210 17375 26213
rect 12617 26208 17375 26210
rect 12617 26152 12622 26208
rect 12678 26152 17314 26208
rect 17370 26152 17375 26208
rect 12617 26150 17375 26152
rect 21590 26210 21650 26286
rect 21766 26284 21772 26286
rect 21836 26284 21883 26288
rect 21817 26283 21883 26284
rect 21958 26344 22251 26346
rect 21958 26288 22190 26344
rect 22246 26288 22251 26344
rect 21958 26286 22251 26288
rect 21958 26210 22018 26286
rect 22185 26283 22251 26286
rect 22369 26346 22435 26349
rect 23013 26346 23079 26349
rect 22369 26344 23079 26346
rect 22369 26288 22374 26344
rect 22430 26288 23018 26344
rect 23074 26288 23079 26344
rect 22369 26286 23079 26288
rect 22369 26283 22435 26286
rect 23013 26283 23079 26286
rect 27797 26346 27863 26349
rect 28022 26346 28028 26348
rect 27797 26344 28028 26346
rect 27797 26288 27802 26344
rect 27858 26288 28028 26344
rect 27797 26286 28028 26288
rect 27797 26283 27863 26286
rect 28022 26284 28028 26286
rect 28092 26284 28098 26348
rect 28390 26284 28396 26348
rect 28460 26346 28466 26348
rect 28809 26346 28875 26349
rect 28460 26344 28875 26346
rect 28460 26288 28814 26344
rect 28870 26288 28875 26344
rect 28460 26286 28875 26288
rect 28460 26284 28466 26286
rect 28809 26283 28875 26286
rect 30782 26284 30788 26348
rect 30852 26346 30858 26348
rect 30925 26346 30991 26349
rect 30852 26344 30991 26346
rect 30852 26288 30930 26344
rect 30986 26288 30991 26344
rect 30852 26286 30991 26288
rect 30852 26284 30858 26286
rect 30925 26283 30991 26286
rect 31661 26346 31727 26349
rect 31845 26346 31911 26349
rect 31661 26344 31911 26346
rect 31661 26288 31666 26344
rect 31722 26288 31850 26344
rect 31906 26288 31911 26344
rect 31661 26286 31911 26288
rect 31661 26283 31727 26286
rect 31845 26283 31911 26286
rect 32489 26346 32555 26349
rect 38377 26346 38443 26349
rect 38510 26346 38516 26348
rect 32489 26344 38516 26346
rect 32489 26288 32494 26344
rect 32550 26288 38382 26344
rect 38438 26288 38516 26344
rect 32489 26286 38516 26288
rect 32489 26283 32555 26286
rect 38377 26283 38443 26286
rect 38510 26284 38516 26286
rect 38580 26284 38586 26348
rect 21590 26150 22018 26210
rect 27889 26210 27955 26213
rect 28625 26210 28691 26213
rect 27889 26208 28691 26210
rect 27889 26152 27894 26208
rect 27950 26152 28630 26208
rect 28686 26152 28691 26208
rect 27889 26150 28691 26152
rect 12617 26147 12683 26150
rect 17309 26147 17375 26150
rect 27889 26147 27955 26150
rect 28625 26147 28691 26150
rect 34697 26210 34763 26213
rect 35157 26210 35223 26213
rect 34697 26208 35223 26210
rect 34697 26152 34702 26208
rect 34758 26152 35162 26208
rect 35218 26152 35223 26208
rect 34697 26150 35223 26152
rect 34697 26147 34763 26150
rect 35157 26147 35223 26150
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 13629 25940 13695 25941
rect 13629 25938 13676 25940
rect 13584 25936 13676 25938
rect 13584 25880 13634 25936
rect 13584 25878 13676 25880
rect 13629 25876 13676 25878
rect 13740 25876 13746 25940
rect 14181 25938 14247 25941
rect 39941 25938 40007 25941
rect 40957 25938 41757 25968
rect 14181 25936 14290 25938
rect 14181 25880 14186 25936
rect 14242 25880 14290 25936
rect 13629 25875 13695 25876
rect 14181 25875 14290 25880
rect 39941 25936 41757 25938
rect 39941 25880 39946 25936
rect 40002 25880 41757 25936
rect 39941 25878 41757 25880
rect 39941 25875 40007 25878
rect 14230 25669 14290 25875
rect 40957 25848 41757 25878
rect 29361 25804 29427 25805
rect 29310 25740 29316 25804
rect 29380 25802 29427 25804
rect 29380 25800 29472 25802
rect 29422 25744 29472 25800
rect 29380 25742 29472 25744
rect 29380 25740 29427 25742
rect 29361 25739 29427 25740
rect 14181 25664 14290 25669
rect 14181 25608 14186 25664
rect 14242 25608 14290 25664
rect 14181 25606 14290 25608
rect 23289 25666 23355 25669
rect 32254 25666 32260 25668
rect 23289 25664 32260 25666
rect 23289 25608 23294 25664
rect 23350 25608 32260 25664
rect 23289 25606 32260 25608
rect 14181 25603 14247 25606
rect 23289 25603 23355 25606
rect 32254 25604 32260 25606
rect 32324 25604 32330 25668
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 17350 25468 17356 25532
rect 17420 25530 17426 25532
rect 18321 25530 18387 25533
rect 24853 25532 24919 25533
rect 24853 25530 24900 25532
rect 17420 25528 18387 25530
rect 17420 25472 18326 25528
rect 18382 25472 18387 25528
rect 17420 25470 18387 25472
rect 24808 25528 24900 25530
rect 24808 25472 24858 25528
rect 24808 25470 24900 25472
rect 17420 25468 17426 25470
rect 18321 25467 18387 25470
rect 24853 25468 24900 25470
rect 24964 25468 24970 25532
rect 24853 25467 24919 25468
rect 4654 25332 4660 25396
rect 4724 25394 4730 25396
rect 4797 25394 4863 25397
rect 4724 25392 4863 25394
rect 4724 25336 4802 25392
rect 4858 25336 4863 25392
rect 4724 25334 4863 25336
rect 4724 25332 4730 25334
rect 4797 25331 4863 25334
rect 16246 25332 16252 25396
rect 16316 25394 16322 25396
rect 26693 25394 26759 25397
rect 26969 25394 27035 25397
rect 16316 25392 27035 25394
rect 16316 25336 26698 25392
rect 26754 25336 26974 25392
rect 27030 25336 27035 25392
rect 16316 25334 27035 25336
rect 16316 25332 16322 25334
rect 26693 25331 26759 25334
rect 26969 25331 27035 25334
rect 31937 25394 32003 25397
rect 36813 25394 36879 25397
rect 31937 25392 36879 25394
rect 31937 25336 31942 25392
rect 31998 25336 36818 25392
rect 36874 25336 36879 25392
rect 31937 25334 36879 25336
rect 31937 25331 32003 25334
rect 36813 25331 36879 25334
rect 7097 25258 7163 25261
rect 8201 25258 8267 25261
rect 7097 25256 8267 25258
rect 7097 25200 7102 25256
rect 7158 25200 8206 25256
rect 8262 25200 8267 25256
rect 7097 25198 8267 25200
rect 7097 25195 7163 25198
rect 8201 25195 8267 25198
rect 17125 25258 17191 25261
rect 33685 25260 33751 25261
rect 21214 25258 21220 25260
rect 17125 25256 21220 25258
rect 17125 25200 17130 25256
rect 17186 25200 21220 25256
rect 17125 25198 21220 25200
rect 17125 25195 17191 25198
rect 21214 25196 21220 25198
rect 21284 25196 21290 25260
rect 33685 25258 33732 25260
rect 33640 25256 33732 25258
rect 33640 25200 33690 25256
rect 33640 25198 33732 25200
rect 33685 25196 33732 25198
rect 33796 25196 33802 25260
rect 35382 25196 35388 25260
rect 35452 25258 35458 25260
rect 35525 25258 35591 25261
rect 35452 25256 35591 25258
rect 35452 25200 35530 25256
rect 35586 25200 35591 25256
rect 35452 25198 35591 25200
rect 35452 25196 35458 25198
rect 33685 25195 33751 25196
rect 35525 25195 35591 25198
rect 6085 25124 6151 25125
rect 8385 25124 8451 25125
rect 6085 25120 6132 25124
rect 6196 25122 6202 25124
rect 6085 25064 6090 25120
rect 6085 25060 6132 25064
rect 6196 25062 6242 25122
rect 6196 25060 6202 25062
rect 8334 25060 8340 25124
rect 8404 25122 8451 25124
rect 8404 25120 8496 25122
rect 8446 25064 8496 25120
rect 8404 25062 8496 25064
rect 8404 25060 8451 25062
rect 21398 25060 21404 25124
rect 21468 25122 21474 25124
rect 27613 25122 27679 25125
rect 21468 25120 27679 25122
rect 21468 25064 27618 25120
rect 27674 25064 27679 25120
rect 21468 25062 27679 25064
rect 21468 25060 21474 25062
rect 6085 25059 6151 25060
rect 8385 25059 8451 25060
rect 27613 25059 27679 25062
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 13905 24986 13971 24989
rect 14222 24986 14228 24988
rect 13905 24984 14228 24986
rect 13905 24928 13910 24984
rect 13966 24928 14228 24984
rect 13905 24926 14228 24928
rect 13905 24923 13971 24926
rect 14222 24924 14228 24926
rect 14292 24924 14298 24988
rect 20161 24986 20227 24989
rect 24526 24986 24532 24988
rect 20161 24984 24532 24986
rect 20161 24928 20166 24984
rect 20222 24928 24532 24984
rect 20161 24926 24532 24928
rect 20161 24923 20227 24926
rect 24526 24924 24532 24926
rect 24596 24924 24602 24988
rect 32489 24986 32555 24989
rect 32990 24986 32996 24988
rect 32489 24984 32996 24986
rect 32489 24928 32494 24984
rect 32550 24928 32996 24984
rect 32489 24926 32996 24928
rect 32489 24923 32555 24926
rect 32990 24924 32996 24926
rect 33060 24924 33066 24988
rect 10409 24850 10475 24853
rect 11973 24850 12039 24853
rect 10409 24848 12039 24850
rect 10409 24792 10414 24848
rect 10470 24792 11978 24848
rect 12034 24792 12039 24848
rect 10409 24790 12039 24792
rect 10409 24787 10475 24790
rect 11973 24787 12039 24790
rect 21081 24850 21147 24853
rect 22134 24850 22140 24852
rect 21081 24848 22140 24850
rect 21081 24792 21086 24848
rect 21142 24792 22140 24848
rect 21081 24790 22140 24792
rect 21081 24787 21147 24790
rect 22134 24788 22140 24790
rect 22204 24850 22210 24852
rect 23657 24850 23723 24853
rect 24761 24850 24827 24853
rect 22204 24848 24827 24850
rect 22204 24792 23662 24848
rect 23718 24792 24766 24848
rect 24822 24792 24827 24848
rect 22204 24790 24827 24792
rect 22204 24788 22210 24790
rect 23657 24787 23723 24790
rect 24761 24787 24827 24790
rect 25405 24850 25471 24853
rect 26233 24850 26299 24853
rect 32397 24852 32463 24853
rect 32397 24850 32444 24852
rect 25405 24848 26299 24850
rect 25405 24792 25410 24848
rect 25466 24792 26238 24848
rect 26294 24792 26299 24848
rect 25405 24790 26299 24792
rect 32352 24848 32444 24850
rect 32508 24850 32514 24852
rect 38193 24850 38259 24853
rect 32508 24848 38259 24850
rect 32352 24792 32402 24848
rect 32508 24792 38198 24848
rect 38254 24792 38259 24848
rect 32352 24790 32444 24792
rect 25405 24787 25471 24790
rect 26233 24787 26299 24790
rect 32397 24788 32444 24790
rect 32508 24790 38259 24792
rect 32508 24788 32514 24790
rect 32397 24787 32463 24788
rect 38193 24787 38259 24790
rect 34646 24652 34652 24716
rect 34716 24714 34722 24716
rect 35249 24714 35315 24717
rect 34716 24712 35315 24714
rect 34716 24656 35254 24712
rect 35310 24656 35315 24712
rect 34716 24654 35315 24656
rect 34716 24652 34722 24654
rect 35249 24651 35315 24654
rect 6545 24578 6611 24581
rect 9029 24578 9095 24581
rect 11789 24578 11855 24581
rect 14733 24578 14799 24581
rect 6545 24576 14799 24578
rect 6545 24520 6550 24576
rect 6606 24520 9034 24576
rect 9090 24520 11794 24576
rect 11850 24520 14738 24576
rect 14794 24520 14799 24576
rect 6545 24518 14799 24520
rect 6545 24515 6611 24518
rect 9029 24515 9095 24518
rect 11789 24515 11855 24518
rect 14733 24515 14799 24518
rect 40217 24578 40283 24581
rect 40957 24578 41757 24608
rect 40217 24576 41757 24578
rect 40217 24520 40222 24576
rect 40278 24520 41757 24576
rect 40217 24518 41757 24520
rect 40217 24515 40283 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 40957 24488 41757 24518
rect 34930 24447 35246 24448
rect 6361 24442 6427 24445
rect 7925 24442 7991 24445
rect 9305 24442 9371 24445
rect 6361 24440 9371 24442
rect 6361 24384 6366 24440
rect 6422 24384 7930 24440
rect 7986 24384 9310 24440
rect 9366 24384 9371 24440
rect 6361 24382 9371 24384
rect 6361 24379 6427 24382
rect 7925 24379 7991 24382
rect 9305 24379 9371 24382
rect 8109 24306 8175 24309
rect 9213 24306 9279 24309
rect 8109 24304 9279 24306
rect 8109 24248 8114 24304
rect 8170 24248 9218 24304
rect 9274 24248 9279 24304
rect 8109 24246 9279 24248
rect 8109 24243 8175 24246
rect 9213 24243 9279 24246
rect 9673 24306 9739 24309
rect 9990 24306 9996 24308
rect 9673 24304 9996 24306
rect 9673 24248 9678 24304
rect 9734 24248 9996 24304
rect 9673 24246 9996 24248
rect 9673 24243 9739 24246
rect 9990 24244 9996 24246
rect 10060 24244 10066 24308
rect 26417 24306 26483 24309
rect 28165 24306 28231 24309
rect 26417 24304 28231 24306
rect 26417 24248 26422 24304
rect 26478 24248 28170 24304
rect 28226 24248 28231 24304
rect 26417 24246 28231 24248
rect 26417 24243 26483 24246
rect 28165 24243 28231 24246
rect 28533 24306 28599 24309
rect 28758 24306 28764 24308
rect 28533 24304 28764 24306
rect 28533 24248 28538 24304
rect 28594 24248 28764 24304
rect 28533 24246 28764 24248
rect 28533 24243 28599 24246
rect 28758 24244 28764 24246
rect 28828 24244 28834 24308
rect 24894 24108 24900 24172
rect 24964 24170 24970 24172
rect 25129 24170 25195 24173
rect 24964 24168 25195 24170
rect 24964 24112 25134 24168
rect 25190 24112 25195 24168
rect 24964 24110 25195 24112
rect 24964 24108 24970 24110
rect 25129 24107 25195 24110
rect 25865 24170 25931 24173
rect 25998 24170 26004 24172
rect 25865 24168 26004 24170
rect 25865 24112 25870 24168
rect 25926 24112 26004 24168
rect 25865 24110 26004 24112
rect 25865 24107 25931 24110
rect 25998 24108 26004 24110
rect 26068 24108 26074 24172
rect 8661 24034 8727 24037
rect 8937 24034 9003 24037
rect 8661 24032 9003 24034
rect 8661 23976 8666 24032
rect 8722 23976 8942 24032
rect 8998 23976 9003 24032
rect 8661 23974 9003 23976
rect 8661 23971 8727 23974
rect 8937 23971 9003 23974
rect 19885 24034 19951 24037
rect 20437 24034 20503 24037
rect 19885 24032 20503 24034
rect 19885 23976 19890 24032
rect 19946 23976 20442 24032
rect 20498 23976 20503 24032
rect 19885 23974 20503 23976
rect 19885 23971 19951 23974
rect 20437 23971 20503 23974
rect 22093 24034 22159 24037
rect 24025 24034 24091 24037
rect 22093 24032 24091 24034
rect 22093 23976 22098 24032
rect 22154 23976 24030 24032
rect 24086 23976 24091 24032
rect 22093 23974 24091 23976
rect 22093 23971 22159 23974
rect 24025 23971 24091 23974
rect 24209 24034 24275 24037
rect 28257 24034 28323 24037
rect 24209 24032 28323 24034
rect 24209 23976 24214 24032
rect 24270 23976 28262 24032
rect 28318 23976 28323 24032
rect 24209 23974 28323 23976
rect 24209 23971 24275 23974
rect 28257 23971 28323 23974
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 35590 23903 35906 23904
rect 6085 23898 6151 23901
rect 6545 23898 6611 23901
rect 8661 23898 8727 23901
rect 6085 23896 8727 23898
rect 6085 23840 6090 23896
rect 6146 23840 6550 23896
rect 6606 23840 8666 23896
rect 8722 23840 8727 23896
rect 6085 23838 8727 23840
rect 6085 23835 6151 23838
rect 6545 23835 6611 23838
rect 8661 23835 8727 23838
rect 19517 23898 19583 23901
rect 22553 23898 22619 23901
rect 23013 23898 23079 23901
rect 23473 23898 23539 23901
rect 19517 23896 23539 23898
rect 19517 23840 19522 23896
rect 19578 23840 22558 23896
rect 22614 23840 23018 23896
rect 23074 23840 23478 23896
rect 23534 23840 23539 23896
rect 19517 23838 23539 23840
rect 19517 23835 19583 23838
rect 22553 23835 22619 23838
rect 23013 23835 23079 23838
rect 23473 23835 23539 23838
rect 27981 23898 28047 23901
rect 39665 23898 39731 23901
rect 40957 23898 41757 23928
rect 27981 23896 31770 23898
rect 27981 23840 27986 23896
rect 28042 23840 31770 23896
rect 27981 23838 31770 23840
rect 27981 23835 28047 23838
rect 5073 23762 5139 23765
rect 7465 23762 7531 23765
rect 5073 23760 7531 23762
rect 5073 23704 5078 23760
rect 5134 23704 7470 23760
rect 7526 23704 7531 23760
rect 5073 23702 7531 23704
rect 5073 23699 5139 23702
rect 7465 23699 7531 23702
rect 8569 23762 8635 23765
rect 9121 23762 9187 23765
rect 8569 23760 9187 23762
rect 8569 23704 8574 23760
rect 8630 23704 9126 23760
rect 9182 23704 9187 23760
rect 8569 23702 9187 23704
rect 8569 23699 8635 23702
rect 9121 23699 9187 23702
rect 19333 23762 19399 23765
rect 22737 23762 22803 23765
rect 25313 23762 25379 23765
rect 28441 23762 28507 23765
rect 19333 23760 28507 23762
rect 19333 23704 19338 23760
rect 19394 23704 22742 23760
rect 22798 23704 25318 23760
rect 25374 23704 28446 23760
rect 28502 23704 28507 23760
rect 19333 23702 28507 23704
rect 19333 23699 19399 23702
rect 22737 23699 22803 23702
rect 25313 23699 25379 23702
rect 28441 23699 28507 23702
rect 5758 23564 5764 23628
rect 5828 23626 5834 23628
rect 6177 23626 6243 23629
rect 5828 23624 6243 23626
rect 5828 23568 6182 23624
rect 6238 23568 6243 23624
rect 5828 23566 6243 23568
rect 5828 23564 5834 23566
rect 6177 23563 6243 23566
rect 18413 23626 18479 23629
rect 19149 23626 19215 23629
rect 18413 23624 19215 23626
rect 18413 23568 18418 23624
rect 18474 23568 19154 23624
rect 19210 23568 19215 23624
rect 18413 23566 19215 23568
rect 18413 23563 18479 23566
rect 19149 23563 19215 23566
rect 5441 23490 5507 23493
rect 5942 23490 5948 23492
rect 5441 23488 5948 23490
rect 5441 23432 5446 23488
rect 5502 23432 5948 23488
rect 5441 23430 5948 23432
rect 5441 23427 5507 23430
rect 5942 23428 5948 23430
rect 6012 23428 6018 23492
rect 23381 23490 23447 23493
rect 23974 23490 23980 23492
rect 23381 23488 23980 23490
rect 23381 23432 23386 23488
rect 23442 23432 23980 23488
rect 23381 23430 23980 23432
rect 23381 23427 23447 23430
rect 23974 23428 23980 23430
rect 24044 23428 24050 23492
rect 31710 23490 31770 23838
rect 39665 23896 41757 23898
rect 39665 23840 39670 23896
rect 39726 23840 41757 23896
rect 39665 23838 41757 23840
rect 39665 23835 39731 23838
rect 40957 23808 41757 23838
rect 33133 23762 33199 23765
rect 34881 23762 34947 23765
rect 33133 23760 34947 23762
rect 33133 23704 33138 23760
rect 33194 23704 34886 23760
rect 34942 23704 34947 23760
rect 33133 23702 34947 23704
rect 33133 23699 33199 23702
rect 34881 23699 34947 23702
rect 32305 23626 32371 23629
rect 34789 23626 34855 23629
rect 32305 23624 34855 23626
rect 32305 23568 32310 23624
rect 32366 23568 34794 23624
rect 34850 23568 34855 23624
rect 32305 23566 34855 23568
rect 32305 23563 32371 23566
rect 34789 23563 34855 23566
rect 34462 23490 34468 23492
rect 31710 23430 34468 23490
rect 34462 23428 34468 23430
rect 34532 23428 34538 23492
rect 37273 23490 37339 23493
rect 37406 23490 37412 23492
rect 37273 23488 37412 23490
rect 37273 23432 37278 23488
rect 37334 23432 37412 23488
rect 37273 23430 37412 23432
rect 37273 23427 37339 23430
rect 37406 23428 37412 23430
rect 37476 23428 37482 23492
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 10225 23354 10291 23357
rect 10182 23352 10291 23354
rect 10182 23296 10230 23352
rect 10286 23296 10291 23352
rect 10182 23291 10291 23296
rect 15377 23354 15443 23357
rect 21817 23354 21883 23357
rect 15377 23352 21883 23354
rect 15377 23296 15382 23352
rect 15438 23296 21822 23352
rect 21878 23296 21883 23352
rect 15377 23294 21883 23296
rect 15377 23291 15443 23294
rect 21817 23291 21883 23294
rect 10182 23085 10242 23291
rect 18689 23218 18755 23221
rect 10412 23216 18755 23218
rect 10412 23160 18694 23216
rect 18750 23160 18755 23216
rect 10412 23158 18755 23160
rect 10412 23085 10472 23158
rect 18689 23155 18755 23158
rect 33225 23218 33291 23221
rect 38745 23218 38811 23221
rect 33225 23216 38811 23218
rect 33225 23160 33230 23216
rect 33286 23160 38750 23216
rect 38806 23160 38811 23216
rect 33225 23158 38811 23160
rect 33225 23155 33291 23158
rect 38745 23155 38811 23158
rect 9765 23084 9831 23085
rect 9765 23082 9812 23084
rect 9720 23080 9812 23082
rect 9720 23024 9770 23080
rect 9720 23022 9812 23024
rect 9765 23020 9812 23022
rect 9876 23020 9882 23084
rect 10182 23080 10291 23085
rect 10182 23024 10230 23080
rect 10286 23024 10291 23080
rect 10182 23022 10291 23024
rect 9765 23019 9874 23020
rect 10225 23019 10291 23022
rect 10409 23080 10475 23085
rect 10409 23024 10414 23080
rect 10470 23024 10475 23080
rect 10409 23019 10475 23024
rect 10685 23084 10751 23085
rect 10685 23080 10732 23084
rect 10796 23082 10802 23084
rect 11973 23082 12039 23085
rect 18045 23082 18111 23085
rect 18638 23082 18644 23084
rect 10685 23024 10690 23080
rect 10685 23020 10732 23024
rect 10796 23022 10842 23082
rect 11973 23080 18644 23082
rect 11973 23024 11978 23080
rect 12034 23024 18050 23080
rect 18106 23024 18644 23080
rect 11973 23022 18644 23024
rect 10796 23020 10802 23022
rect 10685 23019 10751 23020
rect 11973 23019 12039 23022
rect 18045 23019 18111 23022
rect 18638 23020 18644 23022
rect 18708 23020 18714 23084
rect 28993 23082 29059 23085
rect 29637 23082 29703 23085
rect 36445 23082 36511 23085
rect 38009 23082 38075 23085
rect 28993 23080 36511 23082
rect 28993 23024 28998 23080
rect 29054 23024 29642 23080
rect 29698 23024 36450 23080
rect 36506 23024 36511 23080
rect 28993 23022 36511 23024
rect 28993 23019 29059 23022
rect 29637 23019 29703 23022
rect 36445 23019 36511 23022
rect 37966 23080 38075 23082
rect 37966 23024 38014 23080
rect 38070 23024 38075 23080
rect 37966 23019 38075 23024
rect 9814 22946 9874 23019
rect 13813 22948 13879 22949
rect 13813 22946 13860 22948
rect 9814 22944 13860 22946
rect 9814 22888 13818 22944
rect 9814 22886 13860 22888
rect 13813 22884 13860 22886
rect 13924 22884 13930 22948
rect 13813 22883 13879 22884
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 31845 22810 31911 22813
rect 35249 22810 35315 22813
rect 31845 22808 35315 22810
rect 31845 22752 31850 22808
rect 31906 22752 35254 22808
rect 35310 22752 35315 22808
rect 31845 22750 35315 22752
rect 31845 22747 31911 22750
rect 35249 22747 35315 22750
rect 11973 22676 12039 22677
rect 18781 22676 18847 22677
rect 11973 22674 12020 22676
rect 11928 22672 12020 22674
rect 11928 22616 11978 22672
rect 11928 22614 12020 22616
rect 11973 22612 12020 22614
rect 12084 22612 12090 22676
rect 18781 22672 18828 22676
rect 18892 22674 18898 22676
rect 36169 22674 36235 22677
rect 18781 22616 18786 22672
rect 18781 22612 18828 22616
rect 18892 22614 18938 22674
rect 22050 22672 36235 22674
rect 22050 22616 36174 22672
rect 36230 22616 36235 22672
rect 22050 22614 36235 22616
rect 18892 22612 18898 22614
rect 11973 22611 12039 22612
rect 18781 22611 18847 22612
rect 8201 22402 8267 22405
rect 9029 22402 9095 22405
rect 8201 22400 9095 22402
rect 8201 22344 8206 22400
rect 8262 22344 9034 22400
rect 9090 22344 9095 22400
rect 8201 22342 9095 22344
rect 8201 22339 8267 22342
rect 9029 22339 9095 22342
rect 14038 22340 14044 22404
rect 14108 22402 14114 22404
rect 14733 22402 14799 22405
rect 14108 22400 14799 22402
rect 14108 22344 14738 22400
rect 14794 22344 14799 22400
rect 14108 22342 14799 22344
rect 14108 22340 14114 22342
rect 14733 22339 14799 22342
rect 20437 22402 20503 22405
rect 21817 22402 21883 22405
rect 20437 22400 21883 22402
rect 20437 22344 20442 22400
rect 20498 22344 21822 22400
rect 21878 22344 21883 22400
rect 20437 22342 21883 22344
rect 20437 22339 20503 22342
rect 21817 22339 21883 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 8753 22266 8819 22269
rect 9581 22266 9647 22269
rect 8753 22264 9647 22266
rect 8753 22208 8758 22264
rect 8814 22208 9586 22264
rect 9642 22208 9647 22264
rect 8753 22206 9647 22208
rect 8753 22203 8819 22206
rect 9581 22203 9647 22206
rect 19885 22266 19951 22269
rect 21909 22266 21975 22269
rect 19885 22264 21975 22266
rect 19885 22208 19890 22264
rect 19946 22208 21914 22264
rect 21970 22208 21975 22264
rect 19885 22206 21975 22208
rect 19885 22203 19951 22206
rect 21909 22203 21975 22206
rect 10501 22130 10567 22133
rect 12801 22130 12867 22133
rect 14365 22130 14431 22133
rect 10501 22128 14431 22130
rect 10501 22072 10506 22128
rect 10562 22072 12806 22128
rect 12862 22072 14370 22128
rect 14426 22072 14431 22128
rect 10501 22070 14431 22072
rect 10501 22067 10567 22070
rect 12801 22067 12867 22070
rect 14365 22067 14431 22070
rect 20529 22130 20595 22133
rect 22050 22130 22110 22614
rect 36169 22611 36235 22614
rect 37966 22541 38026 23019
rect 24025 22538 24091 22541
rect 24158 22538 24164 22540
rect 24025 22536 24164 22538
rect 24025 22480 24030 22536
rect 24086 22480 24164 22536
rect 24025 22478 24164 22480
rect 24025 22475 24091 22478
rect 24158 22476 24164 22478
rect 24228 22476 24234 22540
rect 29269 22538 29335 22541
rect 30005 22538 30071 22541
rect 36118 22538 36124 22540
rect 29269 22536 36124 22538
rect 29269 22480 29274 22536
rect 29330 22480 30010 22536
rect 30066 22480 36124 22536
rect 29269 22478 36124 22480
rect 29269 22475 29335 22478
rect 30005 22475 30071 22478
rect 36118 22476 36124 22478
rect 36188 22476 36194 22540
rect 37966 22536 38075 22541
rect 37966 22480 38014 22536
rect 38070 22480 38075 22536
rect 37966 22478 38075 22480
rect 38009 22475 38075 22478
rect 29913 22404 29979 22405
rect 29862 22402 29868 22404
rect 29822 22342 29868 22402
rect 29932 22400 29979 22404
rect 29974 22344 29979 22400
rect 29862 22340 29868 22342
rect 29932 22340 29979 22344
rect 29913 22339 29979 22340
rect 31845 22402 31911 22405
rect 33501 22402 33567 22405
rect 31845 22400 33567 22402
rect 31845 22344 31850 22400
rect 31906 22344 33506 22400
rect 33562 22344 33567 22400
rect 31845 22342 33567 22344
rect 31845 22339 31911 22342
rect 33501 22339 33567 22342
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 23933 22266 23999 22269
rect 31017 22266 31083 22269
rect 23933 22264 31083 22266
rect 23933 22208 23938 22264
rect 23994 22208 31022 22264
rect 31078 22208 31083 22264
rect 23933 22206 31083 22208
rect 23933 22203 23999 22206
rect 31017 22203 31083 22206
rect 20529 22128 22110 22130
rect 20529 22072 20534 22128
rect 20590 22072 22110 22128
rect 20529 22070 22110 22072
rect 24761 22130 24827 22133
rect 27797 22130 27863 22133
rect 29821 22130 29887 22133
rect 24761 22128 29887 22130
rect 24761 22072 24766 22128
rect 24822 22072 27802 22128
rect 27858 22072 29826 22128
rect 29882 22072 29887 22128
rect 24761 22070 29887 22072
rect 20529 22067 20595 22070
rect 24761 22067 24827 22070
rect 27797 22067 27863 22070
rect 29821 22067 29887 22070
rect 4613 21994 4679 21997
rect 22001 21994 22067 21997
rect 22461 21996 22527 21997
rect 22461 21994 22508 21996
rect 4613 21992 22067 21994
rect 4613 21936 4618 21992
rect 4674 21936 22006 21992
rect 22062 21936 22067 21992
rect 4613 21934 22067 21936
rect 22416 21992 22508 21994
rect 22416 21936 22466 21992
rect 22416 21934 22508 21936
rect 4613 21931 4679 21934
rect 22001 21931 22067 21934
rect 22461 21932 22508 21934
rect 22572 21932 22578 21996
rect 22461 21931 22527 21932
rect 21214 21796 21220 21860
rect 21284 21858 21290 21860
rect 21357 21858 21423 21861
rect 21284 21856 21423 21858
rect 21284 21800 21362 21856
rect 21418 21800 21423 21856
rect 21284 21798 21423 21800
rect 21284 21796 21290 21798
rect 21357 21795 21423 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 35590 21727 35906 21728
rect 19793 21722 19859 21725
rect 21357 21722 21423 21725
rect 19793 21720 21423 21722
rect 19793 21664 19798 21720
rect 19854 21664 21362 21720
rect 21418 21664 21423 21720
rect 19793 21662 21423 21664
rect 19793 21659 19859 21662
rect 21357 21659 21423 21662
rect 3509 21586 3575 21589
rect 5165 21586 5231 21589
rect 3509 21584 5231 21586
rect 3509 21528 3514 21584
rect 3570 21528 5170 21584
rect 5226 21528 5231 21584
rect 3509 21526 5231 21528
rect 3509 21523 3575 21526
rect 5165 21523 5231 21526
rect 10501 21586 10567 21589
rect 13445 21586 13511 21589
rect 10501 21584 13511 21586
rect 10501 21528 10506 21584
rect 10562 21528 13450 21584
rect 13506 21528 13511 21584
rect 10501 21526 13511 21528
rect 10501 21523 10567 21526
rect 13445 21523 13511 21526
rect 17953 21586 18019 21589
rect 23381 21586 23447 21589
rect 27981 21588 28047 21589
rect 28993 21588 29059 21589
rect 27981 21586 28028 21588
rect 17953 21584 23447 21586
rect 17953 21528 17958 21584
rect 18014 21528 23386 21584
rect 23442 21528 23447 21584
rect 17953 21526 23447 21528
rect 27936 21584 28028 21586
rect 27936 21528 27986 21584
rect 27936 21526 28028 21528
rect 17953 21523 18019 21526
rect 23381 21523 23447 21526
rect 27981 21524 28028 21526
rect 28092 21524 28098 21588
rect 28942 21524 28948 21588
rect 29012 21586 29059 21588
rect 29012 21584 29104 21586
rect 29054 21528 29104 21584
rect 29012 21526 29104 21528
rect 29012 21524 29059 21526
rect 27981 21523 28047 21524
rect 28993 21523 29059 21524
rect 3601 21450 3667 21453
rect 7097 21450 7163 21453
rect 3601 21448 7163 21450
rect 3601 21392 3606 21448
rect 3662 21392 7102 21448
rect 7158 21392 7163 21448
rect 3601 21390 7163 21392
rect 3601 21387 3667 21390
rect 7097 21387 7163 21390
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 5717 21178 5783 21181
rect 6729 21178 6795 21181
rect 5717 21176 6795 21178
rect 5717 21120 5722 21176
rect 5778 21120 6734 21176
rect 6790 21120 6795 21176
rect 5717 21118 6795 21120
rect 5717 21115 5783 21118
rect 6729 21115 6795 21118
rect 4654 20980 4660 21044
rect 4724 21042 4730 21044
rect 4889 21042 4955 21045
rect 4724 21040 4955 21042
rect 4724 20984 4894 21040
rect 4950 20984 4955 21040
rect 4724 20982 4955 20984
rect 4724 20980 4730 20982
rect 4889 20979 4955 20982
rect 5073 21042 5139 21045
rect 7465 21042 7531 21045
rect 5073 21040 7531 21042
rect 5073 20984 5078 21040
rect 5134 20984 7470 21040
rect 7526 20984 7531 21040
rect 5073 20982 7531 20984
rect 5073 20979 5139 20982
rect 7465 20979 7531 20982
rect 8201 21042 8267 21045
rect 8334 21042 8340 21044
rect 8201 21040 8340 21042
rect 8201 20984 8206 21040
rect 8262 20984 8340 21040
rect 8201 20982 8340 20984
rect 8201 20979 8267 20982
rect 8334 20980 8340 20982
rect 8404 20980 8410 21044
rect 36302 20980 36308 21044
rect 36372 21042 36378 21044
rect 38101 21042 38167 21045
rect 36372 21040 38167 21042
rect 36372 20984 38106 21040
rect 38162 20984 38167 21040
rect 36372 20982 38167 20984
rect 36372 20980 36378 20982
rect 38101 20979 38167 20982
rect 3417 20906 3483 20909
rect 20805 20906 20871 20909
rect 27470 20906 27476 20908
rect 3417 20904 20871 20906
rect 3417 20848 3422 20904
rect 3478 20848 20810 20904
rect 20866 20848 20871 20904
rect 3417 20846 20871 20848
rect 3417 20843 3483 20846
rect 20805 20843 20871 20846
rect 21038 20846 27476 20906
rect 16062 20708 16068 20772
rect 16132 20770 16138 20772
rect 17493 20770 17559 20773
rect 16132 20768 17559 20770
rect 16132 20712 17498 20768
rect 17554 20712 17559 20768
rect 16132 20710 17559 20712
rect 16132 20708 16138 20710
rect 17493 20707 17559 20710
rect 20805 20770 20871 20773
rect 21038 20770 21098 20846
rect 27470 20844 27476 20846
rect 27540 20906 27546 20908
rect 28901 20906 28967 20909
rect 27540 20904 28967 20906
rect 27540 20848 28906 20904
rect 28962 20848 28967 20904
rect 27540 20846 28967 20848
rect 27540 20844 27546 20846
rect 28901 20843 28967 20846
rect 30465 20906 30531 20909
rect 34646 20906 34652 20908
rect 30465 20904 34652 20906
rect 30465 20848 30470 20904
rect 30526 20848 34652 20904
rect 30465 20846 34652 20848
rect 30465 20843 30531 20846
rect 34646 20844 34652 20846
rect 34716 20844 34722 20908
rect 22001 20772 22067 20773
rect 21950 20770 21956 20772
rect 20805 20768 21098 20770
rect 20805 20712 20810 20768
rect 20866 20712 21098 20768
rect 20805 20710 21098 20712
rect 21910 20710 21956 20770
rect 22020 20768 22067 20772
rect 22062 20712 22067 20768
rect 20805 20707 20871 20710
rect 21950 20708 21956 20710
rect 22020 20708 22067 20712
rect 23238 20708 23244 20772
rect 23308 20770 23314 20772
rect 23749 20770 23815 20773
rect 23308 20768 23815 20770
rect 23308 20712 23754 20768
rect 23810 20712 23815 20768
rect 23308 20710 23815 20712
rect 23308 20708 23314 20710
rect 22001 20707 22067 20708
rect 23749 20707 23815 20710
rect 24025 20770 24091 20773
rect 24342 20770 24348 20772
rect 24025 20768 24348 20770
rect 24025 20712 24030 20768
rect 24086 20712 24348 20768
rect 24025 20710 24348 20712
rect 24025 20707 24091 20710
rect 24342 20708 24348 20710
rect 24412 20708 24418 20772
rect 29821 20770 29887 20773
rect 30414 20770 30420 20772
rect 29821 20768 30420 20770
rect 29821 20712 29826 20768
rect 29882 20712 30420 20768
rect 29821 20710 30420 20712
rect 29821 20707 29887 20710
rect 30414 20708 30420 20710
rect 30484 20708 30490 20772
rect 34462 20708 34468 20772
rect 34532 20770 34538 20772
rect 34605 20770 34671 20773
rect 34532 20768 34671 20770
rect 34532 20712 34610 20768
rect 34666 20712 34671 20768
rect 34532 20710 34671 20712
rect 34532 20708 34538 20710
rect 34605 20707 34671 20710
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 5533 20634 5599 20637
rect 8569 20634 8635 20637
rect 5533 20632 8635 20634
rect 5533 20576 5538 20632
rect 5594 20576 8574 20632
rect 8630 20576 8635 20632
rect 5533 20574 8635 20576
rect 5533 20571 5599 20574
rect 8569 20571 8635 20574
rect 21398 20572 21404 20636
rect 21468 20634 21474 20636
rect 21817 20634 21883 20637
rect 21468 20632 21883 20634
rect 21468 20576 21822 20632
rect 21878 20576 21883 20632
rect 21468 20574 21883 20576
rect 21468 20572 21474 20574
rect 21817 20571 21883 20574
rect 25589 20634 25655 20637
rect 27613 20634 27679 20637
rect 25589 20632 27679 20634
rect 25589 20576 25594 20632
rect 25650 20576 27618 20632
rect 27674 20576 27679 20632
rect 25589 20574 27679 20576
rect 25589 20571 25655 20574
rect 27613 20571 27679 20574
rect 6361 20498 6427 20501
rect 7005 20498 7071 20501
rect 6361 20496 7071 20498
rect 6361 20440 6366 20496
rect 6422 20440 7010 20496
rect 7066 20440 7071 20496
rect 6361 20438 7071 20440
rect 6361 20435 6427 20438
rect 7005 20435 7071 20438
rect 16297 20498 16363 20501
rect 28717 20498 28783 20501
rect 16297 20496 28783 20498
rect 16297 20440 16302 20496
rect 16358 20440 28722 20496
rect 28778 20440 28783 20496
rect 16297 20438 28783 20440
rect 16297 20435 16363 20438
rect 28717 20435 28783 20438
rect 29729 20498 29795 20501
rect 31753 20498 31819 20501
rect 29729 20496 31819 20498
rect 29729 20440 29734 20496
rect 29790 20440 31758 20496
rect 31814 20440 31819 20496
rect 29729 20438 31819 20440
rect 29729 20435 29795 20438
rect 31753 20435 31819 20438
rect 5993 20362 6059 20365
rect 8109 20362 8175 20365
rect 5993 20360 8175 20362
rect 5993 20304 5998 20360
rect 6054 20304 8114 20360
rect 8170 20304 8175 20360
rect 5993 20302 8175 20304
rect 5993 20299 6059 20302
rect 8109 20299 8175 20302
rect 20478 20300 20484 20364
rect 20548 20362 20554 20364
rect 20621 20362 20687 20365
rect 20548 20360 20687 20362
rect 20548 20304 20626 20360
rect 20682 20304 20687 20360
rect 20548 20302 20687 20304
rect 20548 20300 20554 20302
rect 20621 20299 20687 20302
rect 25313 20362 25379 20365
rect 27245 20362 27311 20365
rect 25313 20360 27311 20362
rect 25313 20304 25318 20360
rect 25374 20304 27250 20360
rect 27306 20304 27311 20360
rect 25313 20302 27311 20304
rect 25313 20299 25379 20302
rect 27245 20299 27311 20302
rect 28574 20300 28580 20364
rect 28644 20362 28650 20364
rect 29453 20362 29519 20365
rect 28644 20360 29519 20362
rect 28644 20304 29458 20360
rect 29514 20304 29519 20360
rect 28644 20302 29519 20304
rect 28644 20300 28650 20302
rect 29453 20299 29519 20302
rect 17718 20164 17724 20228
rect 17788 20226 17794 20228
rect 20437 20226 20503 20229
rect 17788 20224 20503 20226
rect 17788 20168 20442 20224
rect 20498 20168 20503 20224
rect 17788 20166 20503 20168
rect 17788 20164 17794 20166
rect 20437 20163 20503 20166
rect 23105 20226 23171 20229
rect 27521 20226 27587 20229
rect 23105 20224 27587 20226
rect 23105 20168 23110 20224
rect 23166 20168 27526 20224
rect 27582 20168 27587 20224
rect 23105 20166 27587 20168
rect 23105 20163 23171 20166
rect 27521 20163 27587 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 6177 19956 6243 19957
rect 6126 19954 6132 19956
rect 6086 19894 6132 19954
rect 6196 19952 6243 19956
rect 6238 19896 6243 19952
rect 6126 19892 6132 19894
rect 6196 19892 6243 19896
rect 6177 19891 6243 19892
rect 13629 19954 13695 19957
rect 14917 19954 14983 19957
rect 15561 19954 15627 19957
rect 13629 19952 15627 19954
rect 13629 19896 13634 19952
rect 13690 19896 14922 19952
rect 14978 19896 15566 19952
rect 15622 19896 15627 19952
rect 13629 19894 15627 19896
rect 13629 19891 13695 19894
rect 14917 19891 14983 19894
rect 15561 19891 15627 19894
rect 21582 19892 21588 19956
rect 21652 19954 21658 19956
rect 21725 19954 21791 19957
rect 21652 19952 21791 19954
rect 21652 19896 21730 19952
rect 21786 19896 21791 19952
rect 21652 19894 21791 19896
rect 21652 19892 21658 19894
rect 21725 19891 21791 19894
rect 23197 19954 23263 19957
rect 28717 19954 28783 19957
rect 23197 19952 28783 19954
rect 23197 19896 23202 19952
rect 23258 19896 28722 19952
rect 28778 19896 28783 19952
rect 23197 19894 28783 19896
rect 23197 19891 23263 19894
rect 28717 19891 28783 19894
rect 38101 19954 38167 19957
rect 38510 19954 38516 19956
rect 38101 19952 38516 19954
rect 38101 19896 38106 19952
rect 38162 19896 38516 19952
rect 38101 19894 38516 19896
rect 38101 19891 38167 19894
rect 38510 19892 38516 19894
rect 38580 19892 38586 19956
rect 12985 19818 13051 19821
rect 14181 19818 14247 19821
rect 12985 19816 14247 19818
rect 12985 19760 12990 19816
rect 13046 19760 14186 19816
rect 14242 19760 14247 19816
rect 12985 19758 14247 19760
rect 12985 19755 13051 19758
rect 14181 19755 14247 19758
rect 14365 19818 14431 19821
rect 15285 19818 15351 19821
rect 14365 19816 15351 19818
rect 14365 19760 14370 19816
rect 14426 19760 15290 19816
rect 15346 19760 15351 19816
rect 14365 19758 15351 19760
rect 14365 19755 14431 19758
rect 15285 19755 15351 19758
rect 20069 19818 20135 19821
rect 24853 19818 24919 19821
rect 20069 19816 24919 19818
rect 20069 19760 20074 19816
rect 20130 19760 24858 19816
rect 24914 19760 24919 19816
rect 20069 19758 24919 19760
rect 20069 19755 20135 19758
rect 24853 19755 24919 19758
rect 30097 19818 30163 19821
rect 37181 19818 37247 19821
rect 30097 19816 37247 19818
rect 30097 19760 30102 19816
rect 30158 19760 37186 19816
rect 37242 19760 37247 19816
rect 30097 19758 37247 19760
rect 30097 19755 30163 19758
rect 37181 19755 37247 19758
rect 20529 19682 20595 19685
rect 21265 19682 21331 19685
rect 20529 19680 21331 19682
rect 20529 19624 20534 19680
rect 20590 19624 21270 19680
rect 21326 19624 21331 19680
rect 20529 19622 21331 19624
rect 20529 19619 20595 19622
rect 21265 19619 21331 19622
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 23105 19546 23171 19549
rect 23565 19546 23631 19549
rect 23105 19544 23631 19546
rect 23105 19488 23110 19544
rect 23166 19488 23570 19544
rect 23626 19488 23631 19544
rect 23105 19486 23631 19488
rect 23105 19483 23171 19486
rect 23565 19483 23631 19486
rect 21265 19410 21331 19413
rect 21909 19410 21975 19413
rect 21265 19408 21975 19410
rect 21265 19352 21270 19408
rect 21326 19352 21914 19408
rect 21970 19352 21975 19408
rect 21265 19350 21975 19352
rect 21265 19347 21331 19350
rect 21909 19347 21975 19350
rect 24301 19410 24367 19413
rect 27061 19410 27127 19413
rect 24301 19408 27127 19410
rect 24301 19352 24306 19408
rect 24362 19352 27066 19408
rect 27122 19352 27127 19408
rect 24301 19350 27127 19352
rect 24301 19347 24367 19350
rect 27061 19347 27127 19350
rect 30925 19410 30991 19413
rect 34697 19410 34763 19413
rect 30925 19408 34763 19410
rect 30925 19352 30930 19408
rect 30986 19352 34702 19408
rect 34758 19352 34763 19408
rect 30925 19350 34763 19352
rect 30925 19347 30991 19350
rect 34697 19347 34763 19350
rect 35382 19348 35388 19412
rect 35452 19410 35458 19412
rect 35525 19410 35591 19413
rect 35452 19408 35591 19410
rect 35452 19352 35530 19408
rect 35586 19352 35591 19408
rect 35452 19350 35591 19352
rect 35452 19348 35458 19350
rect 35525 19347 35591 19350
rect 21725 19274 21791 19277
rect 27705 19274 27771 19277
rect 21725 19272 27771 19274
rect 21725 19216 21730 19272
rect 21786 19216 27710 19272
rect 27766 19216 27771 19272
rect 21725 19214 27771 19216
rect 21725 19211 21791 19214
rect 27705 19211 27771 19214
rect 32806 19212 32812 19276
rect 32876 19274 32882 19276
rect 35893 19274 35959 19277
rect 32876 19272 35959 19274
rect 32876 19216 35898 19272
rect 35954 19216 35959 19272
rect 32876 19214 35959 19216
rect 32876 19212 32882 19214
rect 35893 19211 35959 19214
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 24393 19002 24459 19005
rect 28901 19002 28967 19005
rect 24393 19000 28967 19002
rect 24393 18944 24398 19000
rect 24454 18944 28906 19000
rect 28962 18944 28967 19000
rect 24393 18942 28967 18944
rect 24393 18939 24459 18942
rect 28901 18939 28967 18942
rect 22921 18866 22987 18869
rect 30230 18866 30236 18868
rect 22921 18864 30236 18866
rect 22921 18808 22926 18864
rect 22982 18808 30236 18864
rect 22921 18806 30236 18808
rect 22921 18803 22987 18806
rect 30230 18804 30236 18806
rect 30300 18866 30306 18868
rect 35893 18866 35959 18869
rect 30300 18864 35959 18866
rect 30300 18808 35898 18864
rect 35954 18808 35959 18864
rect 30300 18806 35959 18808
rect 30300 18804 30306 18806
rect 35893 18803 35959 18806
rect 21173 18730 21239 18733
rect 25957 18730 26023 18733
rect 27245 18730 27311 18733
rect 28717 18732 28783 18733
rect 28717 18730 28764 18732
rect 21173 18728 27311 18730
rect 21173 18672 21178 18728
rect 21234 18672 25962 18728
rect 26018 18672 27250 18728
rect 27306 18672 27311 18728
rect 21173 18670 27311 18672
rect 28672 18728 28764 18730
rect 28672 18672 28722 18728
rect 28672 18670 28764 18672
rect 21173 18667 21239 18670
rect 25957 18667 26023 18670
rect 27245 18667 27311 18670
rect 28717 18668 28764 18670
rect 28828 18668 28834 18732
rect 29678 18668 29684 18732
rect 29748 18730 29754 18732
rect 29913 18730 29979 18733
rect 29748 18728 29979 18730
rect 29748 18672 29918 18728
rect 29974 18672 29979 18728
rect 29748 18670 29979 18672
rect 29748 18668 29754 18670
rect 28717 18667 28783 18668
rect 29913 18667 29979 18670
rect 34278 18668 34284 18732
rect 34348 18730 34354 18732
rect 38285 18730 38351 18733
rect 34348 18728 38351 18730
rect 34348 18672 38290 18728
rect 38346 18672 38351 18728
rect 34348 18670 38351 18672
rect 34348 18668 34354 18670
rect 38285 18667 38351 18670
rect 21817 18594 21883 18597
rect 27429 18594 27495 18597
rect 28349 18596 28415 18597
rect 28349 18594 28396 18596
rect 21817 18592 27495 18594
rect 21817 18536 21822 18592
rect 21878 18536 27434 18592
rect 27490 18536 27495 18592
rect 21817 18534 27495 18536
rect 28308 18592 28396 18594
rect 28460 18594 28466 18596
rect 28758 18594 28764 18596
rect 28308 18536 28354 18592
rect 28308 18534 28396 18536
rect 21817 18531 21883 18534
rect 27429 18531 27495 18534
rect 28349 18532 28396 18534
rect 28460 18534 28764 18594
rect 28460 18532 28466 18534
rect 28758 18532 28764 18534
rect 28828 18532 28834 18596
rect 28349 18531 28415 18532
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 15561 18322 15627 18325
rect 18454 18322 18460 18324
rect 15561 18320 18460 18322
rect 15561 18264 15566 18320
rect 15622 18264 18460 18320
rect 15561 18262 18460 18264
rect 15561 18259 15627 18262
rect 18454 18260 18460 18262
rect 18524 18260 18530 18324
rect 26049 18322 26115 18325
rect 27613 18322 27679 18325
rect 34421 18324 34487 18325
rect 34421 18322 34468 18324
rect 26049 18320 27679 18322
rect 26049 18264 26054 18320
rect 26110 18264 27618 18320
rect 27674 18264 27679 18320
rect 26049 18262 27679 18264
rect 34376 18320 34468 18322
rect 34376 18264 34426 18320
rect 34376 18262 34468 18264
rect 26049 18259 26115 18262
rect 27613 18259 27679 18262
rect 34421 18260 34468 18262
rect 34532 18260 34538 18324
rect 34421 18259 34487 18260
rect 3693 18186 3759 18189
rect 4705 18186 4771 18189
rect 3693 18184 4771 18186
rect 3693 18128 3698 18184
rect 3754 18128 4710 18184
rect 4766 18128 4771 18184
rect 3693 18126 4771 18128
rect 3693 18123 3759 18126
rect 4705 18123 4771 18126
rect 30465 18186 30531 18189
rect 36302 18186 36308 18188
rect 30465 18184 36308 18186
rect 30465 18128 30470 18184
rect 30526 18128 36308 18184
rect 30465 18126 36308 18128
rect 30465 18123 30531 18126
rect 36302 18124 36308 18126
rect 36372 18124 36378 18188
rect 37958 17988 37964 18052
rect 38028 18050 38034 18052
rect 38285 18050 38351 18053
rect 38028 18048 38351 18050
rect 38028 17992 38290 18048
rect 38346 17992 38351 18048
rect 38028 17990 38351 17992
rect 38028 17988 38034 17990
rect 38285 17987 38351 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 8753 17914 8819 17917
rect 8886 17914 8892 17916
rect 8753 17912 8892 17914
rect 8753 17856 8758 17912
rect 8814 17856 8892 17912
rect 8753 17854 8892 17856
rect 8753 17851 8819 17854
rect 8886 17852 8892 17854
rect 8956 17852 8962 17916
rect 26141 17914 26207 17917
rect 27613 17914 27679 17917
rect 26141 17912 27679 17914
rect 26141 17856 26146 17912
rect 26202 17856 27618 17912
rect 27674 17856 27679 17912
rect 26141 17854 27679 17856
rect 26141 17851 26207 17854
rect 27613 17851 27679 17854
rect 30414 17852 30420 17916
rect 30484 17914 30490 17916
rect 31845 17914 31911 17917
rect 30484 17912 31911 17914
rect 30484 17856 31850 17912
rect 31906 17856 31911 17912
rect 30484 17854 31911 17856
rect 30484 17852 30490 17854
rect 31845 17851 31911 17854
rect 16941 17778 17007 17781
rect 17350 17778 17356 17780
rect 16941 17776 17356 17778
rect 16941 17720 16946 17776
rect 17002 17720 17356 17776
rect 16941 17718 17356 17720
rect 16941 17715 17007 17718
rect 17350 17716 17356 17718
rect 17420 17716 17426 17780
rect 26141 17778 26207 17781
rect 28022 17778 28028 17780
rect 26141 17776 28028 17778
rect 26141 17720 26146 17776
rect 26202 17720 28028 17776
rect 26141 17718 28028 17720
rect 26141 17715 26207 17718
rect 28022 17716 28028 17718
rect 28092 17716 28098 17780
rect 28993 17778 29059 17781
rect 29545 17778 29611 17781
rect 37273 17778 37339 17781
rect 28993 17776 37339 17778
rect 28993 17720 28998 17776
rect 29054 17720 29550 17776
rect 29606 17720 37278 17776
rect 37334 17720 37339 17776
rect 28993 17718 37339 17720
rect 28993 17715 29059 17718
rect 29545 17715 29611 17718
rect 37273 17715 37339 17718
rect 39389 17778 39455 17781
rect 40957 17778 41757 17808
rect 39389 17776 41757 17778
rect 39389 17720 39394 17776
rect 39450 17720 41757 17776
rect 39389 17718 41757 17720
rect 39389 17715 39455 17718
rect 40957 17688 41757 17718
rect 32765 17642 32831 17645
rect 34881 17642 34947 17645
rect 32765 17640 34947 17642
rect 32765 17584 32770 17640
rect 32826 17584 34886 17640
rect 34942 17584 34947 17640
rect 32765 17582 34947 17584
rect 32765 17579 32831 17582
rect 34881 17579 34947 17582
rect 31293 17506 31359 17509
rect 35341 17506 35407 17509
rect 31293 17504 35407 17506
rect 31293 17448 31298 17504
rect 31354 17448 35346 17504
rect 35402 17448 35407 17504
rect 31293 17446 35407 17448
rect 31293 17443 31359 17446
rect 35341 17443 35407 17446
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 22921 17370 22987 17373
rect 24526 17370 24532 17372
rect 22921 17368 24532 17370
rect 22921 17312 22926 17368
rect 22982 17312 24532 17368
rect 22921 17310 24532 17312
rect 22921 17307 22987 17310
rect 24526 17308 24532 17310
rect 24596 17370 24602 17372
rect 24669 17370 24735 17373
rect 27889 17370 27955 17373
rect 24596 17368 27955 17370
rect 24596 17312 24674 17368
rect 24730 17312 27894 17368
rect 27950 17312 27955 17368
rect 24596 17310 27955 17312
rect 24596 17308 24602 17310
rect 24669 17307 24735 17310
rect 27889 17307 27955 17310
rect 28349 17370 28415 17373
rect 28349 17368 28964 17370
rect 28349 17312 28354 17368
rect 28410 17312 28964 17368
rect 28349 17310 28964 17312
rect 28349 17307 28415 17310
rect 28904 17237 28964 17310
rect 28717 17234 28783 17237
rect 28717 17232 28826 17234
rect 28717 17176 28722 17232
rect 28778 17176 28826 17232
rect 28717 17171 28826 17176
rect 28901 17232 28967 17237
rect 28901 17176 28906 17232
rect 28962 17176 28967 17232
rect 28901 17171 28967 17176
rect 10726 17036 10732 17100
rect 10796 17098 10802 17100
rect 10869 17098 10935 17101
rect 11094 17098 11100 17100
rect 10796 17096 11100 17098
rect 10796 17040 10874 17096
rect 10930 17040 11100 17096
rect 10796 17038 11100 17040
rect 10796 17036 10802 17038
rect 10869 17035 10935 17038
rect 11094 17036 11100 17038
rect 11164 17036 11170 17100
rect 13813 17098 13879 17101
rect 14038 17098 14044 17100
rect 13813 17096 14044 17098
rect 13813 17040 13818 17096
rect 13874 17040 14044 17096
rect 13813 17038 14044 17040
rect 13813 17035 13879 17038
rect 14038 17036 14044 17038
rect 14108 17036 14114 17100
rect 15193 17098 15259 17101
rect 20110 17098 20116 17100
rect 15193 17096 20116 17098
rect 15193 17040 15198 17096
rect 15254 17040 20116 17096
rect 15193 17038 20116 17040
rect 15193 17035 15259 17038
rect 20110 17036 20116 17038
rect 20180 17036 20186 17100
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 22645 16826 22711 16829
rect 22921 16826 22987 16829
rect 22645 16824 22987 16826
rect 22645 16768 22650 16824
rect 22706 16768 22926 16824
rect 22982 16768 22987 16824
rect 22645 16766 22987 16768
rect 22645 16763 22711 16766
rect 22921 16763 22987 16766
rect 28766 16693 28826 17171
rect 32990 17036 32996 17100
rect 33060 17098 33066 17100
rect 33593 17098 33659 17101
rect 33060 17096 33659 17098
rect 33060 17040 33598 17096
rect 33654 17040 33659 17096
rect 33060 17038 33659 17040
rect 33060 17036 33066 17038
rect 33593 17035 33659 17038
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 10501 16692 10567 16693
rect 10501 16690 10548 16692
rect 10456 16688 10548 16690
rect 10456 16632 10506 16688
rect 10456 16630 10548 16632
rect 10501 16628 10548 16630
rect 10612 16628 10618 16692
rect 11697 16690 11763 16693
rect 11830 16690 11836 16692
rect 11697 16688 11836 16690
rect 11697 16632 11702 16688
rect 11758 16632 11836 16688
rect 11697 16630 11836 16632
rect 10501 16627 10567 16628
rect 11697 16627 11763 16630
rect 11830 16628 11836 16630
rect 11900 16628 11906 16692
rect 20437 16690 20503 16693
rect 27337 16690 27403 16693
rect 20437 16688 27403 16690
rect 20437 16632 20442 16688
rect 20498 16632 27342 16688
rect 27398 16632 27403 16688
rect 20437 16630 27403 16632
rect 28766 16688 28875 16693
rect 28766 16632 28814 16688
rect 28870 16632 28875 16688
rect 28766 16630 28875 16632
rect 20437 16627 20503 16630
rect 27337 16627 27403 16630
rect 28809 16627 28875 16630
rect 31569 16690 31635 16693
rect 31886 16690 31892 16692
rect 31569 16688 31892 16690
rect 31569 16632 31574 16688
rect 31630 16632 31892 16688
rect 31569 16630 31892 16632
rect 31569 16627 31635 16630
rect 31886 16628 31892 16630
rect 31956 16690 31962 16692
rect 32581 16690 32647 16693
rect 31956 16688 32647 16690
rect 31956 16632 32586 16688
rect 32642 16632 32647 16688
rect 31956 16630 32647 16632
rect 31956 16628 31962 16630
rect 32581 16627 32647 16630
rect 20805 16554 20871 16557
rect 23381 16554 23447 16557
rect 20805 16552 23447 16554
rect 20805 16496 20810 16552
rect 20866 16496 23386 16552
rect 23442 16496 23447 16552
rect 20805 16494 23447 16496
rect 20805 16491 20871 16494
rect 23381 16491 23447 16494
rect 27521 16554 27587 16557
rect 28625 16554 28691 16557
rect 36813 16554 36879 16557
rect 27521 16552 28691 16554
rect 27521 16496 27526 16552
rect 27582 16496 28630 16552
rect 28686 16496 28691 16552
rect 27521 16494 28691 16496
rect 27521 16491 27587 16494
rect 28625 16491 28691 16494
rect 34286 16552 36879 16554
rect 34286 16496 36818 16552
rect 36874 16496 36879 16552
rect 34286 16494 36879 16496
rect 30373 16418 30439 16421
rect 30598 16418 30604 16420
rect 30373 16416 30604 16418
rect 30373 16360 30378 16416
rect 30434 16360 30604 16416
rect 30373 16358 30604 16360
rect 30373 16355 30439 16358
rect 30598 16356 30604 16358
rect 30668 16418 30674 16420
rect 34286 16418 34346 16494
rect 36813 16491 36879 16494
rect 30668 16358 34346 16418
rect 37273 16418 37339 16421
rect 40957 16418 41757 16448
rect 37273 16416 41757 16418
rect 37273 16360 37278 16416
rect 37334 16360 41757 16416
rect 37273 16358 41757 16360
rect 30668 16356 30674 16358
rect 37273 16355 37339 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 40957 16328 41757 16358
rect 35590 16287 35906 16288
rect 30373 16282 30439 16285
rect 30649 16282 30715 16285
rect 30373 16280 30715 16282
rect 30373 16224 30378 16280
rect 30434 16224 30654 16280
rect 30710 16224 30715 16280
rect 30373 16222 30715 16224
rect 30373 16219 30439 16222
rect 30649 16219 30715 16222
rect 30281 16146 30347 16149
rect 34421 16146 34487 16149
rect 35157 16146 35223 16149
rect 30281 16144 35223 16146
rect 30281 16088 30286 16144
rect 30342 16088 34426 16144
rect 34482 16088 35162 16144
rect 35218 16088 35223 16144
rect 30281 16086 35223 16088
rect 30281 16083 30347 16086
rect 34421 16083 34487 16086
rect 35157 16083 35223 16086
rect 12801 16012 12867 16013
rect 12750 15948 12756 16012
rect 12820 16010 12867 16012
rect 12820 16008 12912 16010
rect 12862 15952 12912 16008
rect 12820 15950 12912 15952
rect 12820 15948 12867 15950
rect 12801 15947 12867 15948
rect 10869 15876 10935 15877
rect 10869 15874 10916 15876
rect 10824 15872 10916 15874
rect 10824 15816 10874 15872
rect 10824 15814 10916 15816
rect 10869 15812 10916 15814
rect 10980 15812 10986 15876
rect 22001 15874 22067 15877
rect 22318 15874 22324 15876
rect 22001 15872 22324 15874
rect 22001 15816 22006 15872
rect 22062 15816 22324 15872
rect 22001 15814 22324 15816
rect 10869 15811 10935 15812
rect 22001 15811 22067 15814
rect 22318 15812 22324 15814
rect 22388 15812 22394 15876
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 22093 15604 22159 15605
rect 22093 15600 22140 15604
rect 22204 15602 22210 15604
rect 22093 15544 22098 15600
rect 22093 15540 22140 15544
rect 22204 15542 22250 15602
rect 22204 15540 22210 15542
rect 22093 15539 22159 15540
rect 31201 15466 31267 15469
rect 31477 15466 31543 15469
rect 31201 15464 31543 15466
rect 31201 15408 31206 15464
rect 31262 15408 31482 15464
rect 31538 15408 31543 15464
rect 31201 15406 31543 15408
rect 31201 15403 31267 15406
rect 31477 15403 31543 15406
rect 29085 15330 29151 15333
rect 27662 15328 29151 15330
rect 27662 15272 29090 15328
rect 29146 15272 29151 15328
rect 27662 15270 29151 15272
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 18638 15132 18644 15196
rect 18708 15194 18714 15196
rect 20110 15194 20116 15196
rect 18708 15134 20116 15194
rect 18708 15132 18714 15134
rect 20110 15132 20116 15134
rect 20180 15132 20186 15196
rect 25814 15132 25820 15196
rect 25884 15194 25890 15196
rect 27662 15194 27722 15270
rect 29085 15267 29151 15270
rect 36905 15330 36971 15333
rect 37406 15330 37412 15332
rect 36905 15328 37412 15330
rect 36905 15272 36910 15328
rect 36966 15272 37412 15328
rect 36905 15270 37412 15272
rect 36905 15267 36971 15270
rect 37406 15268 37412 15270
rect 37476 15268 37482 15332
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 25884 15134 27722 15194
rect 25884 15132 25890 15134
rect 24669 15058 24735 15061
rect 25630 15058 25636 15060
rect 24669 15056 25636 15058
rect 24669 15000 24674 15056
rect 24730 15000 25636 15056
rect 24669 14998 25636 15000
rect 24669 14995 24735 14998
rect 25630 14996 25636 14998
rect 25700 15058 25706 15060
rect 27429 15058 27495 15061
rect 25700 15056 27495 15058
rect 25700 15000 27434 15056
rect 27490 15000 27495 15056
rect 25700 14998 27495 15000
rect 25700 14996 25706 14998
rect 27429 14995 27495 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19793 14650 19859 14653
rect 19926 14650 19932 14652
rect 19793 14648 19932 14650
rect 19793 14592 19798 14648
rect 19854 14592 19932 14648
rect 19793 14590 19932 14592
rect 19793 14587 19859 14590
rect 19926 14588 19932 14590
rect 19996 14588 20002 14652
rect 21766 14588 21772 14652
rect 21836 14650 21842 14652
rect 22185 14650 22251 14653
rect 21836 14648 22251 14650
rect 21836 14592 22190 14648
rect 22246 14592 22251 14648
rect 21836 14590 22251 14592
rect 21836 14588 21842 14590
rect 22185 14587 22251 14590
rect 27981 14650 28047 14653
rect 28533 14650 28599 14653
rect 27981 14648 28599 14650
rect 27981 14592 27986 14648
rect 28042 14592 28538 14648
rect 28594 14592 28599 14648
rect 27981 14590 28599 14592
rect 27981 14587 28047 14590
rect 28533 14587 28599 14590
rect 7557 14514 7623 14517
rect 8017 14514 8083 14517
rect 8753 14514 8819 14517
rect 7557 14512 8819 14514
rect 7557 14456 7562 14512
rect 7618 14456 8022 14512
rect 8078 14456 8758 14512
rect 8814 14456 8819 14512
rect 7557 14454 8819 14456
rect 7557 14451 7623 14454
rect 8017 14451 8083 14454
rect 8753 14451 8819 14454
rect 20161 14514 20227 14517
rect 23933 14514 23999 14517
rect 20161 14512 23999 14514
rect 20161 14456 20166 14512
rect 20222 14456 23938 14512
rect 23994 14456 23999 14512
rect 20161 14454 23999 14456
rect 20161 14451 20227 14454
rect 23933 14451 23999 14454
rect 25037 14512 25103 14517
rect 25037 14456 25042 14512
rect 25098 14456 25103 14512
rect 25037 14451 25103 14456
rect 27797 14514 27863 14517
rect 28901 14514 28967 14517
rect 27797 14512 28967 14514
rect 27797 14456 27802 14512
rect 27858 14456 28906 14512
rect 28962 14456 28967 14512
rect 27797 14454 28967 14456
rect 27797 14451 27863 14454
rect 28901 14451 28967 14454
rect 25040 14378 25100 14451
rect 25313 14378 25379 14381
rect 25040 14376 25379 14378
rect 25040 14320 25318 14376
rect 25374 14320 25379 14376
rect 25040 14318 25379 14320
rect 25313 14315 25379 14318
rect 28073 14378 28139 14381
rect 28901 14378 28967 14381
rect 28073 14376 28967 14378
rect 28073 14320 28078 14376
rect 28134 14320 28906 14376
rect 28962 14320 28967 14376
rect 28073 14318 28967 14320
rect 28073 14315 28139 14318
rect 28901 14315 28967 14318
rect 30465 14378 30531 14381
rect 30966 14378 30972 14380
rect 30465 14376 30972 14378
rect 30465 14320 30470 14376
rect 30526 14320 30972 14376
rect 30465 14318 30972 14320
rect 30465 14315 30531 14318
rect 30966 14316 30972 14318
rect 31036 14316 31042 14380
rect 22369 14242 22435 14245
rect 26509 14242 26575 14245
rect 22369 14240 26575 14242
rect 22369 14184 22374 14240
rect 22430 14184 26514 14240
rect 26570 14184 26575 14240
rect 22369 14182 26575 14184
rect 22369 14179 22435 14182
rect 26509 14179 26575 14182
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 23933 14108 23999 14109
rect 23933 14106 23980 14108
rect 23888 14104 23980 14106
rect 24044 14106 24050 14108
rect 24485 14106 24551 14109
rect 27061 14108 27127 14109
rect 25814 14106 25820 14108
rect 24044 14104 25820 14106
rect 23888 14048 23938 14104
rect 24044 14048 24490 14104
rect 24546 14048 25820 14104
rect 23888 14046 23980 14048
rect 23933 14044 23980 14046
rect 24044 14046 25820 14048
rect 24044 14044 24050 14046
rect 23933 14043 23999 14044
rect 24485 14043 24551 14046
rect 25814 14044 25820 14046
rect 25884 14044 25890 14108
rect 27061 14106 27108 14108
rect 27016 14104 27108 14106
rect 27016 14048 27066 14104
rect 27016 14046 27108 14048
rect 27061 14044 27108 14046
rect 27172 14044 27178 14108
rect 27705 14106 27771 14109
rect 28901 14106 28967 14109
rect 27705 14104 28967 14106
rect 27705 14048 27710 14104
rect 27766 14048 28906 14104
rect 28962 14048 28967 14104
rect 27705 14046 28967 14048
rect 27061 14043 27127 14044
rect 27705 14043 27771 14046
rect 28901 14043 28967 14046
rect 24669 13970 24735 13973
rect 27654 13970 27660 13972
rect 24669 13968 27660 13970
rect 24669 13912 24674 13968
rect 24730 13912 27660 13968
rect 24669 13910 27660 13912
rect 24669 13907 24735 13910
rect 27654 13908 27660 13910
rect 27724 13908 27730 13972
rect 25446 13772 25452 13836
rect 25516 13834 25522 13836
rect 28574 13834 28580 13836
rect 25516 13774 28580 13834
rect 25516 13772 25522 13774
rect 28574 13772 28580 13774
rect 28644 13772 28650 13836
rect 28942 13636 28948 13700
rect 29012 13698 29018 13700
rect 29085 13698 29151 13701
rect 29012 13696 29151 13698
rect 29012 13640 29090 13696
rect 29146 13640 29151 13696
rect 29012 13638 29151 13640
rect 29012 13636 29018 13638
rect 29085 13635 29151 13638
rect 32213 13698 32279 13701
rect 32438 13698 32444 13700
rect 32213 13696 32444 13698
rect 32213 13640 32218 13696
rect 32274 13640 32444 13696
rect 32213 13638 32444 13640
rect 32213 13635 32279 13638
rect 32438 13636 32444 13638
rect 32508 13636 32514 13700
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 31845 13564 31911 13565
rect 31845 13562 31892 13564
rect 31800 13560 31892 13562
rect 31800 13504 31850 13560
rect 31800 13502 31892 13504
rect 31845 13500 31892 13502
rect 31956 13500 31962 13564
rect 31845 13499 31954 13500
rect 20713 13426 20779 13429
rect 22737 13426 22803 13429
rect 20713 13424 22803 13426
rect 20713 13368 20718 13424
rect 20774 13368 22742 13424
rect 22798 13368 22803 13424
rect 20713 13366 22803 13368
rect 31894 13426 31954 13499
rect 32397 13426 32463 13429
rect 31894 13424 32463 13426
rect 31894 13368 32402 13424
rect 32458 13368 32463 13424
rect 31894 13366 32463 13368
rect 20713 13363 20779 13366
rect 22737 13363 22803 13366
rect 32397 13363 32463 13366
rect 22093 13290 22159 13293
rect 26233 13290 26299 13293
rect 22093 13288 26299 13290
rect 22093 13232 22098 13288
rect 22154 13232 26238 13288
rect 26294 13232 26299 13288
rect 22093 13230 26299 13232
rect 22093 13227 22159 13230
rect 26233 13227 26299 13230
rect 19701 13154 19767 13157
rect 22001 13154 22067 13157
rect 34697 13156 34763 13157
rect 34646 13154 34652 13156
rect 19701 13152 22067 13154
rect 19701 13096 19706 13152
rect 19762 13096 22006 13152
rect 22062 13096 22067 13152
rect 19701 13094 22067 13096
rect 34606 13094 34652 13154
rect 34716 13152 34763 13156
rect 34758 13096 34763 13152
rect 19701 13091 19767 13094
rect 22001 13091 22067 13094
rect 34646 13092 34652 13094
rect 34716 13092 34763 13096
rect 34697 13091 34763 13092
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 30189 13018 30255 13021
rect 30833 13018 30899 13021
rect 30189 13016 30899 13018
rect 30189 12960 30194 13016
rect 30250 12960 30838 13016
rect 30894 12960 30899 13016
rect 30189 12958 30899 12960
rect 30189 12955 30255 12958
rect 30833 12955 30899 12958
rect 4889 12882 4955 12885
rect 7465 12882 7531 12885
rect 4889 12880 7531 12882
rect 4889 12824 4894 12880
rect 4950 12824 7470 12880
rect 7526 12824 7531 12880
rect 4889 12822 7531 12824
rect 4889 12819 4955 12822
rect 7465 12819 7531 12822
rect 17125 12882 17191 12885
rect 17585 12882 17651 12885
rect 17125 12880 17651 12882
rect 17125 12824 17130 12880
rect 17186 12824 17590 12880
rect 17646 12824 17651 12880
rect 17125 12822 17651 12824
rect 17125 12819 17191 12822
rect 17585 12819 17651 12822
rect 22737 12882 22803 12885
rect 33685 12882 33751 12885
rect 22737 12880 33751 12882
rect 22737 12824 22742 12880
rect 22798 12824 33690 12880
rect 33746 12824 33751 12880
rect 22737 12822 33751 12824
rect 22737 12819 22803 12822
rect 33685 12819 33751 12822
rect 5901 12746 5967 12749
rect 6821 12746 6887 12749
rect 8937 12746 9003 12749
rect 5901 12744 9003 12746
rect 5901 12688 5906 12744
rect 5962 12688 6826 12744
rect 6882 12688 8942 12744
rect 8998 12688 9003 12744
rect 5901 12686 9003 12688
rect 5901 12683 5967 12686
rect 6821 12683 6887 12686
rect 8937 12683 9003 12686
rect 18689 12746 18755 12749
rect 29729 12746 29795 12749
rect 18689 12744 29795 12746
rect 18689 12688 18694 12744
rect 18750 12688 29734 12744
rect 29790 12688 29795 12744
rect 18689 12686 29795 12688
rect 18689 12683 18755 12686
rect 29729 12683 29795 12686
rect 30465 12746 30531 12749
rect 34278 12746 34284 12748
rect 30465 12744 34284 12746
rect 30465 12688 30470 12744
rect 30526 12688 34284 12744
rect 30465 12686 34284 12688
rect 30465 12683 30531 12686
rect 34278 12684 34284 12686
rect 34348 12684 34354 12748
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 23657 12474 23723 12477
rect 23841 12474 23907 12477
rect 23657 12472 23907 12474
rect 23657 12416 23662 12472
rect 23718 12416 23846 12472
rect 23902 12416 23907 12472
rect 23657 12414 23907 12416
rect 23657 12411 23723 12414
rect 23841 12411 23907 12414
rect 30230 12412 30236 12476
rect 30300 12474 30306 12476
rect 30465 12474 30531 12477
rect 30300 12472 30531 12474
rect 30300 12416 30470 12472
rect 30526 12416 30531 12472
rect 30300 12414 30531 12416
rect 30300 12412 30306 12414
rect 30465 12411 30531 12414
rect 24342 12276 24348 12340
rect 24412 12338 24418 12340
rect 29729 12338 29795 12341
rect 32990 12338 32996 12340
rect 24412 12336 32996 12338
rect 24412 12280 29734 12336
rect 29790 12280 32996 12336
rect 24412 12278 32996 12280
rect 24412 12276 24418 12278
rect 29729 12275 29795 12278
rect 32990 12276 32996 12278
rect 33060 12276 33066 12340
rect 33501 12202 33567 12205
rect 38193 12202 38259 12205
rect 33501 12200 38259 12202
rect 33501 12144 33506 12200
rect 33562 12144 38198 12200
rect 38254 12144 38259 12200
rect 33501 12142 38259 12144
rect 33501 12139 33567 12142
rect 38193 12139 38259 12142
rect 11830 12004 11836 12068
rect 11900 12066 11906 12068
rect 12893 12066 12959 12069
rect 11900 12064 12959 12066
rect 11900 12008 12898 12064
rect 12954 12008 12959 12064
rect 11900 12006 12959 12008
rect 11900 12004 11906 12006
rect 12893 12003 12959 12006
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 22001 11932 22067 11933
rect 19374 11868 19380 11932
rect 19444 11930 19450 11932
rect 21950 11930 21956 11932
rect 19444 11870 21956 11930
rect 22020 11928 22067 11932
rect 22062 11872 22067 11928
rect 19444 11868 19450 11870
rect 21950 11868 21956 11870
rect 22020 11868 22067 11872
rect 22001 11867 22067 11868
rect 24485 11930 24551 11933
rect 28349 11930 28415 11933
rect 24485 11928 28415 11930
rect 24485 11872 24490 11928
rect 24546 11872 28354 11928
rect 28410 11872 28415 11928
rect 24485 11870 28415 11872
rect 24485 11867 24551 11870
rect 28349 11867 28415 11870
rect 22277 11794 22343 11797
rect 22502 11794 22508 11796
rect 22277 11792 22508 11794
rect 22277 11736 22282 11792
rect 22338 11736 22508 11792
rect 22277 11734 22508 11736
rect 22277 11731 22343 11734
rect 22502 11732 22508 11734
rect 22572 11732 22578 11796
rect 25446 11732 25452 11796
rect 25516 11794 25522 11796
rect 25589 11794 25655 11797
rect 33593 11796 33659 11797
rect 25516 11792 25655 11794
rect 25516 11736 25594 11792
rect 25650 11736 25655 11792
rect 25516 11734 25655 11736
rect 25516 11732 25522 11734
rect 25589 11731 25655 11734
rect 32254 11732 32260 11796
rect 32324 11794 32330 11796
rect 33542 11794 33548 11796
rect 32324 11734 33548 11794
rect 33612 11792 33659 11796
rect 33654 11736 33659 11792
rect 32324 11732 32330 11734
rect 33542 11732 33548 11734
rect 33612 11732 33659 11736
rect 33593 11731 33659 11732
rect 34329 11794 34395 11797
rect 34789 11794 34855 11797
rect 34329 11792 34855 11794
rect 34329 11736 34334 11792
rect 34390 11736 34794 11792
rect 34850 11736 34855 11792
rect 34329 11734 34855 11736
rect 34329 11731 34395 11734
rect 34789 11731 34855 11734
rect 19517 11658 19583 11661
rect 26877 11658 26943 11661
rect 36813 11658 36879 11661
rect 19517 11656 26943 11658
rect 19517 11600 19522 11656
rect 19578 11600 26882 11656
rect 26938 11600 26943 11656
rect 19517 11598 26943 11600
rect 19517 11595 19583 11598
rect 26877 11595 26943 11598
rect 31710 11656 36879 11658
rect 31710 11600 36818 11656
rect 36874 11600 36879 11656
rect 31710 11598 36879 11600
rect 23105 11522 23171 11525
rect 25313 11522 25379 11525
rect 27705 11522 27771 11525
rect 23105 11520 27771 11522
rect 23105 11464 23110 11520
rect 23166 11464 25318 11520
rect 25374 11464 27710 11520
rect 27766 11464 27771 11520
rect 23105 11462 27771 11464
rect 23105 11459 23171 11462
rect 25313 11459 25379 11462
rect 27705 11459 27771 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 28073 11386 28139 11389
rect 31710 11386 31770 11598
rect 36813 11595 36879 11598
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 22050 11384 31770 11386
rect 22050 11328 28078 11384
rect 28134 11328 31770 11384
rect 22050 11326 31770 11328
rect 18505 11250 18571 11253
rect 22050 11250 22110 11326
rect 28073 11323 28139 11326
rect 18505 11248 22110 11250
rect 18505 11192 18510 11248
rect 18566 11192 22110 11248
rect 18505 11190 22110 11192
rect 18505 11187 18571 11190
rect 24710 11188 24716 11252
rect 24780 11250 24786 11252
rect 25998 11250 26004 11252
rect 24780 11190 26004 11250
rect 24780 11188 24786 11190
rect 25998 11188 26004 11190
rect 26068 11188 26074 11252
rect 29545 11250 29611 11253
rect 30782 11250 30788 11252
rect 29545 11248 30788 11250
rect 29545 11192 29550 11248
rect 29606 11192 30788 11248
rect 29545 11190 30788 11192
rect 29545 11187 29611 11190
rect 30782 11188 30788 11190
rect 30852 11188 30858 11252
rect 30925 11250 30991 11253
rect 34973 11250 35039 11253
rect 30925 11248 35039 11250
rect 30925 11192 30930 11248
rect 30986 11192 34978 11248
rect 35034 11192 35039 11248
rect 30925 11190 35039 11192
rect 30925 11187 30991 11190
rect 34973 11187 35039 11190
rect 24853 11114 24919 11117
rect 25405 11114 25471 11117
rect 32857 11114 32923 11117
rect 24853 11112 32923 11114
rect 24853 11056 24858 11112
rect 24914 11056 25410 11112
rect 25466 11056 32862 11112
rect 32918 11056 32923 11112
rect 24853 11054 32923 11056
rect 24853 11051 24919 11054
rect 25405 11051 25471 11054
rect 32857 11051 32923 11054
rect 33593 11114 33659 11117
rect 36629 11114 36695 11117
rect 33593 11112 36695 11114
rect 33593 11056 33598 11112
rect 33654 11056 36634 11112
rect 36690 11056 36695 11112
rect 33593 11054 36695 11056
rect 33593 11051 33659 11054
rect 36629 11051 36695 11054
rect 0 10978 800 11008
rect 1853 10978 1919 10981
rect 0 10976 1919 10978
rect 0 10920 1858 10976
rect 1914 10920 1919 10976
rect 0 10918 1919 10920
rect 0 10888 800 10918
rect 1853 10915 1919 10918
rect 29453 10978 29519 10981
rect 34881 10978 34947 10981
rect 29453 10976 34947 10978
rect 29453 10920 29458 10976
rect 29514 10920 34886 10976
rect 34942 10920 34947 10976
rect 29453 10918 34947 10920
rect 29453 10915 29519 10918
rect 34881 10915 34947 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 35590 10847 35906 10848
rect 25814 10780 25820 10844
rect 25884 10842 25890 10844
rect 26049 10842 26115 10845
rect 25884 10840 26115 10842
rect 25884 10784 26054 10840
rect 26110 10784 26115 10840
rect 25884 10782 26115 10784
rect 25884 10780 25890 10782
rect 26049 10779 26115 10782
rect 20805 10706 20871 10709
rect 21357 10706 21423 10709
rect 21582 10706 21588 10708
rect 20805 10704 21588 10706
rect 20805 10648 20810 10704
rect 20866 10648 21362 10704
rect 21418 10648 21588 10704
rect 20805 10646 21588 10648
rect 20805 10643 20871 10646
rect 21357 10643 21423 10646
rect 21582 10644 21588 10646
rect 21652 10644 21658 10708
rect 21817 10706 21883 10709
rect 25037 10706 25103 10709
rect 25313 10706 25379 10709
rect 21817 10704 25379 10706
rect 21817 10648 21822 10704
rect 21878 10648 25042 10704
rect 25098 10648 25318 10704
rect 25374 10648 25379 10704
rect 21817 10646 25379 10648
rect 21817 10643 21883 10646
rect 25037 10643 25103 10646
rect 25313 10643 25379 10646
rect 22921 10570 22987 10573
rect 27613 10570 27679 10573
rect 28901 10570 28967 10573
rect 22921 10568 28967 10570
rect 22921 10512 22926 10568
rect 22982 10512 27618 10568
rect 27674 10512 28906 10568
rect 28962 10512 28967 10568
rect 22921 10510 28967 10512
rect 22921 10507 22987 10510
rect 27613 10507 27679 10510
rect 28901 10507 28967 10510
rect 31201 10570 31267 10573
rect 31569 10570 31635 10573
rect 31201 10568 31635 10570
rect 31201 10512 31206 10568
rect 31262 10512 31574 10568
rect 31630 10512 31635 10568
rect 31201 10510 31635 10512
rect 31201 10507 31267 10510
rect 31569 10507 31635 10510
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 5717 10300 5783 10301
rect 5717 10298 5764 10300
rect 5672 10296 5764 10298
rect 5672 10240 5722 10296
rect 5672 10238 5764 10240
rect 5717 10236 5764 10238
rect 5828 10236 5834 10300
rect 16849 10298 16915 10301
rect 16982 10298 16988 10300
rect 16849 10296 16988 10298
rect 16849 10240 16854 10296
rect 16910 10240 16988 10296
rect 16849 10238 16988 10240
rect 5717 10235 5783 10236
rect 16849 10235 16915 10238
rect 16982 10236 16988 10238
rect 17052 10236 17058 10300
rect 17217 10162 17283 10165
rect 29545 10162 29611 10165
rect 30598 10162 30604 10164
rect 17217 10160 30604 10162
rect 17217 10104 17222 10160
rect 17278 10104 29550 10160
rect 29606 10104 30604 10160
rect 17217 10102 30604 10104
rect 17217 10099 17283 10102
rect 29545 10099 29611 10102
rect 30598 10100 30604 10102
rect 30668 10100 30674 10164
rect 19793 10026 19859 10029
rect 25589 10028 25655 10029
rect 25589 10026 25636 10028
rect 19793 10024 25636 10026
rect 19793 9968 19798 10024
rect 19854 9968 25594 10024
rect 19793 9966 25636 9968
rect 19793 9963 19859 9966
rect 25589 9964 25636 9966
rect 25700 9964 25706 10028
rect 25589 9963 25655 9964
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 19374 9754 19380 9756
rect 16438 9694 19380 9754
rect 16438 9621 16498 9694
rect 19374 9692 19380 9694
rect 19444 9692 19450 9756
rect 22829 9754 22895 9757
rect 26509 9754 26575 9757
rect 22829 9752 26575 9754
rect 22829 9696 22834 9752
rect 22890 9696 26514 9752
rect 26570 9696 26575 9752
rect 22829 9694 26575 9696
rect 22829 9691 22895 9694
rect 26509 9691 26575 9694
rect 30833 9754 30899 9757
rect 34462 9754 34468 9756
rect 30833 9752 34468 9754
rect 30833 9696 30838 9752
rect 30894 9696 34468 9752
rect 30833 9694 34468 9696
rect 30833 9691 30899 9694
rect 34462 9692 34468 9694
rect 34532 9754 34538 9756
rect 35065 9754 35131 9757
rect 34532 9752 35131 9754
rect 34532 9696 35070 9752
rect 35126 9696 35131 9752
rect 34532 9694 35131 9696
rect 34532 9692 34538 9694
rect 35065 9691 35131 9694
rect 16438 9616 16547 9621
rect 16438 9560 16486 9616
rect 16542 9560 16547 9616
rect 16438 9558 16547 9560
rect 16481 9555 16547 9558
rect 20805 9618 20871 9621
rect 25497 9618 25563 9621
rect 29085 9618 29151 9621
rect 20805 9616 21098 9618
rect 20805 9560 20810 9616
rect 20866 9560 21098 9616
rect 20805 9558 21098 9560
rect 20805 9555 20871 9558
rect 16246 9420 16252 9484
rect 16316 9482 16322 9484
rect 20897 9482 20963 9485
rect 16316 9480 20963 9482
rect 16316 9424 20902 9480
rect 20958 9424 20963 9480
rect 16316 9422 20963 9424
rect 21038 9482 21098 9558
rect 25497 9616 29151 9618
rect 25497 9560 25502 9616
rect 25558 9560 29090 9616
rect 29146 9560 29151 9616
rect 25497 9558 29151 9560
rect 25497 9555 25563 9558
rect 29085 9555 29151 9558
rect 30966 9556 30972 9620
rect 31036 9618 31042 9620
rect 32121 9618 32187 9621
rect 31036 9616 32187 9618
rect 31036 9560 32126 9616
rect 32182 9560 32187 9616
rect 31036 9558 32187 9560
rect 31036 9556 31042 9558
rect 32121 9555 32187 9558
rect 34513 9618 34579 9621
rect 35985 9618 36051 9621
rect 34513 9616 36051 9618
rect 34513 9560 34518 9616
rect 34574 9560 35990 9616
rect 36046 9560 36051 9616
rect 34513 9558 36051 9560
rect 34513 9555 34579 9558
rect 35985 9555 36051 9558
rect 22134 9482 22140 9484
rect 21038 9422 22140 9482
rect 16316 9420 16322 9422
rect 20897 9419 20963 9422
rect 22134 9420 22140 9422
rect 22204 9482 22210 9484
rect 28257 9482 28323 9485
rect 22204 9480 28323 9482
rect 22204 9424 28262 9480
rect 28318 9424 28323 9480
rect 22204 9422 28323 9424
rect 22204 9420 22210 9422
rect 28257 9419 28323 9422
rect 28901 9482 28967 9485
rect 37958 9482 37964 9484
rect 28901 9480 37964 9482
rect 28901 9424 28906 9480
rect 28962 9424 37964 9480
rect 28901 9422 37964 9424
rect 28901 9419 28967 9422
rect 37958 9420 37964 9422
rect 38028 9420 38034 9484
rect 24761 9346 24827 9349
rect 31569 9346 31635 9349
rect 24761 9344 31635 9346
rect 24761 9288 24766 9344
rect 24822 9288 31574 9344
rect 31630 9288 31635 9344
rect 24761 9286 31635 9288
rect 24761 9283 24827 9286
rect 31569 9283 31635 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 21173 9210 21239 9213
rect 26785 9210 26851 9213
rect 27245 9210 27311 9213
rect 27705 9212 27771 9213
rect 38009 9212 38075 9213
rect 21173 9208 27311 9210
rect 21173 9152 21178 9208
rect 21234 9152 26790 9208
rect 26846 9152 27250 9208
rect 27306 9152 27311 9208
rect 21173 9150 27311 9152
rect 21173 9147 21239 9150
rect 26785 9147 26851 9150
rect 27245 9147 27311 9150
rect 27654 9148 27660 9212
rect 27724 9210 27771 9212
rect 27724 9208 27816 9210
rect 27766 9152 27816 9208
rect 27724 9150 27816 9152
rect 27724 9148 27771 9150
rect 37958 9148 37964 9212
rect 38028 9210 38075 9212
rect 38028 9208 38120 9210
rect 38070 9152 38120 9208
rect 38028 9150 38120 9152
rect 38028 9148 38075 9150
rect 27705 9147 27771 9148
rect 38009 9147 38075 9148
rect 20897 9074 20963 9077
rect 21214 9074 21220 9076
rect 20897 9072 21220 9074
rect 20897 9016 20902 9072
rect 20958 9016 21220 9072
rect 20897 9014 21220 9016
rect 20897 9011 20963 9014
rect 21214 9012 21220 9014
rect 21284 9074 21290 9076
rect 25037 9074 25103 9077
rect 21284 9072 25103 9074
rect 21284 9016 25042 9072
rect 25098 9016 25103 9072
rect 21284 9014 25103 9016
rect 21284 9012 21290 9014
rect 25037 9011 25103 9014
rect 29729 9074 29795 9077
rect 29862 9074 29868 9076
rect 29729 9072 29868 9074
rect 29729 9016 29734 9072
rect 29790 9016 29868 9072
rect 29729 9014 29868 9016
rect 29729 9011 29795 9014
rect 29862 9012 29868 9014
rect 29932 9012 29938 9076
rect 31109 9074 31175 9077
rect 35341 9074 35407 9077
rect 31109 9072 35407 9074
rect 31109 9016 31114 9072
rect 31170 9016 35346 9072
rect 35402 9016 35407 9072
rect 31109 9014 35407 9016
rect 31109 9011 31175 9014
rect 35341 9011 35407 9014
rect 7005 8938 7071 8941
rect 8201 8938 8267 8941
rect 7005 8936 8267 8938
rect 7005 8880 7010 8936
rect 7066 8880 8206 8936
rect 8262 8880 8267 8936
rect 7005 8878 8267 8880
rect 7005 8875 7071 8878
rect 8201 8875 8267 8878
rect 11094 8876 11100 8940
rect 11164 8938 11170 8940
rect 11881 8938 11947 8941
rect 11164 8936 11947 8938
rect 11164 8880 11886 8936
rect 11942 8880 11947 8936
rect 11164 8878 11947 8880
rect 11164 8876 11170 8878
rect 11881 8875 11947 8878
rect 24209 8938 24275 8941
rect 34237 8938 34303 8941
rect 24209 8936 34303 8938
rect 24209 8880 24214 8936
rect 24270 8880 34242 8936
rect 34298 8880 34303 8936
rect 24209 8878 34303 8880
rect 24209 8875 24275 8878
rect 34237 8875 34303 8878
rect 24945 8804 25011 8805
rect 24894 8802 24900 8804
rect 24854 8742 24900 8802
rect 24964 8800 25011 8804
rect 25006 8744 25011 8800
rect 24894 8740 24900 8742
rect 24964 8740 25011 8744
rect 24945 8739 25011 8740
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 23289 8668 23355 8669
rect 23238 8604 23244 8668
rect 23308 8666 23355 8668
rect 24209 8666 24275 8669
rect 28809 8666 28875 8669
rect 23308 8664 23400 8666
rect 23350 8608 23400 8664
rect 23308 8606 23400 8608
rect 24209 8664 28875 8666
rect 24209 8608 24214 8664
rect 24270 8608 28814 8664
rect 28870 8608 28875 8664
rect 24209 8606 28875 8608
rect 23308 8604 23355 8606
rect 23289 8603 23355 8604
rect 24209 8603 24275 8606
rect 28809 8603 28875 8606
rect 29729 8666 29795 8669
rect 29729 8664 31770 8666
rect 29729 8608 29734 8664
rect 29790 8608 31770 8664
rect 29729 8606 31770 8608
rect 29729 8603 29795 8606
rect 15653 8530 15719 8533
rect 30373 8530 30439 8533
rect 15653 8528 30439 8530
rect 15653 8472 15658 8528
rect 15714 8472 30378 8528
rect 30434 8472 30439 8528
rect 15653 8470 30439 8472
rect 31710 8530 31770 8606
rect 37733 8530 37799 8533
rect 31710 8528 37799 8530
rect 31710 8472 37738 8528
rect 37794 8472 37799 8528
rect 31710 8470 37799 8472
rect 15653 8467 15719 8470
rect 30373 8467 30439 8470
rect 37733 8467 37799 8470
rect 7005 8394 7071 8397
rect 7925 8394 7991 8397
rect 7005 8392 7991 8394
rect 7005 8336 7010 8392
rect 7066 8336 7930 8392
rect 7986 8336 7991 8392
rect 7005 8334 7991 8336
rect 7005 8331 7071 8334
rect 7925 8331 7991 8334
rect 18822 8332 18828 8396
rect 18892 8394 18898 8396
rect 19425 8394 19491 8397
rect 18892 8392 19491 8394
rect 18892 8336 19430 8392
rect 19486 8336 19491 8392
rect 18892 8334 19491 8336
rect 18892 8332 18898 8334
rect 19425 8331 19491 8334
rect 20069 8394 20135 8397
rect 22185 8394 22251 8397
rect 20069 8392 22251 8394
rect 20069 8336 20074 8392
rect 20130 8336 22190 8392
rect 22246 8336 22251 8392
rect 20069 8334 22251 8336
rect 20069 8331 20135 8334
rect 22185 8331 22251 8334
rect 23841 8394 23907 8397
rect 27245 8394 27311 8397
rect 23841 8392 27311 8394
rect 23841 8336 23846 8392
rect 23902 8336 27250 8392
rect 27306 8336 27311 8392
rect 23841 8334 27311 8336
rect 23841 8331 23907 8334
rect 27245 8331 27311 8334
rect 28993 8394 29059 8397
rect 34329 8394 34395 8397
rect 28993 8392 34395 8394
rect 28993 8336 28998 8392
rect 29054 8336 34334 8392
rect 34390 8336 34395 8392
rect 28993 8334 34395 8336
rect 28993 8331 29059 8334
rect 34329 8331 34395 8334
rect 10542 8196 10548 8260
rect 10612 8258 10618 8260
rect 11605 8258 11671 8261
rect 10612 8256 11671 8258
rect 10612 8200 11610 8256
rect 11666 8200 11671 8256
rect 10612 8198 11671 8200
rect 10612 8196 10618 8198
rect 11605 8195 11671 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 15561 8122 15627 8125
rect 24669 8124 24735 8125
rect 16062 8122 16068 8124
rect 15561 8120 16068 8122
rect 15561 8064 15566 8120
rect 15622 8064 16068 8120
rect 15561 8062 16068 8064
rect 15561 8059 15627 8062
rect 16062 8060 16068 8062
rect 16132 8060 16138 8124
rect 24669 8122 24716 8124
rect 24624 8120 24716 8122
rect 24624 8064 24674 8120
rect 24624 8062 24716 8064
rect 24669 8060 24716 8062
rect 24780 8060 24786 8124
rect 24669 8059 24735 8060
rect 14089 7986 14155 7989
rect 33501 7988 33567 7989
rect 14222 7986 14228 7988
rect 14089 7984 14228 7986
rect 14089 7928 14094 7984
rect 14150 7928 14228 7984
rect 14089 7926 14228 7928
rect 14089 7923 14155 7926
rect 14222 7924 14228 7926
rect 14292 7924 14298 7988
rect 33501 7986 33548 7988
rect 33456 7984 33548 7986
rect 33456 7928 33506 7984
rect 33456 7926 33548 7928
rect 33501 7924 33548 7926
rect 33612 7924 33618 7988
rect 33501 7923 33567 7924
rect 24117 7850 24183 7853
rect 27153 7850 27219 7853
rect 24117 7848 27219 7850
rect 24117 7792 24122 7848
rect 24178 7792 27158 7848
rect 27214 7792 27219 7848
rect 24117 7790 27219 7792
rect 24117 7787 24183 7790
rect 27153 7787 27219 7790
rect 20437 7714 20503 7717
rect 23841 7714 23907 7717
rect 20437 7712 23907 7714
rect 20437 7656 20442 7712
rect 20498 7656 23846 7712
rect 23902 7656 23907 7712
rect 20437 7654 23907 7656
rect 20437 7651 20503 7654
rect 23841 7651 23907 7654
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 29545 7578 29611 7581
rect 29678 7578 29684 7580
rect 29545 7576 29684 7578
rect 29545 7520 29550 7576
rect 29606 7520 29684 7576
rect 29545 7518 29684 7520
rect 29545 7515 29611 7518
rect 29678 7516 29684 7518
rect 29748 7516 29754 7580
rect 12525 7442 12591 7445
rect 12750 7442 12756 7444
rect 12525 7440 12756 7442
rect 12525 7384 12530 7440
rect 12586 7384 12756 7440
rect 12525 7382 12756 7384
rect 12525 7379 12591 7382
rect 12750 7380 12756 7382
rect 12820 7380 12826 7444
rect 21081 7442 21147 7445
rect 29177 7442 29243 7445
rect 21081 7440 29243 7442
rect 21081 7384 21086 7440
rect 21142 7384 29182 7440
rect 29238 7384 29243 7440
rect 21081 7382 29243 7384
rect 21081 7379 21147 7382
rect 29177 7379 29243 7382
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 24209 7036 24275 7037
rect 24158 6972 24164 7036
rect 24228 7034 24275 7036
rect 24228 7032 24320 7034
rect 24270 6976 24320 7032
rect 24228 6974 24320 6976
rect 24228 6972 24275 6974
rect 24209 6971 24275 6972
rect 10910 6836 10916 6900
rect 10980 6898 10986 6900
rect 11513 6898 11579 6901
rect 10980 6896 11579 6898
rect 10980 6840 11518 6896
rect 11574 6840 11579 6896
rect 10980 6838 11579 6840
rect 10980 6836 10986 6838
rect 11513 6835 11579 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 16389 6492 16455 6493
rect 16389 6490 16436 6492
rect 16344 6488 16436 6490
rect 16344 6432 16394 6488
rect 16344 6430 16436 6432
rect 16389 6428 16436 6430
rect 16500 6428 16506 6492
rect 16389 6427 16455 6428
rect 29545 6354 29611 6357
rect 36118 6354 36124 6356
rect 29545 6352 36124 6354
rect 29545 6296 29550 6352
rect 29606 6296 36124 6352
rect 29545 6294 36124 6296
rect 29545 6291 29611 6294
rect 36118 6292 36124 6294
rect 36188 6292 36194 6356
rect 22369 6218 22435 6221
rect 33726 6218 33732 6220
rect 22369 6216 33732 6218
rect 22369 6160 22374 6216
rect 22430 6160 33732 6216
rect 22369 6158 33732 6160
rect 22369 6155 22435 6158
rect 33726 6156 33732 6158
rect 33796 6156 33802 6220
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19977 5946 20043 5949
rect 28717 5948 28783 5949
rect 20110 5946 20116 5948
rect 19977 5944 20116 5946
rect 19977 5888 19982 5944
rect 20038 5888 20116 5944
rect 19977 5886 20116 5888
rect 19977 5883 20043 5886
rect 20110 5884 20116 5886
rect 20180 5884 20186 5948
rect 28717 5946 28764 5948
rect 28672 5944 28764 5946
rect 28672 5888 28722 5944
rect 28672 5886 28764 5888
rect 28717 5884 28764 5886
rect 28828 5884 28834 5948
rect 28717 5883 28783 5884
rect 24485 5812 24551 5813
rect 24485 5810 24532 5812
rect 24440 5808 24532 5810
rect 24440 5752 24490 5808
rect 24440 5750 24532 5752
rect 24485 5748 24532 5750
rect 24596 5748 24602 5812
rect 24485 5747 24551 5748
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 19190 5340 19196 5404
rect 19260 5402 19266 5404
rect 21357 5402 21423 5405
rect 19260 5400 21423 5402
rect 19260 5344 21362 5400
rect 21418 5344 21423 5400
rect 19260 5342 21423 5344
rect 19260 5340 19266 5342
rect 21357 5339 21423 5342
rect 29177 5266 29243 5269
rect 29310 5266 29316 5268
rect 29177 5264 29316 5266
rect 29177 5208 29182 5264
rect 29238 5208 29316 5264
rect 29177 5206 29316 5208
rect 29177 5203 29243 5206
rect 29310 5204 29316 5206
rect 29380 5204 29386 5268
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 13905 4180 13971 4181
rect 13854 4116 13860 4180
rect 13924 4178 13971 4180
rect 13924 4176 14016 4178
rect 13966 4120 14016 4176
rect 13924 4118 14016 4120
rect 13924 4116 13971 4118
rect 13905 4115 13971 4116
rect 20478 3980 20484 4044
rect 20548 4042 20554 4044
rect 21357 4042 21423 4045
rect 21817 4042 21883 4045
rect 20548 4040 21883 4042
rect 20548 3984 21362 4040
rect 21418 3984 21822 4040
rect 21878 3984 21883 4040
rect 20548 3982 21883 3984
rect 20548 3980 20554 3982
rect 21357 3979 21423 3982
rect 21817 3979 21883 3982
rect 17718 3844 17724 3908
rect 17788 3906 17794 3908
rect 22829 3906 22895 3909
rect 17788 3904 22895 3906
rect 17788 3848 22834 3904
rect 22890 3848 22895 3904
rect 17788 3846 22895 3848
rect 17788 3844 17794 3846
rect 22829 3843 22895 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 40125 3498 40191 3501
rect 40957 3498 41757 3528
rect 40125 3496 41757 3498
rect 40125 3440 40130 3496
rect 40186 3440 41757 3496
rect 40125 3438 41757 3440
rect 40125 3435 40191 3438
rect 40957 3408 41757 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
<< via3 >>
rect 4876 41372 4940 41376
rect 4876 41316 4880 41372
rect 4880 41316 4936 41372
rect 4936 41316 4940 41372
rect 4876 41312 4940 41316
rect 4956 41372 5020 41376
rect 4956 41316 4960 41372
rect 4960 41316 5016 41372
rect 5016 41316 5020 41372
rect 4956 41312 5020 41316
rect 5036 41372 5100 41376
rect 5036 41316 5040 41372
rect 5040 41316 5096 41372
rect 5096 41316 5100 41372
rect 5036 41312 5100 41316
rect 5116 41372 5180 41376
rect 5116 41316 5120 41372
rect 5120 41316 5176 41372
rect 5176 41316 5180 41372
rect 5116 41312 5180 41316
rect 35596 41372 35660 41376
rect 35596 41316 35600 41372
rect 35600 41316 35656 41372
rect 35656 41316 35660 41372
rect 35596 41312 35660 41316
rect 35676 41372 35740 41376
rect 35676 41316 35680 41372
rect 35680 41316 35736 41372
rect 35736 41316 35740 41372
rect 35676 41312 35740 41316
rect 35756 41372 35820 41376
rect 35756 41316 35760 41372
rect 35760 41316 35816 41372
rect 35816 41316 35820 41372
rect 35756 41312 35820 41316
rect 35836 41372 35900 41376
rect 35836 41316 35840 41372
rect 35840 41316 35896 41372
rect 35896 41316 35900 41372
rect 35836 41312 35900 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 4876 40284 4940 40288
rect 4876 40228 4880 40284
rect 4880 40228 4936 40284
rect 4936 40228 4940 40284
rect 4876 40224 4940 40228
rect 4956 40284 5020 40288
rect 4956 40228 4960 40284
rect 4960 40228 5016 40284
rect 5016 40228 5020 40284
rect 4956 40224 5020 40228
rect 5036 40284 5100 40288
rect 5036 40228 5040 40284
rect 5040 40228 5096 40284
rect 5096 40228 5100 40284
rect 5036 40224 5100 40228
rect 5116 40284 5180 40288
rect 5116 40228 5120 40284
rect 5120 40228 5176 40284
rect 5176 40228 5180 40284
rect 5116 40224 5180 40228
rect 35596 40284 35660 40288
rect 35596 40228 35600 40284
rect 35600 40228 35656 40284
rect 35656 40228 35660 40284
rect 35596 40224 35660 40228
rect 35676 40284 35740 40288
rect 35676 40228 35680 40284
rect 35680 40228 35736 40284
rect 35736 40228 35740 40284
rect 35676 40224 35740 40228
rect 35756 40284 35820 40288
rect 35756 40228 35760 40284
rect 35760 40228 35816 40284
rect 35816 40228 35820 40284
rect 35756 40224 35820 40228
rect 35836 40284 35900 40288
rect 35836 40228 35840 40284
rect 35840 40228 35896 40284
rect 35896 40228 35900 40284
rect 35836 40224 35900 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 4876 39196 4940 39200
rect 4876 39140 4880 39196
rect 4880 39140 4936 39196
rect 4936 39140 4940 39196
rect 4876 39136 4940 39140
rect 4956 39196 5020 39200
rect 4956 39140 4960 39196
rect 4960 39140 5016 39196
rect 5016 39140 5020 39196
rect 4956 39136 5020 39140
rect 5036 39196 5100 39200
rect 5036 39140 5040 39196
rect 5040 39140 5096 39196
rect 5096 39140 5100 39196
rect 5036 39136 5100 39140
rect 5116 39196 5180 39200
rect 5116 39140 5120 39196
rect 5120 39140 5176 39196
rect 5176 39140 5180 39196
rect 5116 39136 5180 39140
rect 35596 39196 35660 39200
rect 35596 39140 35600 39196
rect 35600 39140 35656 39196
rect 35656 39140 35660 39196
rect 35596 39136 35660 39140
rect 35676 39196 35740 39200
rect 35676 39140 35680 39196
rect 35680 39140 35736 39196
rect 35736 39140 35740 39196
rect 35676 39136 35740 39140
rect 35756 39196 35820 39200
rect 35756 39140 35760 39196
rect 35760 39140 35816 39196
rect 35816 39140 35820 39196
rect 35756 39136 35820 39140
rect 35836 39196 35900 39200
rect 35836 39140 35840 39196
rect 35840 39140 35896 39196
rect 35896 39140 35900 39196
rect 35836 39136 35900 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 35596 38108 35660 38112
rect 35596 38052 35600 38108
rect 35600 38052 35656 38108
rect 35656 38052 35660 38108
rect 35596 38048 35660 38052
rect 35676 38108 35740 38112
rect 35676 38052 35680 38108
rect 35680 38052 35736 38108
rect 35736 38052 35740 38108
rect 35676 38048 35740 38052
rect 35756 38108 35820 38112
rect 35756 38052 35760 38108
rect 35760 38052 35816 38108
rect 35816 38052 35820 38108
rect 35756 38048 35820 38052
rect 35836 38108 35900 38112
rect 35836 38052 35840 38108
rect 35840 38052 35896 38108
rect 35896 38052 35900 38108
rect 35836 38048 35900 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 8156 35260 8220 35324
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 22508 32948 22572 33012
rect 30420 32948 30484 33012
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 9812 32540 9876 32604
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 18460 31996 18524 32060
rect 24532 32056 24596 32060
rect 24532 32000 24546 32056
rect 24546 32000 24596 32056
rect 24532 31996 24596 32000
rect 13676 31724 13740 31788
rect 27476 31724 27540 31788
rect 30604 31784 30668 31788
rect 30604 31728 30654 31784
rect 30654 31728 30668 31784
rect 30604 31724 30668 31728
rect 12020 31588 12084 31652
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 24900 31316 24964 31380
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 34652 30968 34716 30972
rect 34652 30912 34666 30968
rect 34666 30912 34716 30968
rect 34652 30908 34716 30912
rect 36124 30500 36188 30564
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 22140 30364 22204 30428
rect 29684 30364 29748 30428
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 30420 29880 30484 29884
rect 30420 29824 30470 29880
rect 30470 29824 30484 29880
rect 30420 29820 30484 29824
rect 35388 29820 35452 29884
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 35388 29276 35452 29340
rect 36124 29200 36188 29204
rect 36124 29144 36138 29200
rect 36138 29144 36188 29200
rect 36124 29140 36188 29144
rect 20116 29004 20180 29068
rect 34652 28928 34716 28932
rect 34652 28872 34702 28928
rect 34702 28872 34716 28928
rect 34652 28868 34716 28872
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 27108 28460 27172 28524
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 30604 28188 30668 28252
rect 5948 28112 6012 28116
rect 5948 28056 5998 28112
rect 5998 28056 6012 28112
rect 5948 28052 6012 28056
rect 9996 27916 10060 27980
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19932 27644 19996 27708
rect 32812 27296 32876 27300
rect 32812 27240 32826 27296
rect 32826 27240 32876 27296
rect 32812 27236 32876 27240
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 22324 26828 22388 26892
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 8340 26556 8404 26620
rect 8892 26616 8956 26620
rect 8892 26560 8942 26616
rect 8942 26560 8956 26616
rect 8892 26556 8956 26560
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 22140 26616 22204 26620
rect 22140 26560 22190 26616
rect 22190 26560 22204 26616
rect 22140 26556 22204 26560
rect 22508 26616 22572 26620
rect 22508 26560 22522 26616
rect 22522 26560 22572 26616
rect 22508 26556 22572 26560
rect 16436 26284 16500 26348
rect 16988 26344 17052 26348
rect 16988 26288 17002 26344
rect 17002 26288 17052 26344
rect 16988 26284 17052 26288
rect 19196 26284 19260 26348
rect 21772 26344 21836 26348
rect 21772 26288 21822 26344
rect 21822 26288 21836 26344
rect 21772 26284 21836 26288
rect 28028 26284 28092 26348
rect 28396 26284 28460 26348
rect 30788 26284 30852 26348
rect 38516 26284 38580 26348
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 13676 25936 13740 25940
rect 13676 25880 13690 25936
rect 13690 25880 13740 25936
rect 13676 25876 13740 25880
rect 29316 25800 29380 25804
rect 29316 25744 29366 25800
rect 29366 25744 29380 25800
rect 29316 25740 29380 25744
rect 32260 25604 32324 25668
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 17356 25468 17420 25532
rect 24900 25528 24964 25532
rect 24900 25472 24914 25528
rect 24914 25472 24964 25528
rect 24900 25468 24964 25472
rect 4660 25332 4724 25396
rect 16252 25332 16316 25396
rect 21220 25196 21284 25260
rect 33732 25256 33796 25260
rect 33732 25200 33746 25256
rect 33746 25200 33796 25256
rect 33732 25196 33796 25200
rect 35388 25196 35452 25260
rect 6132 25120 6196 25124
rect 6132 25064 6146 25120
rect 6146 25064 6196 25120
rect 6132 25060 6196 25064
rect 8340 25120 8404 25124
rect 8340 25064 8390 25120
rect 8390 25064 8404 25120
rect 8340 25060 8404 25064
rect 21404 25060 21468 25124
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 14228 24924 14292 24988
rect 24532 24924 24596 24988
rect 32996 24924 33060 24988
rect 22140 24788 22204 24852
rect 32444 24848 32508 24852
rect 32444 24792 32458 24848
rect 32458 24792 32508 24848
rect 32444 24788 32508 24792
rect 34652 24652 34716 24716
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 9996 24244 10060 24308
rect 28764 24244 28828 24308
rect 24900 24108 24964 24172
rect 26004 24108 26068 24172
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 5764 23564 5828 23628
rect 5948 23428 6012 23492
rect 23980 23428 24044 23492
rect 34468 23428 34532 23492
rect 37412 23428 37476 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 9812 23080 9876 23084
rect 9812 23024 9826 23080
rect 9826 23024 9876 23080
rect 9812 23020 9876 23024
rect 10732 23080 10796 23084
rect 10732 23024 10746 23080
rect 10746 23024 10796 23080
rect 10732 23020 10796 23024
rect 18644 23020 18708 23084
rect 13860 22944 13924 22948
rect 13860 22888 13874 22944
rect 13874 22888 13924 22944
rect 13860 22884 13924 22888
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 12020 22672 12084 22676
rect 12020 22616 12034 22672
rect 12034 22616 12084 22672
rect 12020 22612 12084 22616
rect 18828 22672 18892 22676
rect 18828 22616 18842 22672
rect 18842 22616 18892 22672
rect 18828 22612 18892 22616
rect 14044 22340 14108 22404
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 24164 22476 24228 22540
rect 36124 22476 36188 22540
rect 29868 22400 29932 22404
rect 29868 22344 29918 22400
rect 29918 22344 29932 22400
rect 29868 22340 29932 22344
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 22508 21992 22572 21996
rect 22508 21936 22522 21992
rect 22522 21936 22572 21992
rect 22508 21932 22572 21936
rect 21220 21796 21284 21860
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 28028 21584 28092 21588
rect 28028 21528 28042 21584
rect 28042 21528 28092 21584
rect 28028 21524 28092 21528
rect 28948 21584 29012 21588
rect 28948 21528 28998 21584
rect 28998 21528 29012 21584
rect 28948 21524 29012 21528
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 4660 20980 4724 21044
rect 8340 20980 8404 21044
rect 36308 20980 36372 21044
rect 16068 20708 16132 20772
rect 27476 20844 27540 20908
rect 34652 20844 34716 20908
rect 21956 20768 22020 20772
rect 21956 20712 22006 20768
rect 22006 20712 22020 20768
rect 21956 20708 22020 20712
rect 23244 20708 23308 20772
rect 24348 20708 24412 20772
rect 30420 20708 30484 20772
rect 34468 20708 34532 20772
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 21404 20572 21468 20636
rect 20484 20300 20548 20364
rect 28580 20300 28644 20364
rect 17724 20164 17788 20228
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 6132 19952 6196 19956
rect 6132 19896 6182 19952
rect 6182 19896 6196 19952
rect 6132 19892 6196 19896
rect 21588 19892 21652 19956
rect 38516 19892 38580 19956
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 35388 19348 35452 19412
rect 32812 19212 32876 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 30236 18804 30300 18868
rect 28764 18728 28828 18732
rect 28764 18672 28778 18728
rect 28778 18672 28828 18728
rect 28764 18668 28828 18672
rect 29684 18668 29748 18732
rect 34284 18668 34348 18732
rect 28396 18592 28460 18596
rect 28396 18536 28410 18592
rect 28410 18536 28460 18592
rect 28396 18532 28460 18536
rect 28764 18532 28828 18596
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 18460 18260 18524 18324
rect 34468 18320 34532 18324
rect 34468 18264 34482 18320
rect 34482 18264 34532 18320
rect 34468 18260 34532 18264
rect 36308 18124 36372 18188
rect 37964 17988 38028 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 8892 17852 8956 17916
rect 30420 17852 30484 17916
rect 17356 17716 17420 17780
rect 28028 17716 28092 17780
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 24532 17308 24596 17372
rect 10732 17036 10796 17100
rect 11100 17036 11164 17100
rect 14044 17036 14108 17100
rect 20116 17036 20180 17100
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 32996 17036 33060 17100
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 10548 16688 10612 16692
rect 10548 16632 10562 16688
rect 10562 16632 10612 16688
rect 10548 16628 10612 16632
rect 11836 16628 11900 16692
rect 31892 16628 31956 16692
rect 30604 16356 30668 16420
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 12756 16008 12820 16012
rect 12756 15952 12806 16008
rect 12806 15952 12820 16008
rect 12756 15948 12820 15952
rect 10916 15872 10980 15876
rect 10916 15816 10930 15872
rect 10930 15816 10980 15872
rect 10916 15812 10980 15816
rect 22324 15812 22388 15876
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 22140 15600 22204 15604
rect 22140 15544 22154 15600
rect 22154 15544 22204 15600
rect 22140 15540 22204 15544
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 18644 15132 18708 15196
rect 20116 15132 20180 15196
rect 25820 15132 25884 15196
rect 37412 15268 37476 15332
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 25636 14996 25700 15060
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19932 14588 19996 14652
rect 21772 14588 21836 14652
rect 30972 14316 31036 14380
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 23980 14104 24044 14108
rect 23980 14048 23994 14104
rect 23994 14048 24044 14104
rect 23980 14044 24044 14048
rect 25820 14044 25884 14108
rect 27108 14104 27172 14108
rect 27108 14048 27122 14104
rect 27122 14048 27172 14104
rect 27108 14044 27172 14048
rect 27660 13908 27724 13972
rect 25452 13772 25516 13836
rect 28580 13772 28644 13836
rect 28948 13636 29012 13700
rect 32444 13636 32508 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 31892 13560 31956 13564
rect 31892 13504 31906 13560
rect 31906 13504 31956 13560
rect 31892 13500 31956 13504
rect 34652 13152 34716 13156
rect 34652 13096 34702 13152
rect 34702 13096 34716 13152
rect 34652 13092 34716 13096
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 34284 12684 34348 12748
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 30236 12412 30300 12476
rect 24348 12276 24412 12340
rect 32996 12276 33060 12340
rect 11836 12004 11900 12068
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 19380 11868 19444 11932
rect 21956 11928 22020 11932
rect 21956 11872 22006 11928
rect 22006 11872 22020 11928
rect 21956 11868 22020 11872
rect 22508 11732 22572 11796
rect 25452 11732 25516 11796
rect 32260 11732 32324 11796
rect 33548 11792 33612 11796
rect 33548 11736 33598 11792
rect 33598 11736 33612 11792
rect 33548 11732 33612 11736
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 24716 11188 24780 11252
rect 26004 11188 26068 11252
rect 30788 11188 30852 11252
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 25820 10780 25884 10844
rect 21588 10644 21652 10708
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 5764 10296 5828 10300
rect 5764 10240 5778 10296
rect 5778 10240 5828 10296
rect 5764 10236 5828 10240
rect 16988 10236 17052 10300
rect 30604 10100 30668 10164
rect 25636 10024 25700 10028
rect 25636 9968 25650 10024
rect 25650 9968 25700 10024
rect 25636 9964 25700 9968
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 19380 9692 19444 9756
rect 34468 9692 34532 9756
rect 16252 9420 16316 9484
rect 30972 9556 31036 9620
rect 22140 9420 22204 9484
rect 37964 9420 38028 9484
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 27660 9208 27724 9212
rect 27660 9152 27710 9208
rect 27710 9152 27724 9208
rect 27660 9148 27724 9152
rect 37964 9208 38028 9212
rect 37964 9152 38014 9208
rect 38014 9152 38028 9208
rect 37964 9148 38028 9152
rect 21220 9012 21284 9076
rect 29868 9012 29932 9076
rect 11100 8876 11164 8940
rect 24900 8800 24964 8804
rect 24900 8744 24950 8800
rect 24950 8744 24964 8800
rect 24900 8740 24964 8744
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 23244 8664 23308 8668
rect 23244 8608 23294 8664
rect 23294 8608 23308 8664
rect 23244 8604 23308 8608
rect 18828 8332 18892 8396
rect 10548 8196 10612 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 16068 8060 16132 8124
rect 24716 8120 24780 8124
rect 24716 8064 24730 8120
rect 24730 8064 24780 8120
rect 24716 8060 24780 8064
rect 14228 7924 14292 7988
rect 33548 7984 33612 7988
rect 33548 7928 33562 7984
rect 33562 7928 33612 7984
rect 33548 7924 33612 7928
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 29684 7516 29748 7580
rect 12756 7380 12820 7444
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 24164 7032 24228 7036
rect 24164 6976 24214 7032
rect 24214 6976 24228 7032
rect 24164 6972 24228 6976
rect 10916 6836 10980 6900
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 16436 6488 16500 6492
rect 16436 6432 16450 6488
rect 16450 6432 16500 6488
rect 16436 6428 16500 6432
rect 36124 6292 36188 6356
rect 33732 6156 33796 6220
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 20116 5884 20180 5948
rect 28764 5944 28828 5948
rect 28764 5888 28778 5944
rect 28778 5888 28828 5944
rect 28764 5884 28828 5888
rect 24532 5808 24596 5812
rect 24532 5752 24546 5808
rect 24546 5752 24596 5808
rect 24532 5748 24596 5752
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 19196 5340 19260 5404
rect 29316 5204 29380 5268
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 13860 4176 13924 4180
rect 13860 4120 13910 4176
rect 13910 4120 13924 4176
rect 13860 4116 13924 4120
rect 20484 3980 20548 4044
rect 17724 3844 17788 3908
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
<< metal4 >>
rect 4208 40832 4528 41392
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4868 41376 5188 41392
rect 4868 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5188 41376
rect 4868 40288 5188 41312
rect 4868 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5188 40288
rect 4868 39200 5188 40224
rect 4868 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5188 39200
rect 4868 38112 5188 39136
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 35936 5188 36960
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 34928 40832 35248 41392
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 8155 35324 8221 35325
rect 8155 35260 8156 35324
rect 8220 35260 8221 35324
rect 8155 35259 8221 35260
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 8158 29610 8218 35259
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 22507 33012 22573 33013
rect 22507 32948 22508 33012
rect 22572 32948 22573 33012
rect 22507 32947 22573 32948
rect 30419 33012 30485 33013
rect 30419 32948 30420 33012
rect 30484 32948 30485 33012
rect 30419 32947 30485 32948
rect 9811 32604 9877 32605
rect 9811 32540 9812 32604
rect 9876 32540 9877 32604
rect 9811 32539 9877 32540
rect 8158 29550 8402 29610
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 5947 28116 6013 28117
rect 5947 28052 5948 28116
rect 6012 28052 6013 28116
rect 5947 28051 6013 28052
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4659 25396 4725 25397
rect 4659 25332 4660 25396
rect 4724 25332 4725 25396
rect 4659 25331 4725 25332
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4662 21045 4722 25331
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 5763 23628 5829 23629
rect 5763 23564 5764 23628
rect 5828 23564 5829 23628
rect 5763 23563 5829 23564
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4659 21044 4725 21045
rect 4659 20980 4660 21044
rect 4724 20980 4725 21044
rect 4659 20979 4725 20980
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 5766 10301 5826 23563
rect 5950 23493 6010 28051
rect 8342 26621 8402 29550
rect 8339 26620 8405 26621
rect 8339 26556 8340 26620
rect 8404 26556 8405 26620
rect 8339 26555 8405 26556
rect 8891 26620 8957 26621
rect 8891 26556 8892 26620
rect 8956 26556 8957 26620
rect 8891 26555 8957 26556
rect 6131 25124 6197 25125
rect 6131 25060 6132 25124
rect 6196 25060 6197 25124
rect 6131 25059 6197 25060
rect 8339 25124 8405 25125
rect 8339 25060 8340 25124
rect 8404 25060 8405 25124
rect 8339 25059 8405 25060
rect 5947 23492 6013 23493
rect 5947 23428 5948 23492
rect 6012 23428 6013 23492
rect 5947 23427 6013 23428
rect 6134 19957 6194 25059
rect 8342 21045 8402 25059
rect 8339 21044 8405 21045
rect 8339 20980 8340 21044
rect 8404 20980 8405 21044
rect 8339 20979 8405 20980
rect 6131 19956 6197 19957
rect 6131 19892 6132 19956
rect 6196 19892 6197 19956
rect 6131 19891 6197 19892
rect 8894 17917 8954 26555
rect 9814 23085 9874 32539
rect 18459 32060 18525 32061
rect 18459 31996 18460 32060
rect 18524 31996 18525 32060
rect 18459 31995 18525 31996
rect 13675 31788 13741 31789
rect 13675 31724 13676 31788
rect 13740 31724 13741 31788
rect 13675 31723 13741 31724
rect 12019 31652 12085 31653
rect 12019 31588 12020 31652
rect 12084 31588 12085 31652
rect 12019 31587 12085 31588
rect 9995 27980 10061 27981
rect 9995 27916 9996 27980
rect 10060 27916 10061 27980
rect 9995 27915 10061 27916
rect 9998 24309 10058 27915
rect 9995 24308 10061 24309
rect 9995 24244 9996 24308
rect 10060 24244 10061 24308
rect 9995 24243 10061 24244
rect 9811 23084 9877 23085
rect 9811 23020 9812 23084
rect 9876 23020 9877 23084
rect 9811 23019 9877 23020
rect 10731 23084 10797 23085
rect 10731 23020 10732 23084
rect 10796 23020 10797 23084
rect 10731 23019 10797 23020
rect 8891 17916 8957 17917
rect 8891 17852 8892 17916
rect 8956 17852 8957 17916
rect 8891 17851 8957 17852
rect 10734 17101 10794 23019
rect 12022 22677 12082 31587
rect 13678 25941 13738 31723
rect 16435 26348 16501 26349
rect 16435 26284 16436 26348
rect 16500 26284 16501 26348
rect 16435 26283 16501 26284
rect 16987 26348 17053 26349
rect 16987 26284 16988 26348
rect 17052 26284 17053 26348
rect 16987 26283 17053 26284
rect 13675 25940 13741 25941
rect 13675 25876 13676 25940
rect 13740 25876 13741 25940
rect 13675 25875 13741 25876
rect 16251 25396 16317 25397
rect 16251 25332 16252 25396
rect 16316 25332 16317 25396
rect 16251 25331 16317 25332
rect 14227 24988 14293 24989
rect 14227 24924 14228 24988
rect 14292 24924 14293 24988
rect 14227 24923 14293 24924
rect 13859 22948 13925 22949
rect 13859 22884 13860 22948
rect 13924 22884 13925 22948
rect 13859 22883 13925 22884
rect 12019 22676 12085 22677
rect 12019 22612 12020 22676
rect 12084 22612 12085 22676
rect 12019 22611 12085 22612
rect 10731 17100 10797 17101
rect 10731 17036 10732 17100
rect 10796 17036 10797 17100
rect 10731 17035 10797 17036
rect 11099 17100 11165 17101
rect 11099 17036 11100 17100
rect 11164 17036 11165 17100
rect 11099 17035 11165 17036
rect 10547 16692 10613 16693
rect 10547 16628 10548 16692
rect 10612 16628 10613 16692
rect 10547 16627 10613 16628
rect 5763 10300 5829 10301
rect 5763 10236 5764 10300
rect 5828 10236 5829 10300
rect 5763 10235 5829 10236
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 10550 8261 10610 16627
rect 10915 15876 10981 15877
rect 10915 15812 10916 15876
rect 10980 15812 10981 15876
rect 10915 15811 10981 15812
rect 10547 8260 10613 8261
rect 10547 8196 10548 8260
rect 10612 8196 10613 8260
rect 10547 8195 10613 8196
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 10918 6901 10978 15811
rect 11102 8941 11162 17035
rect 11835 16692 11901 16693
rect 11835 16628 11836 16692
rect 11900 16628 11901 16692
rect 11835 16627 11901 16628
rect 11838 12069 11898 16627
rect 12755 16012 12821 16013
rect 12755 15948 12756 16012
rect 12820 15948 12821 16012
rect 12755 15947 12821 15948
rect 11835 12068 11901 12069
rect 11835 12004 11836 12068
rect 11900 12004 11901 12068
rect 11835 12003 11901 12004
rect 11099 8940 11165 8941
rect 11099 8876 11100 8940
rect 11164 8876 11165 8940
rect 11099 8875 11165 8876
rect 12758 7445 12818 15947
rect 12755 7444 12821 7445
rect 12755 7380 12756 7444
rect 12820 7380 12821 7444
rect 12755 7379 12821 7380
rect 10915 6900 10981 6901
rect 10915 6836 10916 6900
rect 10980 6836 10981 6900
rect 10915 6835 10981 6836
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 13862 4181 13922 22883
rect 14043 22404 14109 22405
rect 14043 22340 14044 22404
rect 14108 22340 14109 22404
rect 14043 22339 14109 22340
rect 14046 17101 14106 22339
rect 14043 17100 14109 17101
rect 14043 17036 14044 17100
rect 14108 17036 14109 17100
rect 14043 17035 14109 17036
rect 14230 7989 14290 24923
rect 16067 20772 16133 20773
rect 16067 20708 16068 20772
rect 16132 20708 16133 20772
rect 16067 20707 16133 20708
rect 16070 8125 16130 20707
rect 16254 9485 16314 25331
rect 16251 9484 16317 9485
rect 16251 9420 16252 9484
rect 16316 9420 16317 9484
rect 16251 9419 16317 9420
rect 16067 8124 16133 8125
rect 16067 8060 16068 8124
rect 16132 8060 16133 8124
rect 16067 8059 16133 8060
rect 14227 7988 14293 7989
rect 14227 7924 14228 7988
rect 14292 7924 14293 7988
rect 14227 7923 14293 7924
rect 16438 6493 16498 26283
rect 16990 10301 17050 26283
rect 17355 25532 17421 25533
rect 17355 25468 17356 25532
rect 17420 25468 17421 25532
rect 17355 25467 17421 25468
rect 17358 17781 17418 25467
rect 17723 20228 17789 20229
rect 17723 20164 17724 20228
rect 17788 20164 17789 20228
rect 17723 20163 17789 20164
rect 17355 17780 17421 17781
rect 17355 17716 17356 17780
rect 17420 17716 17421 17780
rect 17355 17715 17421 17716
rect 16987 10300 17053 10301
rect 16987 10236 16988 10300
rect 17052 10236 17053 10300
rect 16987 10235 17053 10236
rect 16435 6492 16501 6493
rect 16435 6428 16436 6492
rect 16500 6428 16501 6492
rect 16435 6427 16501 6428
rect 13859 4180 13925 4181
rect 13859 4116 13860 4180
rect 13924 4116 13925 4180
rect 13859 4115 13925 4116
rect 17726 3909 17786 20163
rect 18462 18325 18522 31995
rect 22139 30428 22205 30429
rect 22139 30364 22140 30428
rect 22204 30364 22205 30428
rect 22139 30363 22205 30364
rect 20115 29068 20181 29069
rect 20115 29004 20116 29068
rect 20180 29004 20181 29068
rect 20115 29003 20181 29004
rect 19931 27708 19997 27709
rect 19931 27644 19932 27708
rect 19996 27644 19997 27708
rect 19931 27643 19997 27644
rect 19195 26348 19261 26349
rect 19195 26284 19196 26348
rect 19260 26284 19261 26348
rect 19195 26283 19261 26284
rect 18643 23084 18709 23085
rect 18643 23020 18644 23084
rect 18708 23020 18709 23084
rect 18643 23019 18709 23020
rect 18459 18324 18525 18325
rect 18459 18260 18460 18324
rect 18524 18260 18525 18324
rect 18459 18259 18525 18260
rect 18646 15197 18706 23019
rect 18827 22676 18893 22677
rect 18827 22612 18828 22676
rect 18892 22612 18893 22676
rect 18827 22611 18893 22612
rect 18643 15196 18709 15197
rect 18643 15132 18644 15196
rect 18708 15132 18709 15196
rect 18643 15131 18709 15132
rect 18830 8397 18890 22611
rect 18827 8396 18893 8397
rect 18827 8332 18828 8396
rect 18892 8332 18893 8396
rect 18827 8331 18893 8332
rect 19198 5405 19258 26283
rect 19934 14653 19994 27643
rect 20118 17101 20178 29003
rect 22142 26621 22202 30363
rect 22323 26892 22389 26893
rect 22323 26828 22324 26892
rect 22388 26828 22389 26892
rect 22323 26827 22389 26828
rect 22139 26620 22205 26621
rect 22139 26556 22140 26620
rect 22204 26556 22205 26620
rect 22139 26555 22205 26556
rect 21771 26348 21837 26349
rect 21771 26284 21772 26348
rect 21836 26284 21837 26348
rect 21771 26283 21837 26284
rect 21219 25260 21285 25261
rect 21219 25196 21220 25260
rect 21284 25196 21285 25260
rect 21219 25195 21285 25196
rect 21222 21861 21282 25195
rect 21403 25124 21469 25125
rect 21403 25060 21404 25124
rect 21468 25060 21469 25124
rect 21403 25059 21469 25060
rect 21219 21860 21285 21861
rect 21219 21796 21220 21860
rect 21284 21796 21285 21860
rect 21219 21795 21285 21796
rect 20483 20364 20549 20365
rect 20483 20300 20484 20364
rect 20548 20300 20549 20364
rect 20483 20299 20549 20300
rect 20115 17100 20181 17101
rect 20115 17036 20116 17100
rect 20180 17036 20181 17100
rect 20115 17035 20181 17036
rect 20115 15196 20181 15197
rect 20115 15132 20116 15196
rect 20180 15132 20181 15196
rect 20115 15131 20181 15132
rect 19931 14652 19997 14653
rect 19931 14588 19932 14652
rect 19996 14588 19997 14652
rect 19931 14587 19997 14588
rect 19379 11932 19445 11933
rect 19379 11868 19380 11932
rect 19444 11868 19445 11932
rect 19379 11867 19445 11868
rect 19382 9757 19442 11867
rect 19379 9756 19445 9757
rect 19379 9692 19380 9756
rect 19444 9692 19445 9756
rect 19379 9691 19445 9692
rect 20118 5949 20178 15131
rect 20115 5948 20181 5949
rect 20115 5884 20116 5948
rect 20180 5884 20181 5948
rect 20115 5883 20181 5884
rect 19195 5404 19261 5405
rect 19195 5340 19196 5404
rect 19260 5340 19261 5404
rect 19195 5339 19261 5340
rect 20486 4045 20546 20299
rect 21222 9077 21282 21795
rect 21406 20637 21466 25059
rect 21403 20636 21469 20637
rect 21403 20572 21404 20636
rect 21468 20572 21469 20636
rect 21403 20571 21469 20572
rect 21587 19956 21653 19957
rect 21587 19892 21588 19956
rect 21652 19892 21653 19956
rect 21587 19891 21653 19892
rect 21590 10709 21650 19891
rect 21774 14653 21834 26283
rect 22139 24852 22205 24853
rect 22139 24788 22140 24852
rect 22204 24788 22205 24852
rect 22139 24787 22205 24788
rect 21955 20772 22021 20773
rect 21955 20708 21956 20772
rect 22020 20708 22021 20772
rect 21955 20707 22021 20708
rect 21771 14652 21837 14653
rect 21771 14588 21772 14652
rect 21836 14588 21837 14652
rect 21771 14587 21837 14588
rect 21958 11933 22018 20707
rect 22142 15605 22202 24787
rect 22326 15877 22386 26827
rect 22510 26621 22570 32947
rect 24531 32060 24597 32061
rect 24531 31996 24532 32060
rect 24596 31996 24597 32060
rect 24531 31995 24597 31996
rect 22507 26620 22573 26621
rect 22507 26556 22508 26620
rect 22572 26556 22573 26620
rect 22507 26555 22573 26556
rect 24534 24989 24594 31995
rect 27475 31788 27541 31789
rect 27475 31724 27476 31788
rect 27540 31724 27541 31788
rect 27475 31723 27541 31724
rect 24899 31380 24965 31381
rect 24899 31316 24900 31380
rect 24964 31316 24965 31380
rect 24899 31315 24965 31316
rect 24902 25533 24962 31315
rect 27107 28524 27173 28525
rect 27107 28460 27108 28524
rect 27172 28460 27173 28524
rect 27107 28459 27173 28460
rect 24899 25532 24965 25533
rect 24899 25468 24900 25532
rect 24964 25468 24965 25532
rect 24899 25467 24965 25468
rect 24531 24988 24597 24989
rect 24531 24924 24532 24988
rect 24596 24924 24597 24988
rect 24531 24923 24597 24924
rect 24899 24172 24965 24173
rect 24899 24108 24900 24172
rect 24964 24108 24965 24172
rect 24899 24107 24965 24108
rect 26003 24172 26069 24173
rect 26003 24108 26004 24172
rect 26068 24108 26069 24172
rect 26003 24107 26069 24108
rect 23979 23492 24045 23493
rect 23979 23428 23980 23492
rect 24044 23428 24045 23492
rect 23979 23427 24045 23428
rect 22507 21996 22573 21997
rect 22507 21932 22508 21996
rect 22572 21932 22573 21996
rect 22507 21931 22573 21932
rect 22323 15876 22389 15877
rect 22323 15812 22324 15876
rect 22388 15812 22389 15876
rect 22323 15811 22389 15812
rect 22139 15604 22205 15605
rect 22139 15540 22140 15604
rect 22204 15540 22205 15604
rect 22139 15539 22205 15540
rect 21955 11932 22021 11933
rect 21955 11868 21956 11932
rect 22020 11868 22021 11932
rect 21955 11867 22021 11868
rect 21587 10708 21653 10709
rect 21587 10644 21588 10708
rect 21652 10644 21653 10708
rect 21587 10643 21653 10644
rect 22142 9485 22202 15539
rect 22510 11797 22570 21931
rect 23243 20772 23309 20773
rect 23243 20708 23244 20772
rect 23308 20708 23309 20772
rect 23243 20707 23309 20708
rect 22507 11796 22573 11797
rect 22507 11732 22508 11796
rect 22572 11732 22573 11796
rect 22507 11731 22573 11732
rect 22139 9484 22205 9485
rect 22139 9420 22140 9484
rect 22204 9420 22205 9484
rect 22139 9419 22205 9420
rect 21219 9076 21285 9077
rect 21219 9012 21220 9076
rect 21284 9012 21285 9076
rect 21219 9011 21285 9012
rect 23246 8669 23306 20707
rect 23982 14109 24042 23427
rect 24163 22540 24229 22541
rect 24163 22476 24164 22540
rect 24228 22476 24229 22540
rect 24163 22475 24229 22476
rect 23979 14108 24045 14109
rect 23979 14044 23980 14108
rect 24044 14044 24045 14108
rect 23979 14043 24045 14044
rect 23243 8668 23309 8669
rect 23243 8604 23244 8668
rect 23308 8604 23309 8668
rect 23243 8603 23309 8604
rect 24166 7037 24226 22475
rect 24347 20772 24413 20773
rect 24347 20708 24348 20772
rect 24412 20708 24413 20772
rect 24347 20707 24413 20708
rect 24350 12341 24410 20707
rect 24531 17372 24597 17373
rect 24531 17308 24532 17372
rect 24596 17308 24597 17372
rect 24531 17307 24597 17308
rect 24347 12340 24413 12341
rect 24347 12276 24348 12340
rect 24412 12276 24413 12340
rect 24347 12275 24413 12276
rect 24163 7036 24229 7037
rect 24163 6972 24164 7036
rect 24228 6972 24229 7036
rect 24163 6971 24229 6972
rect 24534 5813 24594 17307
rect 24715 11252 24781 11253
rect 24715 11188 24716 11252
rect 24780 11188 24781 11252
rect 24715 11187 24781 11188
rect 24718 8125 24778 11187
rect 24902 8805 24962 24107
rect 25819 15196 25885 15197
rect 25819 15132 25820 15196
rect 25884 15132 25885 15196
rect 25819 15131 25885 15132
rect 25635 15060 25701 15061
rect 25635 14996 25636 15060
rect 25700 14996 25701 15060
rect 25635 14995 25701 14996
rect 25451 13836 25517 13837
rect 25451 13772 25452 13836
rect 25516 13772 25517 13836
rect 25451 13771 25517 13772
rect 25454 11797 25514 13771
rect 25451 11796 25517 11797
rect 25451 11732 25452 11796
rect 25516 11732 25517 11796
rect 25451 11731 25517 11732
rect 25638 10029 25698 14995
rect 25822 14109 25882 15131
rect 25819 14108 25885 14109
rect 25819 14044 25820 14108
rect 25884 14044 25885 14108
rect 25819 14043 25885 14044
rect 25822 10845 25882 14043
rect 26006 11253 26066 24107
rect 27110 14109 27170 28459
rect 27478 20909 27538 31723
rect 29683 30428 29749 30429
rect 29683 30364 29684 30428
rect 29748 30364 29749 30428
rect 29683 30363 29749 30364
rect 28027 26348 28093 26349
rect 28027 26284 28028 26348
rect 28092 26284 28093 26348
rect 28027 26283 28093 26284
rect 28395 26348 28461 26349
rect 28395 26284 28396 26348
rect 28460 26284 28461 26348
rect 28395 26283 28461 26284
rect 28030 21589 28090 26283
rect 28027 21588 28093 21589
rect 28027 21524 28028 21588
rect 28092 21524 28093 21588
rect 28027 21523 28093 21524
rect 27475 20908 27541 20909
rect 27475 20844 27476 20908
rect 27540 20844 27541 20908
rect 27475 20843 27541 20844
rect 28030 17781 28090 21523
rect 28398 18597 28458 26283
rect 29315 25804 29381 25805
rect 29315 25740 29316 25804
rect 29380 25740 29381 25804
rect 29315 25739 29381 25740
rect 28763 24308 28829 24309
rect 28763 24244 28764 24308
rect 28828 24244 28829 24308
rect 28763 24243 28829 24244
rect 28579 20364 28645 20365
rect 28579 20300 28580 20364
rect 28644 20300 28645 20364
rect 28579 20299 28645 20300
rect 28395 18596 28461 18597
rect 28395 18532 28396 18596
rect 28460 18532 28461 18596
rect 28395 18531 28461 18532
rect 28027 17780 28093 17781
rect 28027 17716 28028 17780
rect 28092 17716 28093 17780
rect 28027 17715 28093 17716
rect 27107 14108 27173 14109
rect 27107 14044 27108 14108
rect 27172 14044 27173 14108
rect 27107 14043 27173 14044
rect 27659 13972 27725 13973
rect 27659 13908 27660 13972
rect 27724 13908 27725 13972
rect 27659 13907 27725 13908
rect 26003 11252 26069 11253
rect 26003 11188 26004 11252
rect 26068 11188 26069 11252
rect 26003 11187 26069 11188
rect 25819 10844 25885 10845
rect 25819 10780 25820 10844
rect 25884 10780 25885 10844
rect 25819 10779 25885 10780
rect 25635 10028 25701 10029
rect 25635 9964 25636 10028
rect 25700 9964 25701 10028
rect 25635 9963 25701 9964
rect 27662 9213 27722 13907
rect 28582 13837 28642 20299
rect 28766 18733 28826 24243
rect 28947 21588 29013 21589
rect 28947 21524 28948 21588
rect 29012 21524 29013 21588
rect 28947 21523 29013 21524
rect 28763 18732 28829 18733
rect 28763 18668 28764 18732
rect 28828 18668 28829 18732
rect 28763 18667 28829 18668
rect 28763 18596 28829 18597
rect 28763 18532 28764 18596
rect 28828 18532 28829 18596
rect 28763 18531 28829 18532
rect 28579 13836 28645 13837
rect 28579 13772 28580 13836
rect 28644 13772 28645 13836
rect 28579 13771 28645 13772
rect 27659 9212 27725 9213
rect 27659 9148 27660 9212
rect 27724 9148 27725 9212
rect 27659 9147 27725 9148
rect 24899 8804 24965 8805
rect 24899 8740 24900 8804
rect 24964 8740 24965 8804
rect 24899 8739 24965 8740
rect 24715 8124 24781 8125
rect 24715 8060 24716 8124
rect 24780 8060 24781 8124
rect 24715 8059 24781 8060
rect 28766 5949 28826 18531
rect 28950 13701 29010 21523
rect 28947 13700 29013 13701
rect 28947 13636 28948 13700
rect 29012 13636 29013 13700
rect 28947 13635 29013 13636
rect 28763 5948 28829 5949
rect 28763 5884 28764 5948
rect 28828 5884 28829 5948
rect 28763 5883 28829 5884
rect 24531 5812 24597 5813
rect 24531 5748 24532 5812
rect 24596 5748 24597 5812
rect 24531 5747 24597 5748
rect 29318 5269 29378 25739
rect 29686 18733 29746 30363
rect 30422 29885 30482 32947
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 30603 31788 30669 31789
rect 30603 31724 30604 31788
rect 30668 31724 30669 31788
rect 30603 31723 30669 31724
rect 30419 29884 30485 29885
rect 30419 29820 30420 29884
rect 30484 29820 30485 29884
rect 30419 29819 30485 29820
rect 30606 28253 30666 31723
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34651 30972 34717 30973
rect 34651 30908 34652 30972
rect 34716 30908 34717 30972
rect 34651 30907 34717 30908
rect 34654 28933 34714 30907
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34651 28932 34717 28933
rect 34651 28868 34652 28932
rect 34716 28868 34717 28932
rect 34651 28867 34717 28868
rect 34928 28864 35248 29888
rect 35588 41376 35908 41392
rect 35588 41312 35596 41376
rect 35660 41312 35676 41376
rect 35740 41312 35756 41376
rect 35820 41312 35836 41376
rect 35900 41312 35908 41376
rect 35588 40288 35908 41312
rect 35588 40224 35596 40288
rect 35660 40224 35676 40288
rect 35740 40224 35756 40288
rect 35820 40224 35836 40288
rect 35900 40224 35908 40288
rect 35588 39200 35908 40224
rect 35588 39136 35596 39200
rect 35660 39136 35676 39200
rect 35740 39136 35756 39200
rect 35820 39136 35836 39200
rect 35900 39136 35908 39200
rect 35588 38112 35908 39136
rect 35588 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35908 38112
rect 35588 37024 35908 38048
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 35936 35908 36960
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 36123 30564 36189 30565
rect 36123 30500 36124 30564
rect 36188 30500 36189 30564
rect 36123 30499 36189 30500
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35387 29884 35453 29885
rect 35387 29820 35388 29884
rect 35452 29820 35453 29884
rect 35387 29819 35453 29820
rect 35390 29341 35450 29819
rect 35588 29408 35908 30432
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35387 29340 35453 29341
rect 35387 29276 35388 29340
rect 35452 29276 35453 29340
rect 35387 29275 35453 29276
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 30603 28252 30669 28253
rect 30603 28188 30604 28252
rect 30668 28188 30669 28252
rect 30603 28187 30669 28188
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 32811 27300 32877 27301
rect 32811 27236 32812 27300
rect 32876 27236 32877 27300
rect 32811 27235 32877 27236
rect 30787 26348 30853 26349
rect 30787 26284 30788 26348
rect 30852 26284 30853 26348
rect 30787 26283 30853 26284
rect 29867 22404 29933 22405
rect 29867 22340 29868 22404
rect 29932 22340 29933 22404
rect 29867 22339 29933 22340
rect 29683 18732 29749 18733
rect 29683 18668 29684 18732
rect 29748 18668 29749 18732
rect 29683 18667 29749 18668
rect 29686 7581 29746 18667
rect 29870 9077 29930 22339
rect 30419 20772 30485 20773
rect 30419 20708 30420 20772
rect 30484 20708 30485 20772
rect 30419 20707 30485 20708
rect 30235 18868 30301 18869
rect 30235 18804 30236 18868
rect 30300 18804 30301 18868
rect 30235 18803 30301 18804
rect 30238 12477 30298 18803
rect 30422 17917 30482 20707
rect 30419 17916 30485 17917
rect 30419 17852 30420 17916
rect 30484 17852 30485 17916
rect 30419 17851 30485 17852
rect 30603 16420 30669 16421
rect 30603 16356 30604 16420
rect 30668 16356 30669 16420
rect 30603 16355 30669 16356
rect 30235 12476 30301 12477
rect 30235 12412 30236 12476
rect 30300 12412 30301 12476
rect 30235 12411 30301 12412
rect 30606 10165 30666 16355
rect 30790 11253 30850 26283
rect 32259 25668 32325 25669
rect 32259 25604 32260 25668
rect 32324 25604 32325 25668
rect 32259 25603 32325 25604
rect 31891 16692 31957 16693
rect 31891 16628 31892 16692
rect 31956 16628 31957 16692
rect 31891 16627 31957 16628
rect 30971 14380 31037 14381
rect 30971 14316 30972 14380
rect 31036 14316 31037 14380
rect 30971 14315 31037 14316
rect 30787 11252 30853 11253
rect 30787 11188 30788 11252
rect 30852 11188 30853 11252
rect 30787 11187 30853 11188
rect 30603 10164 30669 10165
rect 30603 10100 30604 10164
rect 30668 10100 30669 10164
rect 30603 10099 30669 10100
rect 30974 9621 31034 14315
rect 31894 13565 31954 16627
rect 31891 13564 31957 13565
rect 31891 13500 31892 13564
rect 31956 13500 31957 13564
rect 31891 13499 31957 13500
rect 32262 11797 32322 25603
rect 32443 24852 32509 24853
rect 32443 24788 32444 24852
rect 32508 24788 32509 24852
rect 32443 24787 32509 24788
rect 32446 13701 32506 24787
rect 32814 19277 32874 27235
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 33731 25260 33797 25261
rect 33731 25196 33732 25260
rect 33796 25196 33797 25260
rect 33731 25195 33797 25196
rect 32995 24988 33061 24989
rect 32995 24924 32996 24988
rect 33060 24924 33061 24988
rect 32995 24923 33061 24924
rect 32811 19276 32877 19277
rect 32811 19212 32812 19276
rect 32876 19212 32877 19276
rect 32811 19211 32877 19212
rect 32998 17101 33058 24923
rect 32995 17100 33061 17101
rect 32995 17036 32996 17100
rect 33060 17036 33061 17100
rect 32995 17035 33061 17036
rect 32443 13700 32509 13701
rect 32443 13636 32444 13700
rect 32508 13636 32509 13700
rect 32443 13635 32509 13636
rect 32998 12341 33058 17035
rect 32995 12340 33061 12341
rect 32995 12276 32996 12340
rect 33060 12276 33061 12340
rect 32995 12275 33061 12276
rect 32259 11796 32325 11797
rect 32259 11732 32260 11796
rect 32324 11732 32325 11796
rect 32259 11731 32325 11732
rect 33547 11796 33613 11797
rect 33547 11732 33548 11796
rect 33612 11732 33613 11796
rect 33547 11731 33613 11732
rect 30971 9620 31037 9621
rect 30971 9556 30972 9620
rect 31036 9556 31037 9620
rect 30971 9555 31037 9556
rect 29867 9076 29933 9077
rect 29867 9012 29868 9076
rect 29932 9012 29933 9076
rect 29867 9011 29933 9012
rect 33550 7989 33610 11731
rect 33547 7988 33613 7989
rect 33547 7924 33548 7988
rect 33612 7924 33613 7988
rect 33547 7923 33613 7924
rect 29683 7580 29749 7581
rect 29683 7516 29684 7580
rect 29748 7516 29749 7580
rect 29683 7515 29749 7516
rect 33734 6221 33794 25195
rect 34651 24716 34717 24717
rect 34651 24652 34652 24716
rect 34716 24652 34717 24716
rect 34651 24651 34717 24652
rect 34467 23492 34533 23493
rect 34467 23428 34468 23492
rect 34532 23428 34533 23492
rect 34467 23427 34533 23428
rect 34470 20773 34530 23427
rect 34654 20909 34714 24651
rect 34928 24512 35248 25536
rect 35588 28320 35908 29344
rect 36126 29205 36186 30499
rect 36123 29204 36189 29205
rect 36123 29140 36124 29204
rect 36188 29140 36189 29204
rect 36123 29139 36189 29140
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35588 27232 35908 28256
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 38515 26348 38581 26349
rect 38515 26284 38516 26348
rect 38580 26284 38581 26348
rect 38515 26283 38581 26284
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35387 25260 35453 25261
rect 35387 25196 35388 25260
rect 35452 25196 35453 25260
rect 35387 25195 35453 25196
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34651 20908 34717 20909
rect 34651 20844 34652 20908
rect 34716 20844 34717 20908
rect 34651 20843 34717 20844
rect 34467 20772 34533 20773
rect 34467 20708 34468 20772
rect 34532 20708 34533 20772
rect 34467 20707 34533 20708
rect 34283 18732 34349 18733
rect 34283 18668 34284 18732
rect 34348 18668 34349 18732
rect 34283 18667 34349 18668
rect 34286 12749 34346 18667
rect 34467 18324 34533 18325
rect 34467 18260 34468 18324
rect 34532 18260 34533 18324
rect 34467 18259 34533 18260
rect 34283 12748 34349 12749
rect 34283 12684 34284 12748
rect 34348 12684 34349 12748
rect 34283 12683 34349 12684
rect 34470 9757 34530 18259
rect 34654 13157 34714 20843
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 35390 19413 35450 25195
rect 35588 25056 35908 26080
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35588 22880 35908 23904
rect 37411 23492 37477 23493
rect 37411 23428 37412 23492
rect 37476 23428 37477 23492
rect 37411 23427 37477 23428
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 36123 22540 36189 22541
rect 36123 22476 36124 22540
rect 36188 22476 36189 22540
rect 36123 22475 36189 22476
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35387 19412 35453 19413
rect 35387 19348 35388 19412
rect 35452 19348 35453 19412
rect 35387 19347 35453 19348
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34651 13156 34717 13157
rect 34651 13092 34652 13156
rect 34716 13092 34717 13156
rect 34651 13091 34717 13092
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34467 9756 34533 9757
rect 34467 9692 34468 9756
rect 34532 9692 34533 9756
rect 34467 9691 34533 9692
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 33731 6220 33797 6221
rect 33731 6156 33732 6220
rect 33796 6156 33797 6220
rect 33731 6155 33797 6156
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 29315 5268 29381 5269
rect 29315 5204 29316 5268
rect 29380 5204 29381 5268
rect 29315 5203 29381 5204
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 20483 4044 20549 4045
rect 20483 3980 20484 4044
rect 20548 3980 20549 4044
rect 20483 3979 20549 3980
rect 17723 3908 17789 3909
rect 17723 3844 17724 3908
rect 17788 3844 17789 3908
rect 17723 3843 17789 3844
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 18528 35908 19552
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35588 14176 35908 15200
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 5472 35908 6496
rect 36126 6357 36186 22475
rect 36307 21044 36373 21045
rect 36307 20980 36308 21044
rect 36372 20980 36373 21044
rect 36307 20979 36373 20980
rect 36310 18189 36370 20979
rect 36307 18188 36373 18189
rect 36307 18124 36308 18188
rect 36372 18124 36373 18188
rect 36307 18123 36373 18124
rect 37414 15333 37474 23427
rect 38518 19957 38578 26283
rect 38515 19956 38581 19957
rect 38515 19892 38516 19956
rect 38580 19892 38581 19956
rect 38515 19891 38581 19892
rect 37963 18052 38029 18053
rect 37963 17988 37964 18052
rect 38028 17988 38029 18052
rect 37963 17987 38029 17988
rect 37411 15332 37477 15333
rect 37411 15268 37412 15332
rect 37476 15268 37477 15332
rect 37411 15267 37477 15268
rect 37966 9485 38026 17987
rect 37963 9484 38029 9485
rect 37963 9420 37964 9484
rect 38028 9420 38029 9484
rect 37963 9419 38029 9420
rect 37966 9213 38026 9419
rect 37963 9212 38029 9213
rect 37963 9148 37964 9212
rect 38028 9148 38029 9212
rect 37963 9147 38029 9148
rect 36123 6356 36189 6357
rect 36123 6292 36124 6356
rect 36188 6292 36189 6356
rect 36123 6291 36189 6292
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
use sky130_fd_sc_hd__inv_2  _1336_
timestamp 18001
transform 1 0 27600 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1337_
timestamp 18001
transform -1 0 28796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1338_
timestamp 18001
transform -1 0 28520 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1339_
timestamp 18001
transform 1 0 24932 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1340_
timestamp 18001
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1341_
timestamp 18001
transform -1 0 18032 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1342_
timestamp 18001
transform -1 0 20148 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1343_
timestamp 18001
transform 1 0 31280 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1344_
timestamp 18001
transform 1 0 20516 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1345_
timestamp 18001
transform -1 0 19504 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1346_
timestamp 18001
transform 1 0 15640 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1347_
timestamp 18001
transform 1 0 34224 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_1  _1348_
timestamp 18001
transform -1 0 32200 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1349_
timestamp 18001
transform 1 0 31188 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1350_
timestamp 18001
transform -1 0 24564 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1351_
timestamp 18001
transform 1 0 21344 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1352_
timestamp 18001
transform 1 0 33304 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_4  _1353_
timestamp 18001
transform 1 0 29808 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__and2b_2  _1354_
timestamp 18001
transform -1 0 29440 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_2  _1355_
timestamp 18001
transform 1 0 32384 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__or4bb_2  _1356_
timestamp 18001
transform 1 0 29624 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _1357_
timestamp 18001
transform -1 0 30360 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1358_
timestamp 18001
transform -1 0 37444 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor4b_1  _1359_
timestamp 18001
transform 1 0 26220 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_2  _1360_
timestamp 18001
transform -1 0 31280 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1361_
timestamp 18001
transform -1 0 30820 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1362_
timestamp 18001
transform -1 0 24748 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1363_
timestamp 18001
transform -1 0 24288 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1364_
timestamp 18001
transform -1 0 34960 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1365_
timestamp 18001
transform -1 0 29716 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1366_
timestamp 18001
transform -1 0 37536 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1367_
timestamp 18001
transform -1 0 29440 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1368_
timestamp 18001
transform -1 0 30544 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1369_
timestamp 18001
transform -1 0 28152 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1370_
timestamp 18001
transform -1 0 34316 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_4  _1371_
timestamp 18001
transform -1 0 30728 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__and4b_4  _1372_
timestamp 18001
transform 1 0 31280 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__and2_1  _1373_
timestamp 18001
transform -1 0 30728 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1374_
timestamp 18001
transform -1 0 27324 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1375_
timestamp 18001
transform -1 0 26036 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1376_
timestamp 18001
transform -1 0 18952 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1377_
timestamp 18001
transform 1 0 25392 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1378_
timestamp 18001
transform 1 0 22540 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _1379_
timestamp 18001
transform 1 0 24012 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_2  _1380_
timestamp 18001
transform 1 0 32752 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__or4bb_2  _1381_
timestamp 18001
transform -1 0 27876 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _1382_
timestamp 18001
transform 1 0 25852 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1383_
timestamp 18001
transform 1 0 29532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1384_
timestamp 18001
transform 1 0 26404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor4b_2  _1385_
timestamp 18001
transform -1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__or4b_4  _1386_
timestamp 18001
transform -1 0 27416 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _1387_
timestamp 18001
transform -1 0 25300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1388_
timestamp 18001
transform -1 0 26312 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1389_
timestamp 18001
transform 1 0 25852 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1390_
timestamp 18001
transform -1 0 26772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _1391_
timestamp 18001
transform -1 0 30820 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_4  _1392_
timestamp 18001
transform -1 0 30452 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_4  _1393_
timestamp 18001
transform 1 0 34684 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__or4bb_4  _1394_
timestamp 18001
transform -1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _1395_
timestamp 18001
transform -1 0 25852 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1396_
timestamp 18001
transform -1 0 25668 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1397_
timestamp 18001
transform 1 0 24196 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1398_
timestamp 18001
transform -1 0 33856 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1399_
timestamp 18001
transform -1 0 30912 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_2  _1400_
timestamp 18001
transform -1 0 33028 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or4_2  _1401_
timestamp 18001
transform -1 0 27324 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1402_
timestamp 18001
transform 1 0 26956 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor4b_2  _1403_
timestamp 18001
transform -1 0 35972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__or4b_2  _1404_
timestamp 18001
transform 1 0 28060 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1405_
timestamp 18001
transform 1 0 28980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1406_
timestamp 18001
transform 1 0 26220 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _1407_
timestamp 18001
transform 1 0 24288 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a311o_1  _1408_
timestamp 18001
transform 1 0 26956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_2  _1409_
timestamp 18001
transform 1 0 23552 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1410_
timestamp 18001
transform -1 0 22632 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1411_
timestamp 18001
transform 1 0 22632 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1412_
timestamp 18001
transform -1 0 22724 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1413_
timestamp 18001
transform 1 0 23184 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1414_
timestamp 18001
transform 1 0 22816 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1415_
timestamp 18001
transform -1 0 17204 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_2  _1416_
timestamp 18001
transform -1 0 34592 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _1417_
timestamp 18001
transform -1 0 36800 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__o31a_1  _1418_
timestamp 18001
transform 1 0 28704 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_2  _1419_
timestamp 18001
transform 1 0 33304 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1420_
timestamp 18001
transform 1 0 37444 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _1421_
timestamp 18001
transform -1 0 28704 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1422_
timestamp 18001
transform -1 0 26404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _1423_
timestamp 18001
transform -1 0 29072 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1424_
timestamp 18001
transform 1 0 25300 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1425_
timestamp 18001
transform -1 0 26404 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1426_
timestamp 18001
transform 1 0 24840 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1427_
timestamp 18001
transform -1 0 25668 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1428_
timestamp 18001
transform -1 0 25944 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1429_
timestamp 18001
transform 1 0 24380 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1430_
timestamp 18001
transform 1 0 24380 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a2111oi_4  _1431_
timestamp 18001
transform 1 0 24748 0 -1 8704
box -38 -48 2062 592
use sky130_fd_sc_hd__and4_2  _1432_
timestamp 18001
transform -1 0 25300 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1433_
timestamp 18001
transform 1 0 25760 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1434_
timestamp 18001
transform -1 0 19320 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _1435_
timestamp 18001
transform -1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1436_
timestamp 18001
transform -1 0 27508 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1437_
timestamp 18001
transform -1 0 30360 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1438_
timestamp 18001
transform -1 0 34960 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1439_
timestamp 18001
transform -1 0 27416 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1440_
timestamp 18001
transform 1 0 24472 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1441_
timestamp 18001
transform -1 0 28244 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1442_
timestamp 18001
transform -1 0 32844 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1443_
timestamp 18001
transform -1 0 30084 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1444_
timestamp 18001
transform 1 0 21804 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1445_
timestamp 18001
transform -1 0 20792 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1446_
timestamp 18001
transform -1 0 22724 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1447_
timestamp 18001
transform -1 0 22448 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1448_
timestamp 18001
transform 1 0 22080 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1449_
timestamp 18001
transform -1 0 30820 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1450_
timestamp 18001
transform -1 0 20240 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1451_
timestamp 18001
transform 1 0 24932 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1452_
timestamp 18001
transform 1 0 25116 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1453_
timestamp 18001
transform -1 0 23460 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_2  _1454_
timestamp 18001
transform -1 0 31648 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1455_
timestamp 18001
transform 1 0 31096 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1456_
timestamp 18001
transform -1 0 24472 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1457_
timestamp 18001
transform -1 0 29348 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1458_
timestamp 18001
transform -1 0 25392 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1459_
timestamp 18001
transform -1 0 25944 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1460_
timestamp 18001
transform 1 0 25116 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1461_
timestamp 18001
transform -1 0 25116 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1462_
timestamp 18001
transform 1 0 25484 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1463_
timestamp 18001
transform 1 0 26220 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1464_
timestamp 18001
transform -1 0 30084 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1465_
timestamp 18001
transform -1 0 31464 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1466_
timestamp 18001
transform 1 0 30268 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1467_
timestamp 18001
transform 1 0 29900 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1468_
timestamp 18001
transform -1 0 31096 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1469_
timestamp 18001
transform 1 0 28060 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1470_
timestamp 18001
transform -1 0 31648 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1471_
timestamp 18001
transform 1 0 28336 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1472_
timestamp 18001
transform 1 0 28336 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1473_
timestamp 18001
transform 1 0 20608 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _1474_
timestamp 18001
transform 1 0 21804 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1475_
timestamp 18001
transform 1 0 30452 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1476_
timestamp 18001
transform 1 0 30084 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1477_
timestamp 18001
transform -1 0 31096 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1478_
timestamp 18001
transform 1 0 26312 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1479_
timestamp 18001
transform -1 0 30820 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1480_
timestamp 18001
transform 1 0 30084 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1481_
timestamp 18001
transform -1 0 31372 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1482_
timestamp 18001
transform -1 0 34224 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1483_
timestamp 18001
transform 1 0 28704 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1484_
timestamp 18001
transform 1 0 28520 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1485_
timestamp 18001
transform -1 0 30544 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _1486_
timestamp 18001
transform -1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1487_
timestamp 18001
transform 1 0 24472 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1488_
timestamp 18001
transform -1 0 25944 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1489_
timestamp 18001
transform -1 0 30636 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1490_
timestamp 18001
transform 1 0 30452 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1491_
timestamp 18001
transform -1 0 30728 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1492_
timestamp 18001
transform 1 0 28980 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1493_
timestamp 18001
transform -1 0 28428 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1494_
timestamp 18001
transform 1 0 28428 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1495_
timestamp 18001
transform -1 0 30176 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1496_
timestamp 18001
transform -1 0 27140 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1497_
timestamp 18001
transform 1 0 23920 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1498_
timestamp 18001
transform 1 0 28520 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1499_
timestamp 18001
transform -1 0 28520 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1500_
timestamp 18001
transform 1 0 27876 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1501_
timestamp 18001
transform 1 0 26220 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1502_
timestamp 18001
transform -1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _1503_
timestamp 18001
transform 1 0 29348 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1504_
timestamp 18001
transform 1 0 30176 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1505_
timestamp 18001
transform 1 0 27508 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1506_
timestamp 18001
transform -1 0 28796 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1507_
timestamp 18001
transform 1 0 24564 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1508_
timestamp 18001
transform -1 0 18860 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _1509_
timestamp 18001
transform -1 0 21988 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_2  _1510_
timestamp 18001
transform -1 0 28704 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1511_
timestamp 18001
transform -1 0 29072 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a32oi_4  _1512_
timestamp 18001
transform 1 0 27140 0 1 29376
box -38 -48 2062 592
use sky130_fd_sc_hd__a32o_1  _1513_
timestamp 18001
transform 1 0 28060 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_2  _1514_
timestamp 18001
transform -1 0 28336 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1515_
timestamp 18001
transform 1 0 25484 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1516_
timestamp 18001
transform 1 0 29532 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_4  _1517_
timestamp 18001
transform -1 0 27140 0 1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_1  _1518_
timestamp 18001
transform 1 0 26404 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_2  _1519_
timestamp 18001
transform -1 0 28060 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__a211oi_4  _1520_
timestamp 18001
transform 1 0 29532 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__a22o_1  _1521_
timestamp 18001
transform 1 0 24472 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1522_
timestamp 18001
transform -1 0 27600 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1523_
timestamp 18001
transform 1 0 28980 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1524_
timestamp 18001
transform 1 0 39468 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1525_
timestamp 18001
transform 1 0 29808 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a311o_1  _1526_
timestamp 18001
transform 1 0 29532 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1527_
timestamp 18001
transform 1 0 28796 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1528_
timestamp 18001
transform 1 0 29532 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1529_
timestamp 18001
transform -1 0 25760 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1530_
timestamp 18001
transform 1 0 26220 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1531_
timestamp 18001
transform 1 0 21252 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _1532_
timestamp 18001
transform -1 0 22908 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _1533_
timestamp 18001
transform 1 0 32108 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _1534_
timestamp 18001
transform 1 0 39192 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1535_
timestamp 18001
transform 1 0 34224 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1536_
timestamp 18001
transform -1 0 30728 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1537_
timestamp 18001
transform 1 0 34408 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1538_
timestamp 18001
transform -1 0 34316 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1539_
timestamp 18001
transform 1 0 37904 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1540_
timestamp 18001
transform 1 0 37260 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1541_
timestamp 18001
transform 1 0 38180 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1542_
timestamp 18001
transform -1 0 38456 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1543_
timestamp 18001
transform -1 0 37812 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1544_
timestamp 18001
transform -1 0 39100 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1545_
timestamp 18001
transform -1 0 33028 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1546_
timestamp 18001
transform -1 0 38824 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _1547_
timestamp 18001
transform -1 0 36892 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1548_
timestamp 18001
transform 1 0 33396 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1549_
timestamp 18001
transform 1 0 35696 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1550_
timestamp 18001
transform 1 0 36892 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1551_
timestamp 18001
transform 1 0 37260 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1552_
timestamp 18001
transform 1 0 36064 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1553_
timestamp 18001
transform -1 0 35236 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1554_
timestamp 18001
transform 1 0 35604 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1555_
timestamp 18001
transform -1 0 36708 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1556_
timestamp 18001
transform 1 0 36708 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1557_
timestamp 18001
transform -1 0 34960 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1558_
timestamp 18001
transform 1 0 37260 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1559_
timestamp 18001
transform 1 0 37352 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1560_
timestamp 18001
transform 1 0 38180 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1561_
timestamp 18001
transform 1 0 32660 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1562_
timestamp 18001
transform 1 0 36248 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1563_
timestamp 18001
transform -1 0 31832 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1564_
timestamp 18001
transform 1 0 30820 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1565_
timestamp 18001
transform -1 0 31464 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1566_
timestamp 18001
transform -1 0 31556 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1567_
timestamp 18001
transform -1 0 31004 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1568_
timestamp 18001
transform -1 0 35696 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1569_
timestamp 18001
transform -1 0 29808 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1570_
timestamp 18001
transform -1 0 29808 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1571_
timestamp 18001
transform 1 0 28520 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1572_
timestamp 18001
transform 1 0 38272 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _1573_
timestamp 18001
transform -1 0 33764 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1574_
timestamp 18001
transform 1 0 32476 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1575_
timestamp 18001
transform -1 0 32016 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1576_
timestamp 18001
transform 1 0 32660 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1577_
timestamp 18001
transform 1 0 32108 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1578_
timestamp 18001
transform 1 0 32844 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1579_
timestamp 18001
transform 1 0 32108 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1580_
timestamp 18001
transform 1 0 32200 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1581_
timestamp 18001
transform -1 0 36064 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1582_
timestamp 18001
transform -1 0 34500 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1583_
timestamp 18001
transform -1 0 32936 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1584_
timestamp 18001
transform 1 0 32568 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1585_
timestamp 18001
transform 1 0 33948 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1586_
timestamp 18001
transform 1 0 29532 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1587_
timestamp 18001
transform -1 0 35144 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1588_
timestamp 18001
transform 1 0 35512 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1589_
timestamp 18001
transform -1 0 31924 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1590_
timestamp 18001
transform 1 0 34224 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1591_
timestamp 18001
transform 1 0 33580 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1592_
timestamp 18001
transform 1 0 33212 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1593_
timestamp 18001
transform 1 0 30912 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1594_
timestamp 18001
transform -1 0 36984 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _1595_
timestamp 18001
transform -1 0 36524 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1596_
timestamp 18001
transform 1 0 30820 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1597_
timestamp 18001
transform 1 0 31648 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1598_
timestamp 18001
transform 1 0 31924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1599_
timestamp 18001
transform 1 0 30176 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1600_
timestamp 18001
transform -1 0 33672 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _1601_
timestamp 18001
transform -1 0 35420 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1602_
timestamp 18001
transform 1 0 31280 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_2  _1603_
timestamp 18001
transform -1 0 38456 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1604_
timestamp 18001
transform -1 0 36800 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1605_
timestamp 18001
transform 1 0 33948 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1606_
timestamp 18001
transform 1 0 34684 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_4  _1607_
timestamp 18001
transform -1 0 31832 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1608_
timestamp 18001
transform 1 0 32108 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1609_
timestamp 18001
transform -1 0 33948 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _1610_
timestamp 18001
transform 1 0 32844 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1611_
timestamp 18001
transform -1 0 33396 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1612_
timestamp 18001
transform -1 0 31648 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1613_
timestamp 18001
transform -1 0 31372 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1614_
timestamp 18001
transform 1 0 31188 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1615_
timestamp 18001
transform 1 0 37260 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1616_
timestamp 18001
transform -1 0 37444 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1617_
timestamp 18001
transform 1 0 31556 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1618_
timestamp 18001
transform 1 0 37260 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1619_
timestamp 18001
transform 1 0 36064 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1620_
timestamp 18001
transform 1 0 37996 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1621_
timestamp 18001
transform 1 0 31372 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1622_
timestamp 18001
transform 1 0 33488 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1623_
timestamp 18001
transform -1 0 32844 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1624_
timestamp 18001
transform -1 0 32568 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1625_
timestamp 18001
transform 1 0 31096 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1626_
timestamp 18001
transform 1 0 32752 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1627_
timestamp 18001
transform -1 0 31280 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _1628_
timestamp 18001
transform -1 0 39100 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1629_
timestamp 18001
transform -1 0 39376 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1630_
timestamp 18001
transform -1 0 36064 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _1631_
timestamp 18001
transform 1 0 35328 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1632_
timestamp 18001
transform -1 0 35696 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1633_
timestamp 18001
transform -1 0 34684 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _1634_
timestamp 18001
transform -1 0 35512 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1635_
timestamp 18001
transform -1 0 34592 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1636_
timestamp 18001
transform -1 0 35328 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1637_
timestamp 18001
transform -1 0 34132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1638_
timestamp 18001
transform -1 0 36524 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1639_
timestamp 18001
transform 1 0 36524 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1640_
timestamp 18001
transform -1 0 38548 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1641_
timestamp 18001
transform 1 0 37996 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1642_
timestamp 18001
transform -1 0 33948 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1643_
timestamp 18001
transform -1 0 35420 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1644_
timestamp 18001
transform 1 0 34776 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1645_
timestamp 18001
transform 1 0 38364 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1646_
timestamp 18001
transform -1 0 31648 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1647_
timestamp 18001
transform 1 0 31004 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1648_
timestamp 18001
transform 1 0 31096 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1649_
timestamp 18001
transform 1 0 32108 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1650_
timestamp 18001
transform -1 0 31924 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1651_
timestamp 18001
transform 1 0 32108 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1652_
timestamp 18001
transform 1 0 32936 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1653_
timestamp 18001
transform 1 0 31648 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1654_
timestamp 18001
transform 1 0 32568 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1655_
timestamp 18001
transform 1 0 33304 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1656_
timestamp 18001
transform 1 0 34224 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1657_
timestamp 18001
transform 1 0 35236 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1658_
timestamp 18001
transform 1 0 34132 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1659_
timestamp 18001
transform 1 0 35788 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1660_
timestamp 18001
transform -1 0 34408 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1661_
timestamp 18001
transform 1 0 37260 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1662_
timestamp 18001
transform -1 0 35328 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1663_
timestamp 18001
transform -1 0 31924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1664_
timestamp 18001
transform 1 0 30820 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1665_
timestamp 18001
transform 1 0 31464 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1666_
timestamp 18001
transform 1 0 32844 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1667_
timestamp 18001
transform 1 0 32108 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1668_
timestamp 18001
transform 1 0 36708 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1669_
timestamp 18001
transform 1 0 36524 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1670_
timestamp 18001
transform -1 0 36984 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1671_
timestamp 18001
transform 1 0 36984 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1672_
timestamp 18001
transform 1 0 38272 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1673_
timestamp 18001
transform -1 0 35236 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1674_
timestamp 18001
transform -1 0 36524 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1675_
timestamp 18001
transform 1 0 36156 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1676_
timestamp 18001
transform 1 0 38088 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1677_
timestamp 18001
transform -1 0 35144 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1678_
timestamp 18001
transform 1 0 33856 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1679_
timestamp 18001
transform -1 0 34868 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1680_
timestamp 18001
transform 1 0 35052 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1681_
timestamp 18001
transform 1 0 35696 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1682_
timestamp 18001
transform 1 0 34500 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1683_
timestamp 18001
transform 1 0 36064 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1684_
timestamp 18001
transform -1 0 31740 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1685_
timestamp 18001
transform -1 0 36156 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1686_
timestamp 18001
transform 1 0 38364 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1687_
timestamp 18001
transform -1 0 35788 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1688_
timestamp 18001
transform 1 0 36432 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1689_
timestamp 18001
transform 1 0 31740 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1690_
timestamp 18001
transform 1 0 32752 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1691_
timestamp 18001
transform 1 0 38088 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1692_
timestamp 18001
transform 1 0 38640 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1693_
timestamp 18001
transform 1 0 38824 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1694_
timestamp 18001
transform 1 0 32108 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1695_
timestamp 18001
transform 1 0 35604 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1696_
timestamp 18001
transform 1 0 38824 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1697_
timestamp 18001
transform -1 0 32844 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1698_
timestamp 18001
transform -1 0 33580 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1699_
timestamp 18001
transform -1 0 39192 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1700_
timestamp 18001
transform 1 0 32476 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1701_
timestamp 18001
transform 1 0 36616 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1702_
timestamp 18001
transform 1 0 36800 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1703_
timestamp 18001
transform -1 0 39008 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1704_
timestamp 18001
transform 1 0 39100 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1705_
timestamp 18001
transform -1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1706_
timestamp 18001
transform 1 0 36708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1707_
timestamp 18001
transform -1 0 34500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1708_
timestamp 18001
transform 1 0 36432 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1709_
timestamp 18001
transform 1 0 37444 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1710_
timestamp 18001
transform 1 0 38824 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1711_
timestamp 18001
transform 1 0 36064 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1712_
timestamp 18001
transform 1 0 38272 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1713_
timestamp 18001
transform 1 0 38640 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1714_
timestamp 18001
transform 1 0 37996 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1715_
timestamp 18001
transform -1 0 39100 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1716_
timestamp 18001
transform 1 0 38824 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1717_
timestamp 18001
transform 1 0 34960 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1718_
timestamp 18001
transform -1 0 38732 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1719_
timestamp 18001
transform 1 0 32384 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1720_
timestamp 18001
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1721_
timestamp 18001
transform 1 0 37904 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1722_
timestamp 18001
transform 1 0 38732 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1723_
timestamp 18001
transform -1 0 38732 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1724_
timestamp 18001
transform -1 0 38824 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1725_
timestamp 18001
transform 1 0 36524 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1726_
timestamp 18001
transform 1 0 37904 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1727_
timestamp 18001
transform 1 0 35420 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1728_
timestamp 18001
transform 1 0 33028 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1729_
timestamp 18001
transform 1 0 36064 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1730_
timestamp 18001
transform -1 0 37812 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1731_
timestamp 18001
transform 1 0 36248 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1732_
timestamp 18001
transform 1 0 37260 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1733_
timestamp 18001
transform 1 0 32568 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1734_
timestamp 18001
transform 1 0 34684 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1735_
timestamp 18001
transform 1 0 36708 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1736_
timestamp 18001
transform 1 0 25300 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1737_
timestamp 18001
transform -1 0 19044 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _1738_
timestamp 18001
transform -1 0 19780 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1739_
timestamp 18001
transform -1 0 18400 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1740_
timestamp 18001
transform 1 0 22632 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_2  _1741_
timestamp 18001
transform 1 0 21804 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1742_
timestamp 18001
transform 1 0 22080 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1743_
timestamp 18001
transform 1 0 19872 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _1744_
timestamp 18001
transform 1 0 16652 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1745_
timestamp 18001
transform -1 0 25392 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1746_
timestamp 18001
transform -1 0 24012 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1747_
timestamp 18001
transform -1 0 24104 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1748_
timestamp 18001
transform -1 0 23644 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1749_
timestamp 18001
transform 1 0 22908 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1750_
timestamp 18001
transform 1 0 21896 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _1751_
timestamp 18001
transform -1 0 21160 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1752_
timestamp 18001
transform -1 0 19412 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1753_
timestamp 18001
transform -1 0 21344 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1754_
timestamp 18001
transform -1 0 24288 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1755_
timestamp 18001
transform 1 0 20148 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1756_
timestamp 18001
transform 1 0 18032 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1757_
timestamp 18001
transform 1 0 17940 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _1758_
timestamp 18001
transform -1 0 24932 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1759_
timestamp 18001
transform 1 0 17756 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1760_
timestamp 18001
transform -1 0 17940 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_4  _1761_
timestamp 18001
transform 1 0 24472 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__nand2_1  _1762_
timestamp 18001
transform -1 0 16928 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _1763_
timestamp 18001
transform -1 0 21528 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1764_
timestamp 18001
transform -1 0 18124 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1765_
timestamp 18001
transform 1 0 17020 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1766_
timestamp 18001
transform -1 0 28704 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1767_
timestamp 18001
transform 1 0 21620 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1768_
timestamp 18001
transform -1 0 20884 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1769_
timestamp 18001
transform 1 0 20884 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1770_
timestamp 18001
transform 1 0 18492 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1771_
timestamp 18001
transform 1 0 19688 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1772_
timestamp 18001
transform 1 0 17480 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1773_
timestamp 18001
transform -1 0 17572 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1774_
timestamp 18001
transform -1 0 17388 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1775_
timestamp 18001
transform -1 0 15180 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1776_
timestamp 18001
transform -1 0 25668 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1777_
timestamp 18001
transform 1 0 23736 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1778_
timestamp 18001
transform 1 0 25944 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1779_
timestamp 18001
transform 1 0 26404 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1780_
timestamp 18001
transform 1 0 23644 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1781_
timestamp 18001
transform 1 0 20056 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1782_
timestamp 18001
transform 1 0 19688 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1783_
timestamp 18001
transform 1 0 19872 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1784_
timestamp 18001
transform 1 0 24012 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1785_
timestamp 18001
transform -1 0 18768 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _1786_
timestamp 18001
transform 1 0 25668 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1787_
timestamp 18001
transform 1 0 16836 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1788_
timestamp 18001
transform -1 0 17020 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1789_
timestamp 18001
transform -1 0 21252 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1790_
timestamp 18001
transform 1 0 17572 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1791_
timestamp 18001
transform -1 0 23276 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1792_
timestamp 18001
transform 1 0 16928 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1793_
timestamp 18001
transform -1 0 17480 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1794_
timestamp 18001
transform -1 0 15824 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1795_
timestamp 18001
transform -1 0 23184 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1796_
timestamp 18001
transform 1 0 23184 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1797_
timestamp 18001
transform 1 0 21804 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1798_
timestamp 18001
transform 1 0 15364 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1799_
timestamp 18001
transform -1 0 8096 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1800_
timestamp 18001
transform -1 0 21252 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1801_
timestamp 18001
transform -1 0 22264 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1802_
timestamp 18001
transform 1 0 21988 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1803_
timestamp 18001
transform -1 0 22264 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1804_
timestamp 18001
transform -1 0 17940 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1805_
timestamp 18001
transform 1 0 27508 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _1806_
timestamp 18001
transform 1 0 27508 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _1807_
timestamp 18001
transform 1 0 24748 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1808_
timestamp 18001
transform -1 0 23092 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1809_
timestamp 18001
transform -1 0 21712 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1810_
timestamp 18001
transform -1 0 20792 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1811_
timestamp 18001
transform 1 0 22816 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1812_
timestamp 18001
transform -1 0 22540 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1813_
timestamp 18001
transform 1 0 21252 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1814_
timestamp 18001
transform -1 0 22632 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_2  _1815_
timestamp 18001
transform -1 0 23000 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _1816_
timestamp 18001
transform -1 0 22908 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_4  _1817_
timestamp 18001
transform 1 0 25852 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__a211oi_4  _1818_
timestamp 18001
transform -1 0 23552 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1819_
timestamp 18001
transform 1 0 12420 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_2  _1820_
timestamp 18001
transform -1 0 21620 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1821_
timestamp 18001
transform -1 0 21344 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1822_
timestamp 18001
transform -1 0 20884 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _1823_
timestamp 18001
transform -1 0 19136 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1824_
timestamp 18001
transform 1 0 20240 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1825_
timestamp 18001
transform -1 0 20056 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1826_
timestamp 18001
transform 1 0 19780 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1827_
timestamp 18001
transform 1 0 20240 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1828_
timestamp 18001
transform -1 0 27048 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1829_
timestamp 18001
transform -1 0 20884 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1830_
timestamp 18001
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1831_
timestamp 18001
transform 1 0 20884 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1832_
timestamp 18001
transform -1 0 20700 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1833_
timestamp 18001
transform -1 0 20884 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1834_
timestamp 18001
transform 1 0 23644 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1835_
timestamp 18001
transform 1 0 20148 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1836_
timestamp 18001
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1837_
timestamp 18001
transform 1 0 19504 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1838_
timestamp 18001
transform -1 0 19872 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1839_
timestamp 18001
transform 1 0 20148 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1840_
timestamp 18001
transform 1 0 19964 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _1841_
timestamp 18001
transform 1 0 19320 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_2  _1842_
timestamp 18001
transform 1 0 21804 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _1843_
timestamp 18001
transform 1 0 20884 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1844_
timestamp 18001
transform -1 0 19136 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1845_
timestamp 18001
transform -1 0 20240 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1846_
timestamp 18001
transform -1 0 19688 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_2  _1847_
timestamp 18001
transform -1 0 18308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nand4b_1  _1848_
timestamp 18001
transform 1 0 18216 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _1849_
timestamp 18001
transform -1 0 19044 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1850_
timestamp 18001
transform -1 0 24472 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1851_
timestamp 18001
transform -1 0 19320 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1852_
timestamp 18001
transform -1 0 17112 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1853_
timestamp 18001
transform 1 0 15916 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1854_
timestamp 18001
transform -1 0 16008 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1855_
timestamp 18001
transform 1 0 11500 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1856_
timestamp 18001
transform -1 0 17572 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _1857_
timestamp 18001
transform -1 0 19964 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1858_
timestamp 18001
transform 1 0 15180 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1859_
timestamp 18001
transform -1 0 18676 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _1860_
timestamp 18001
transform -1 0 19964 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1861_
timestamp 18001
transform -1 0 16100 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1862_
timestamp 18001
transform -1 0 12696 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1863_
timestamp 18001
transform 1 0 11224 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1864_
timestamp 18001
transform 1 0 12236 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1865_
timestamp 18001
transform -1 0 18492 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1866_
timestamp 18001
transform 1 0 19228 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1867_
timestamp 18001
transform -1 0 23828 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1868_
timestamp 18001
transform -1 0 19780 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _1869_
timestamp 18001
transform -1 0 19412 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_1  _1870_
timestamp 18001
transform -1 0 11408 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1871_
timestamp 18001
transform 1 0 9844 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1872_
timestamp 18001
transform -1 0 23276 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1873_
timestamp 18001
transform -1 0 16468 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1874_
timestamp 18001
transform -1 0 16008 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1875_
timestamp 18001
transform -1 0 15640 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1876_
timestamp 18001
transform -1 0 23552 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1877_
timestamp 18001
transform -1 0 24840 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1878_
timestamp 18001
transform -1 0 21252 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1879_
timestamp 18001
transform 1 0 19412 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1880_
timestamp 18001
transform 1 0 21252 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1881_
timestamp 18001
transform -1 0 23552 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1882_
timestamp 18001
transform 1 0 24104 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1883_
timestamp 18001
transform 1 0 22264 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1884_
timestamp 18001
transform 1 0 22816 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _1885_
timestamp 18001
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1886_
timestamp 18001
transform -1 0 14444 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1887_
timestamp 18001
transform 1 0 14260 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1888_
timestamp 18001
transform 1 0 28428 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _1889_
timestamp 18001
transform 1 0 27968 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1890_
timestamp 18001
transform 1 0 29716 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1891_
timestamp 18001
transform 1 0 29072 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _1892_
timestamp 18001
transform -1 0 29348 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1893_
timestamp 18001
transform -1 0 23920 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1894_
timestamp 18001
transform 1 0 18216 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _1895_
timestamp 18001
transform 1 0 29716 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _1896_
timestamp 18001
transform -1 0 19044 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1897_
timestamp 18001
transform -1 0 16008 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1898_
timestamp 18001
transform -1 0 15732 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1899_
timestamp 18001
transform -1 0 15180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1900_
timestamp 18001
transform -1 0 28428 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1901_
timestamp 18001
transform -1 0 28428 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1902_
timestamp 18001
transform 1 0 27600 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1903_
timestamp 18001
transform 1 0 29716 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1904_
timestamp 18001
transform 1 0 21344 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1905_
timestamp 18001
transform -1 0 20976 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1906_
timestamp 18001
transform 1 0 15180 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1907_
timestamp 18001
transform -1 0 14720 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1908_
timestamp 18001
transform -1 0 14996 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1909_
timestamp 18001
transform -1 0 14076 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_4  _1910_
timestamp 18001
transform -1 0 15456 0 -1 20672
box -38 -48 1326 592
use sky130_fd_sc_hd__o21a_1  _1911_
timestamp 18001
transform 1 0 14076 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1912_
timestamp 18001
transform -1 0 15364 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _1913_
timestamp 18001
transform -1 0 13616 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1914_
timestamp 18001
transform -1 0 13984 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _1915_
timestamp 18001
transform -1 0 14168 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _1916_
timestamp 18001
transform -1 0 13984 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1917_
timestamp 18001
transform -1 0 10764 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1918_
timestamp 18001
transform 1 0 10212 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1919_
timestamp 18001
transform -1 0 11408 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1920_
timestamp 18001
transform 1 0 11408 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1921_
timestamp 18001
transform 1 0 27876 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1922_
timestamp 18001
transform 1 0 27600 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1923_
timestamp 18001
transform 1 0 26956 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1924_
timestamp 18001
transform 1 0 28888 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1925_
timestamp 18001
transform -1 0 26864 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1926_
timestamp 18001
transform -1 0 26864 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1927_
timestamp 18001
transform -1 0 27876 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1928_
timestamp 18001
transform 1 0 26956 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1929_
timestamp 18001
transform 1 0 27232 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1930_
timestamp 18001
transform -1 0 28888 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1931_
timestamp 18001
transform -1 0 27876 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1932_
timestamp 18001
transform -1 0 27876 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1933_
timestamp 18001
transform -1 0 28336 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1934_
timestamp 18001
transform -1 0 27968 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1935_
timestamp 18001
transform 1 0 27968 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1936_
timestamp 18001
transform -1 0 23368 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1937_
timestamp 18001
transform -1 0 26220 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1938_
timestamp 18001
transform -1 0 26588 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1939_
timestamp 18001
transform -1 0 26220 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1940_
timestamp 18001
transform 1 0 20516 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1941_
timestamp 18001
transform -1 0 27048 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _1942_
timestamp 18001
transform 1 0 22908 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1943_
timestamp 18001
transform -1 0 23092 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1944_
timestamp 18001
transform 1 0 23276 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1945_
timestamp 18001
transform 1 0 25392 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1946_
timestamp 18001
transform -1 0 23828 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1947_
timestamp 18001
transform 1 0 23736 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1948_
timestamp 18001
transform 1 0 24380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1949_
timestamp 18001
transform -1 0 24932 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1950_
timestamp 18001
transform 1 0 24840 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1951_
timestamp 18001
transform 1 0 25668 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1952_
timestamp 18001
transform -1 0 26404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1953_
timestamp 18001
transform -1 0 24288 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _1954_
timestamp 18001
transform -1 0 18124 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1955_
timestamp 18001
transform -1 0 17940 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _1956_
timestamp 18001
transform -1 0 18584 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_1  _1957_
timestamp 18001
transform -1 0 23828 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1958_
timestamp 18001
transform -1 0 19596 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1959_
timestamp 18001
transform -1 0 20608 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _1960_
timestamp 18001
transform 1 0 19596 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_4  _1961_
timestamp 18001
transform 1 0 16192 0 1 29376
box -38 -48 1786 592
use sky130_fd_sc_hd__a221oi_2  _1962_
timestamp 18001
transform 1 0 14996 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _1963_
timestamp 18001
transform 1 0 11592 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1964_
timestamp 18001
transform 1 0 11500 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1965_
timestamp 18001
transform 1 0 10948 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1966_
timestamp 18001
transform -1 0 11224 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1967_
timestamp 18001
transform 1 0 17572 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1968_
timestamp 18001
transform -1 0 18032 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1969_
timestamp 18001
transform 1 0 18032 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1970_
timestamp 18001
transform -1 0 17388 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  _1971_
timestamp 18001
transform -1 0 18032 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _1972_
timestamp 18001
transform 1 0 16836 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1973_
timestamp 18001
transform 1 0 9384 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1974_
timestamp 18001
transform -1 0 16468 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1975_
timestamp 18001
transform 1 0 16744 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1976_
timestamp 18001
transform 1 0 16928 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1977_
timestamp 18001
transform 1 0 16560 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1978_
timestamp 18001
transform -1 0 16928 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1979_
timestamp 18001
transform 1 0 15824 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1980_
timestamp 18001
transform -1 0 15272 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1981_
timestamp 18001
transform 1 0 11684 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1982_
timestamp 18001
transform 1 0 12420 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1983_
timestamp 18001
transform -1 0 17940 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _1984_
timestamp 18001
transform -1 0 12328 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1985_
timestamp 18001
transform 1 0 18584 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1986_
timestamp 18001
transform 1 0 17756 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1987_
timestamp 18001
transform -1 0 26680 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1988_
timestamp 18001
transform 1 0 25208 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1989_
timestamp 18001
transform 1 0 23000 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1990_
timestamp 18001
transform -1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1991_
timestamp 18001
transform 1 0 23736 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1992_
timestamp 18001
transform 1 0 23000 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1993_
timestamp 18001
transform 1 0 23736 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1994_
timestamp 18001
transform 1 0 24196 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1995_
timestamp 18001
transform -1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1996_
timestamp 18001
transform -1 0 26588 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1997_
timestamp 18001
transform -1 0 23276 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1998_
timestamp 18001
transform -1 0 16652 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1999_
timestamp 18001
transform 1 0 16192 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2000_
timestamp 18001
transform 1 0 26220 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2001_
timestamp 18001
transform -1 0 26864 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_1  _2002_
timestamp 18001
transform 1 0 25944 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2003_
timestamp 18001
transform 1 0 16008 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _2004_
timestamp 18001
transform -1 0 17388 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _2005_
timestamp 18001
transform 1 0 17388 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _2006_
timestamp 18001
transform -1 0 16008 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _2007_
timestamp 18001
transform -1 0 16100 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _2008_
timestamp 18001
transform -1 0 15732 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2009_
timestamp 18001
transform -1 0 11408 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2010_
timestamp 18001
transform 1 0 10488 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _2011_
timestamp 18001
transform -1 0 15640 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2012_
timestamp 18001
transform 1 0 11500 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _2013_
timestamp 18001
transform 1 0 12236 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2014_
timestamp 18001
transform 1 0 11776 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2015_
timestamp 18001
transform 1 0 11500 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2016_
timestamp 18001
transform -1 0 12052 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2017_
timestamp 18001
transform 1 0 11316 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2018_
timestamp 18001
transform 1 0 12972 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _2019_
timestamp 18001
transform -1 0 12420 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2020_
timestamp 18001
transform 1 0 16652 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2021_
timestamp 18001
transform -1 0 17388 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2022_
timestamp 18001
transform -1 0 10764 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _2023_
timestamp 18001
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2024_
timestamp 18001
transform 1 0 6348 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2025_
timestamp 18001
transform -1 0 6256 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2026_
timestamp 18001
transform 1 0 4692 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2027_
timestamp 18001
transform -1 0 5980 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_2  _2028_
timestamp 18001
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__o2bb2a_1  _2029_
timestamp 18001
transform 1 0 10764 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _2030_
timestamp 18001
transform -1 0 10856 0 -1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _2031_
timestamp 18001
transform -1 0 9476 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2032_
timestamp 18001
transform 1 0 6348 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2033_
timestamp 18001
transform 1 0 8004 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _2034_
timestamp 18001
transform -1 0 9384 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_2  _2035_
timestamp 18001
transform 1 0 10580 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2036_
timestamp 18001
transform 1 0 10488 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2037_
timestamp 18001
transform -1 0 8832 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2038_
timestamp 18001
transform 1 0 9384 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _2039_
timestamp 18001
transform 1 0 9476 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _2040_
timestamp 18001
transform 1 0 10028 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _2041_
timestamp 18001
transform -1 0 10028 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2042_
timestamp 18001
transform 1 0 3404 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2043_
timestamp 18001
transform 1 0 5428 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2044_
timestamp 18001
transform 1 0 5520 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2045_
timestamp 18001
transform -1 0 6256 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_2  _2046_
timestamp 18001
transform 1 0 15088 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _2047_
timestamp 18001
transform -1 0 9936 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2048_
timestamp 18001
transform 1 0 13340 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2049_
timestamp 18001
transform -1 0 14720 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2050_
timestamp 18001
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2051_
timestamp 18001
transform 1 0 12972 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2052_
timestamp 18001
transform -1 0 12604 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _2053_
timestamp 18001
transform -1 0 9660 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _2054_
timestamp 18001
transform 1 0 9016 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2055_
timestamp 18001
transform -1 0 8188 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2056_
timestamp 18001
transform -1 0 12420 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2057_
timestamp 18001
transform 1 0 10672 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2058_
timestamp 18001
transform -1 0 8740 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2059_
timestamp 18001
transform -1 0 6992 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2060_
timestamp 18001
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _2061_
timestamp 18001
transform 1 0 6992 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2062_
timestamp 18001
transform 1 0 7084 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _2063_
timestamp 18001
transform 1 0 8004 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2064_
timestamp 18001
transform -1 0 8004 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2065_
timestamp 18001
transform 1 0 7820 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2066_
timestamp 18001
transform 1 0 6808 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2067_
timestamp 18001
transform 1 0 5704 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2068_
timestamp 18001
transform -1 0 7268 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _2069_
timestamp 18001
transform -1 0 6808 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_1  _2070_
timestamp 18001
transform 1 0 15180 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _2071_
timestamp 18001
transform 1 0 11500 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2072_
timestamp 18001
transform -1 0 14996 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2073_
timestamp 18001
transform -1 0 19504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _2074_
timestamp 18001
transform 1 0 18124 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2075_
timestamp 18001
transform -1 0 18216 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _2076_
timestamp 18001
transform 1 0 11684 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _2077_
timestamp 18001
transform 1 0 11500 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _2078_
timestamp 18001
transform -1 0 10764 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _2079_
timestamp 18001
transform -1 0 7820 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _2080_
timestamp 18001
transform 1 0 10948 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2081_
timestamp 18001
transform 1 0 11500 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2082_
timestamp 18001
transform 1 0 10488 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2083_
timestamp 18001
transform 1 0 5336 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2084_
timestamp 18001
transform 1 0 7084 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _2085_
timestamp 18001
transform -1 0 7176 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2086_
timestamp 18001
transform -1 0 7452 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2087_
timestamp 18001
transform -1 0 7728 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2088_
timestamp 18001
transform -1 0 7544 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2089_
timestamp 18001
transform -1 0 7084 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2090_
timestamp 18001
transform -1 0 7084 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2091_
timestamp 18001
transform -1 0 6992 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2092_
timestamp 18001
transform 1 0 6164 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2093_
timestamp 18001
transform 1 0 5336 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2094_
timestamp 18001
transform -1 0 6624 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _2095_
timestamp 18001
transform 1 0 6808 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_2  _2096_
timestamp 18001
transform 1 0 14904 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__o22ai_1  _2097_
timestamp 18001
transform -1 0 9844 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2098_
timestamp 18001
transform 1 0 13524 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2099_
timestamp 18001
transform -1 0 14812 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2100_
timestamp 18001
transform -1 0 10212 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2101_
timestamp 18001
transform 1 0 10120 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _2102_
timestamp 18001
transform 1 0 9384 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_2  _2103_
timestamp 18001
transform 1 0 10488 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2104_
timestamp 18001
transform 1 0 11776 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2105_
timestamp 18001
transform 1 0 9844 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2106_
timestamp 18001
transform 1 0 5612 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2107_
timestamp 18001
transform 1 0 5980 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _2108_
timestamp 18001
transform -1 0 6900 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2109_
timestamp 18001
transform 1 0 6072 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2110_
timestamp 18001
transform 1 0 8924 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor3b_1  _2111_
timestamp 18001
transform 1 0 7452 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2112_
timestamp 18001
transform 1 0 15364 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2113_
timestamp 18001
transform 1 0 16100 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2114_
timestamp 18001
transform -1 0 10396 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _2115_
timestamp 18001
transform 1 0 10580 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2116_
timestamp 18001
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2117_
timestamp 18001
transform -1 0 6992 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2118_
timestamp 18001
transform 1 0 5612 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_4  _2119_
timestamp 18001
transform 1 0 5980 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__a221oi_2  _2120_
timestamp 18001
transform 1 0 15088 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _2121_
timestamp 18001
transform -1 0 10488 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _2122_
timestamp 18001
transform 1 0 10212 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2123_
timestamp 18001
transform 1 0 9660 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _2124_
timestamp 18001
transform -1 0 10948 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2125_
timestamp 18001
transform 1 0 11960 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2126_
timestamp 18001
transform -1 0 12788 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2127_
timestamp 18001
transform 1 0 11316 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2128_
timestamp 18001
transform -1 0 15732 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2129_
timestamp 18001
transform -1 0 8556 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _2130_
timestamp 18001
transform 1 0 8004 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2131_
timestamp 18001
transform 1 0 9200 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _2132_
timestamp 18001
transform 1 0 10396 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _2133_
timestamp 18001
transform 1 0 12788 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2134_
timestamp 18001
transform 1 0 13616 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _2135_
timestamp 18001
transform -1 0 14812 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2136_
timestamp 18001
transform -1 0 13616 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2137_
timestamp 18001
transform -1 0 14444 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2138_
timestamp 18001
transform -1 0 8096 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2139_
timestamp 18001
transform -1 0 9200 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2140_
timestamp 18001
transform 1 0 8096 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2141_
timestamp 18001
transform -1 0 9016 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_4  _2142_
timestamp 18001
transform 1 0 15088 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__o2bb2a_1  _2143_
timestamp 18001
transform 1 0 14076 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _2144_
timestamp 18001
transform 1 0 12788 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _2145_
timestamp 18001
transform -1 0 12880 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _2146_
timestamp 18001
transform -1 0 14904 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2147_
timestamp 18001
transform -1 0 13984 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2148_
timestamp 18001
transform 1 0 13156 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2149_
timestamp 18001
transform 1 0 8924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2150_
timestamp 18001
transform -1 0 11500 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2151_
timestamp 18001
transform -1 0 9844 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _2152_
timestamp 18001
transform 1 0 8924 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2153_
timestamp 18001
transform 1 0 7360 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _2154_
timestamp 18001
transform -1 0 13156 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2155_
timestamp 18001
transform -1 0 12052 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2156_
timestamp 18001
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_2  _2157_
timestamp 18001
transform -1 0 13340 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__a22oi_1  _2158_
timestamp 18001
transform -1 0 13248 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2159_
timestamp 18001
transform -1 0 12972 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2160_
timestamp 18001
transform -1 0 12972 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2161_
timestamp 18001
transform -1 0 17204 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _2162_
timestamp 18001
transform 1 0 16008 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2163_
timestamp 18001
transform 1 0 16652 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2164_
timestamp 18001
transform 1 0 14352 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2165_
timestamp 18001
transform -1 0 15548 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_1  _2166_
timestamp 18001
transform 1 0 14260 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _2167_
timestamp 18001
transform 1 0 16836 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2168_
timestamp 18001
transform 1 0 14628 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2169_
timestamp 18001
transform -1 0 14352 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _2170_
timestamp 18001
transform 1 0 13064 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _2171_
timestamp 18001
transform -1 0 13708 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2172_
timestamp 18001
transform -1 0 14260 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2173_
timestamp 18001
transform 1 0 14628 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2174_
timestamp 18001
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2175_
timestamp 18001
transform -1 0 14260 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _2176_
timestamp 18001
transform -1 0 14628 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _2177_
timestamp 18001
transform -1 0 14812 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_1  _2178_
timestamp 18001
transform 1 0 14444 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _2179_
timestamp 18001
transform -1 0 17204 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _2180_
timestamp 18001
transform 1 0 14904 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2181_
timestamp 18001
transform -1 0 9200 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2182_
timestamp 18001
transform -1 0 14076 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _2183_
timestamp 18001
transform 1 0 13156 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _2184_
timestamp 18001
transform -1 0 14260 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _2185_
timestamp 18001
transform -1 0 13616 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _2186_
timestamp 18001
transform 1 0 12788 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _2187_
timestamp 18001
transform -1 0 22540 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2188_
timestamp 18001
transform -1 0 21528 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2189_
timestamp 18001
transform -1 0 20976 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _2190_
timestamp 18001
transform -1 0 24748 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2191_
timestamp 18001
transform -1 0 21620 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _2192_
timestamp 18001
transform -1 0 21620 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2193_
timestamp 18001
transform 1 0 26956 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2194_
timestamp 18001
transform -1 0 22264 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2195_
timestamp 18001
transform 1 0 20976 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2196_
timestamp 18001
transform 1 0 20516 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2197_
timestamp 18001
transform -1 0 19872 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2198_
timestamp 18001
transform 1 0 12420 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _2199_
timestamp 18001
transform -1 0 12696 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _2200_
timestamp 18001
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2201_
timestamp 18001
transform 1 0 9844 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2202_
timestamp 18001
transform 1 0 10304 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2203_
timestamp 18001
transform 1 0 9200 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _2204_
timestamp 18001
transform -1 0 8740 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _2205_
timestamp 18001
transform 1 0 7268 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2206_
timestamp 18001
transform 1 0 6716 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2207_
timestamp 18001
transform 1 0 6256 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2208_
timestamp 18001
transform -1 0 6256 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2209_
timestamp 18001
transform 1 0 7544 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2210_
timestamp 18001
transform -1 0 9200 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2211_
timestamp 18001
transform 1 0 11316 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _2212_
timestamp 18001
transform -1 0 11408 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2213_
timestamp 18001
transform -1 0 15180 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2214_
timestamp 18001
transform 1 0 14260 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _2215_
timestamp 18001
transform -1 0 14996 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _2216_
timestamp 18001
transform -1 0 14904 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_2  _2217_
timestamp 18001
transform 1 0 19780 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2218_
timestamp 18001
transform 1 0 12512 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2219_
timestamp 18001
transform 1 0 11592 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2220_
timestamp 18001
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _2221_
timestamp 18001
transform -1 0 10304 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _2222_
timestamp 18001
transform -1 0 11500 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _2223_
timestamp 18001
transform 1 0 5060 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2224_
timestamp 18001
transform -1 0 7360 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _2225_
timestamp 18001
transform -1 0 5612 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _2226_
timestamp 18001
transform 1 0 6900 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _2227_
timestamp 18001
transform -1 0 5060 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2228_
timestamp 18001
transform 1 0 6992 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2229_
timestamp 18001
transform -1 0 8648 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _2230_
timestamp 18001
transform 1 0 9476 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2231_
timestamp 18001
transform -1 0 8464 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _2232_
timestamp 18001
transform 1 0 7544 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2233_
timestamp 18001
transform 1 0 6992 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2234_
timestamp 18001
transform 1 0 8556 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _2235_
timestamp 18001
transform 1 0 10764 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _2236_
timestamp 18001
transform -1 0 12696 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _2237_
timestamp 18001
transform -1 0 8464 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2238_
timestamp 18001
transform 1 0 10948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2239_
timestamp 18001
transform 1 0 10304 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _2240_
timestamp 18001
transform -1 0 11224 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2241_
timestamp 18001
transform -1 0 18400 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2242_
timestamp 18001
transform 1 0 20608 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _2243_
timestamp 18001
transform -1 0 18952 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _2244_
timestamp 18001
transform 1 0 16928 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2245_
timestamp 18001
transform 1 0 17204 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2246_
timestamp 18001
transform -1 0 16928 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2247_
timestamp 18001
transform 1 0 15364 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2248_
timestamp 18001
transform 1 0 22264 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _2249_
timestamp 18001
transform 1 0 22080 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _2250_
timestamp 18001
transform 1 0 19964 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2251_
timestamp 18001
transform -1 0 15456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2252_
timestamp 18001
transform 1 0 14536 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2253_
timestamp 18001
transform 1 0 12052 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _2254_
timestamp 18001
transform 1 0 14076 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _2255_
timestamp 18001
transform 1 0 13248 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2256_
timestamp 18001
transform -1 0 15732 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _2257_
timestamp 18001
transform 1 0 18400 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2258_
timestamp 18001
transform -1 0 21712 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2259_
timestamp 18001
transform 1 0 18400 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2260_
timestamp 18001
transform -1 0 14628 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_2  _2261_
timestamp 18001
transform 1 0 30084 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _2262_
timestamp 18001
transform 1 0 14812 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _2263_
timestamp 18001
transform -1 0 15916 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2264_
timestamp 18001
transform 1 0 11500 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2265_
timestamp 18001
transform -1 0 12972 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _2266_
timestamp 18001
transform 1 0 14536 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2267_
timestamp 18001
transform 1 0 17940 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _2268_
timestamp 18001
transform 1 0 17020 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _2269_
timestamp 18001
transform 1 0 18492 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2270_
timestamp 18001
transform 1 0 15916 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _2271_
timestamp 18001
transform -1 0 15732 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _2272_
timestamp 18001
transform 1 0 23184 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _2273_
timestamp 18001
transform -1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2274_
timestamp 18001
transform 1 0 18492 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2275_
timestamp 18001
transform -1 0 21160 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2276_
timestamp 18001
transform -1 0 20700 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2277_
timestamp 18001
transform 1 0 19688 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2278_
timestamp 18001
transform -1 0 29256 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2279_
timestamp 18001
transform 1 0 19320 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2280_
timestamp 18001
transform 1 0 19596 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _2281_
timestamp 18001
transform 1 0 18308 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2282_
timestamp 18001
transform 1 0 17020 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _2283_
timestamp 18001
transform 1 0 20884 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2284_
timestamp 18001
transform -1 0 20516 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2285_
timestamp 18001
transform 1 0 19780 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2286_
timestamp 18001
transform -1 0 19136 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2287_
timestamp 18001
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2288_
timestamp 18001
transform -1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2289_
timestamp 18001
transform 1 0 18216 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2290_
timestamp 18001
transform 1 0 18216 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_4  _2291_
timestamp 18001
transform 1 0 19228 0 1 20672
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _2292_
timestamp 18001
transform 1 0 16652 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2293_
timestamp 18001
transform 1 0 14352 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2294_
timestamp 18001
transform 1 0 12328 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2295_
timestamp 18001
transform 1 0 11500 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2296_
timestamp 18001
transform 1 0 12512 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2297_
timestamp 18001
transform 1 0 12328 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2298_
timestamp 18001
transform 1 0 11500 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2299_
timestamp 18001
transform 1 0 14260 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _2300_
timestamp 18001
transform 1 0 25116 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _2301_
timestamp 18001
transform 1 0 25208 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _2302_
timestamp 18001
transform 1 0 24932 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2303_
timestamp 18001
transform 1 0 24472 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2304_
timestamp 18001
transform 1 0 24564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2305_
timestamp 18001
transform -1 0 26220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2306_
timestamp 18001
transform 1 0 25392 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2307_
timestamp 18001
transform -1 0 27600 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2308_
timestamp 18001
transform 1 0 26588 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _2309_
timestamp 18001
transform -1 0 29348 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _2310_
timestamp 18001
transform 1 0 24932 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2311_
timestamp 18001
transform 1 0 25116 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _2312_
timestamp 18001
transform 1 0 25576 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _2313_
timestamp 18001
transform -1 0 26588 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2314_
timestamp 18001
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2315_
timestamp 18001
transform 1 0 24288 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2316_
timestamp 18001
transform 1 0 24840 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _2317_
timestamp 18001
transform -1 0 23736 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2318_
timestamp 18001
transform -1 0 23644 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _2319_
timestamp 18001
transform 1 0 22816 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _2320_
timestamp 18001
transform 1 0 22540 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2321_
timestamp 18001
transform 1 0 22172 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _2322_
timestamp 18001
transform 1 0 22448 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2323_
timestamp 18001
transform 1 0 15548 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2324_
timestamp 18001
transform 1 0 15272 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2325_
timestamp 18001
transform 1 0 22264 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2326_
timestamp 18001
transform -1 0 11776 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2327_
timestamp 18001
transform 1 0 11776 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2328_
timestamp 18001
transform -1 0 12512 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2329_
timestamp 18001
transform -1 0 11592 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2330_
timestamp 18001
transform 1 0 11500 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2331_
timestamp 18001
transform 1 0 10120 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2332_
timestamp 18001
transform -1 0 10028 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2333_
timestamp 18001
transform 1 0 10212 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2334_
timestamp 18001
transform -1 0 9108 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2335_
timestamp 18001
transform -1 0 9384 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2336_
timestamp 18001
transform 1 0 9384 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2337_
timestamp 18001
transform 1 0 8464 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2338_
timestamp 18001
transform -1 0 8280 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2339_
timestamp 18001
transform 1 0 9292 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2340_
timestamp 18001
transform 1 0 8372 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2341_
timestamp 18001
transform 1 0 9200 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2342_
timestamp 18001
transform -1 0 9200 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2343_
timestamp 18001
transform 1 0 9476 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2344_
timestamp 18001
transform -1 0 10212 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2345_
timestamp 18001
transform -1 0 10580 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2346_
timestamp 18001
transform -1 0 11408 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2347_
timestamp 18001
transform 1 0 12052 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2348_
timestamp 18001
transform -1 0 13156 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2349_
timestamp 18001
transform 1 0 10396 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2350_
timestamp 18001
transform 1 0 9200 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2351_
timestamp 18001
transform 1 0 8280 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2352_
timestamp 18001
transform 1 0 8924 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2353_
timestamp 18001
transform -1 0 9476 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2354_
timestamp 18001
transform -1 0 12052 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2355_
timestamp 18001
transform -1 0 12420 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _2356_
timestamp 18001
transform 1 0 12420 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2357_
timestamp 18001
transform 1 0 12788 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _2358_
timestamp 18001
transform -1 0 8096 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2359_
timestamp 18001
transform -1 0 7452 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2360_
timestamp 18001
transform 1 0 7360 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2361_
timestamp 18001
transform 1 0 8924 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_2  _2362_
timestamp 18001
transform 1 0 18216 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _2363_
timestamp 18001
transform -1 0 13340 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _2364_
timestamp 18001
transform -1 0 11960 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2365_
timestamp 18001
transform 1 0 13064 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2366_
timestamp 18001
transform 1 0 13708 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _2367_
timestamp 18001
transform 1 0 12512 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _2368_
timestamp 18001
transform 1 0 5336 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2369_
timestamp 18001
transform -1 0 6808 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2370_
timestamp 18001
transform 1 0 6256 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2371_
timestamp 18001
transform 1 0 11868 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2372_
timestamp 18001
transform -1 0 12604 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2373_
timestamp 18001
transform 1 0 15180 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _2374_
timestamp 18001
transform 1 0 11960 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2375_
timestamp 18001
transform 1 0 12604 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _2376_
timestamp 18001
transform -1 0 16560 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2377_
timestamp 18001
transform 1 0 5980 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2378_
timestamp 18001
transform 1 0 12604 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2379_
timestamp 18001
transform -1 0 13708 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _2380_
timestamp 18001
transform -1 0 14996 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2381_
timestamp 18001
transform 1 0 13708 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2382_
timestamp 18001
transform 1 0 13340 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _2383_
timestamp 18001
transform 1 0 13708 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_4  _2384_
timestamp 18001
transform -1 0 15456 0 -1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__and4_1  _2385_
timestamp 18001
transform 1 0 12420 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _2386_
timestamp 18001
transform 1 0 13340 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2387_
timestamp 18001
transform 1 0 12696 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2388_
timestamp 18001
transform -1 0 14904 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2389_
timestamp 18001
transform 1 0 14076 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _2390_
timestamp 18001
transform -1 0 16008 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2391_
timestamp 18001
transform 1 0 16008 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2392_
timestamp 18001
transform 1 0 14260 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2393_
timestamp 18001
transform -1 0 16284 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _2394_
timestamp 18001
transform 1 0 14996 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2395_
timestamp 18001
transform 1 0 15548 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2396_
timestamp 18001
transform 1 0 15088 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2397_
timestamp 18001
transform 1 0 14904 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _2398_
timestamp 18001
transform 1 0 15640 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2399_
timestamp 18001
transform -1 0 11408 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _2400_
timestamp 18001
transform 1 0 10580 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_1  _2401_
timestamp 18001
transform 1 0 15548 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2402_
timestamp 18001
transform -1 0 14996 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2403_
timestamp 18001
transform -1 0 16284 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _2404_
timestamp 18001
transform -1 0 18216 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2405_
timestamp 18001
transform 1 0 16284 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2406_
timestamp 18001
transform 1 0 16928 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _2407_
timestamp 18001
transform -1 0 17204 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nand4b_1  _2408_
timestamp 18001
transform 1 0 15548 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2409_
timestamp 18001
transform 1 0 17572 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _2410_
timestamp 18001
transform 1 0 10856 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_2  _2411_
timestamp 18001
transform 1 0 11776 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2412_
timestamp 18001
transform 1 0 18400 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2413_
timestamp 18001
transform -1 0 17572 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2414_
timestamp 18001
transform -1 0 18124 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _2415_
timestamp 18001
transform 1 0 17756 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2416_
timestamp 18001
transform 1 0 20700 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2417_
timestamp 18001
transform 1 0 21252 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2418_
timestamp 18001
transform -1 0 21804 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2419_
timestamp 18001
transform -1 0 21804 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2420_
timestamp 18001
transform 1 0 16652 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _2421_
timestamp 18001
transform -1 0 16652 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2422_
timestamp 18001
transform 1 0 16652 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2423_
timestamp 18001
transform -1 0 21068 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2424_
timestamp 18001
transform 1 0 17848 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2425_
timestamp 18001
transform -1 0 18860 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2426_
timestamp 18001
transform -1 0 11040 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_4  _2427_
timestamp 18001
transform 1 0 11500 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__inv_2  _2428_
timestamp 18001
transform 1 0 22908 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _2429_
timestamp 18001
transform -1 0 19780 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2430_
timestamp 18001
transform 1 0 18676 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2431_
timestamp 18001
transform 1 0 18952 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _2432_
timestamp 18001
transform -1 0 22172 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2433_
timestamp 18001
transform -1 0 22724 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2434_
timestamp 18001
transform 1 0 20976 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2435_
timestamp 18001
transform -1 0 22540 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2436_
timestamp 18001
transform -1 0 22172 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2437_
timestamp 18001
transform 1 0 12696 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _2438_
timestamp 18001
transform -1 0 12788 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2439_
timestamp 18001
transform 1 0 18124 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2440_
timestamp 18001
transform 1 0 16192 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2441_
timestamp 18001
transform -1 0 17664 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2442_
timestamp 18001
transform 1 0 18308 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2443_
timestamp 18001
transform 1 0 17664 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _2444_
timestamp 18001
transform 1 0 19044 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _2445_
timestamp 18001
transform 1 0 20976 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _2446_
timestamp 18001
transform -1 0 21712 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2447_
timestamp 18001
transform 1 0 20700 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2448_
timestamp 18001
transform -1 0 22264 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2449_
timestamp 18001
transform 1 0 16744 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2450_
timestamp 18001
transform -1 0 18584 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2451_
timestamp 18001
transform 1 0 11040 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _2452_
timestamp 18001
transform 1 0 11224 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2453_
timestamp 18001
transform 1 0 18584 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2454_
timestamp 18001
transform -1 0 18768 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _2455_
timestamp 18001
transform 1 0 18768 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _2456_
timestamp 18001
transform 1 0 21804 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2457_
timestamp 18001
transform 1 0 19596 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2458_
timestamp 18001
transform -1 0 20700 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _2459_
timestamp 18001
transform 1 0 17296 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2460_
timestamp 18001
transform -1 0 17664 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2461_
timestamp 18001
transform 1 0 12052 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _2462_
timestamp 18001
transform 1 0 11868 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _2463_
timestamp 18001
transform 1 0 17020 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2464_
timestamp 18001
transform -1 0 17940 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2465_
timestamp 18001
transform 1 0 17572 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _2466_
timestamp 18001
transform -1 0 22724 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_4  _2467_
timestamp 18001
transform 1 0 21620 0 1 17408
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _2468_
timestamp 18001
transform 1 0 12604 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2469_
timestamp 18001
transform 1 0 7912 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2470_
timestamp 18001
transform 1 0 4600 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2471_
timestamp 18001
transform 1 0 2576 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2472_
timestamp 18001
transform 1 0 4508 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2473_
timestamp 18001
transform 1 0 2668 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2474_
timestamp 18001
transform 1 0 2484 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2475_
timestamp 18001
transform -1 0 10212 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _2476_
timestamp 18001
transform 1 0 29624 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _2477_
timestamp 18001
transform -1 0 29256 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _2478_
timestamp 18001
transform 1 0 15732 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2479_
timestamp 18001
transform 1 0 11776 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2480_
timestamp 18001
transform 1 0 7636 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2481_
timestamp 18001
transform 1 0 3956 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2482_
timestamp 18001
transform 1 0 4784 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2483_
timestamp 18001
transform 1 0 4416 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2484_
timestamp 18001
transform 1 0 2668 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2485_
timestamp 18001
transform 1 0 2208 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2486_
timestamp 18001
transform 1 0 9292 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2487_
timestamp 18001
transform 1 0 21620 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2488_
timestamp 18001
transform -1 0 23184 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a2111oi_1  _2489_
timestamp 18001
transform 1 0 26128 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _2490_
timestamp 18001
transform -1 0 26128 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _2491_
timestamp 18001
transform -1 0 29164 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2492_
timestamp 18001
transform -1 0 28428 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2493_
timestamp 18001
transform 1 0 28060 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _2494_
timestamp 18001
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _2495_
timestamp 18001
transform -1 0 26864 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2496_
timestamp 18001
transform 1 0 26588 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2497_
timestamp 18001
transform 1 0 26128 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a22oi_1  _2498_
timestamp 18001
transform 1 0 24656 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_2  _2499_
timestamp 18001
transform 1 0 25668 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2500_
timestamp 18001
transform 1 0 25392 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2501_
timestamp 18001
transform -1 0 26220 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2502_
timestamp 18001
transform 1 0 23000 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2503_
timestamp 18001
transform 1 0 24932 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2504_
timestamp 18001
transform 1 0 23184 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2505_
timestamp 18001
transform 1 0 23460 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2506_
timestamp 18001
transform 1 0 25300 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2507_
timestamp 18001
transform 1 0 24380 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2508_
timestamp 18001
transform 1 0 14168 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2509_
timestamp 18001
transform 1 0 14168 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2510_
timestamp 18001
transform -1 0 8280 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2511_
timestamp 18001
transform -1 0 8832 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2512_
timestamp 18001
transform -1 0 8648 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2513_
timestamp 18001
transform 1 0 8096 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2514_
timestamp 18001
transform -1 0 12052 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2515_
timestamp 18001
transform 1 0 12052 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2516_
timestamp 18001
transform -1 0 11408 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2517_
timestamp 18001
transform -1 0 8004 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2518_
timestamp 18001
transform -1 0 8372 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _2519_
timestamp 18001
transform -1 0 10672 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2520_
timestamp 18001
transform -1 0 10304 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _2521_
timestamp 18001
transform -1 0 7636 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2522_
timestamp 18001
transform 1 0 7636 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2523_
timestamp 18001
transform 1 0 6072 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _2524_
timestamp 18001
transform -1 0 10212 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _2525_
timestamp 18001
transform -1 0 9476 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2526_
timestamp 18001
transform 1 0 5520 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2527_
timestamp 18001
transform 1 0 6348 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2528_
timestamp 18001
transform 1 0 5152 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2529_
timestamp 18001
transform -1 0 8924 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _2530_
timestamp 18001
transform 1 0 8924 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2531_
timestamp 18001
transform 1 0 6348 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _2532_
timestamp 18001
transform 1 0 5980 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2533_
timestamp 18001
transform 1 0 5152 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2534_
timestamp 18001
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2535_
timestamp 18001
transform -1 0 7084 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2536_
timestamp 18001
transform 1 0 6900 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _2537_
timestamp 18001
transform 1 0 6716 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2538_
timestamp 18001
transform 1 0 6348 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2539_
timestamp 18001
transform 1 0 5152 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _2540_
timestamp 18001
transform 1 0 5520 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _2541_
timestamp 18001
transform 1 0 8464 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _2542_
timestamp 18001
transform 1 0 8096 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _2543_
timestamp 18001
transform 1 0 5704 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _2544_
timestamp 18001
transform -1 0 8096 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _2545_
timestamp 18001
transform 1 0 8280 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2546_
timestamp 18001
transform 1 0 5888 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2547_
timestamp 18001
transform -1 0 7728 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2548_
timestamp 18001
transform 1 0 7912 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2549_
timestamp 18001
transform 1 0 6808 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2550_
timestamp 18001
transform 1 0 7268 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2551_
timestamp 18001
transform 1 0 7728 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2552_
timestamp 18001
transform -1 0 8832 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2553_
timestamp 18001
transform -1 0 11500 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _2554_
timestamp 18001
transform 1 0 10580 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _2555_
timestamp 18001
transform 1 0 9568 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2556_
timestamp 18001
transform 1 0 10488 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2557_
timestamp 18001
transform -1 0 11224 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _2558_
timestamp 18001
transform 1 0 10488 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2559_
timestamp 18001
transform 1 0 24564 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2560_
timestamp 18001
transform 1 0 29624 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_4  _2561_
timestamp 18001
transform 1 0 24380 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _2562_
timestamp 18001
transform 1 0 12788 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2563_
timestamp 18001
transform 1 0 7544 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2564_
timestamp 18001
transform 1 0 6348 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2565_
timestamp 18001
transform 1 0 4324 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2566_
timestamp 18001
transform 1 0 5612 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2567_
timestamp 18001
transform 1 0 3956 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2568_
timestamp 18001
transform 1 0 4140 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2569_
timestamp 18001
transform 1 0 8372 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2570_
timestamp 18001
transform -1 0 27968 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2571_
timestamp 18001
transform 1 0 27876 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2572_
timestamp 18001
transform 1 0 28244 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _2573_
timestamp 18001
transform -1 0 28244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2574_
timestamp 18001
transform 1 0 27232 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _2575_
timestamp 18001
transform -1 0 25760 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__a221oi_2  _2576_
timestamp 18001
transform -1 0 24196 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _2577_
timestamp 18001
transform 1 0 24196 0 -1 31552
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _2578_
timestamp 18001
transform 1 0 2760 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2579_
timestamp 18001
transform 1 0 4140 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _2580_
timestamp 18001
transform 1 0 2668 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2581_
timestamp 18001
transform -1 0 2760 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2582_
timestamp 18001
transform 1 0 3036 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2583_
timestamp 18001
transform 1 0 5244 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2584_
timestamp 18001
transform 1 0 1932 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2585_
timestamp 18001
transform 1 0 3772 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _2586_
timestamp 18001
transform 1 0 12880 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2587_
timestamp 18001
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2588_
timestamp 18001
transform -1 0 15456 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2589_
timestamp 18001
transform -1 0 15088 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2590_
timestamp 18001
transform -1 0 17572 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _2591_
timestamp 18001
transform -1 0 19136 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _2592_
timestamp 18001
transform -1 0 16008 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2593_
timestamp 18001
transform 1 0 13708 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _2594_
timestamp 18001
transform -1 0 13708 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _2595_
timestamp 18001
transform 1 0 12788 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _2596_
timestamp 18001
transform 1 0 13708 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _2597_
timestamp 18001
transform 1 0 19780 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _2598_
timestamp 18001
transform -1 0 18124 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2599_
timestamp 18001
transform -1 0 16376 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _2600_
timestamp 18001
transform -1 0 16468 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _2601_
timestamp 18001
transform -1 0 16376 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _2602_
timestamp 18001
transform 1 0 14812 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2603_
timestamp 18001
transform 1 0 4784 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2604_
timestamp 18001
transform 1 0 7544 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _2605_
timestamp 18001
transform 1 0 12512 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _2606_
timestamp 18001
transform 1 0 10212 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2607_
timestamp 18001
transform 1 0 11040 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _2608_
timestamp 18001
transform 1 0 10580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _2609_
timestamp 18001
transform 1 0 7360 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2610_
timestamp 18001
transform 1 0 3772 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2611_
timestamp 18001
transform -1 0 4876 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2612_
timestamp 18001
transform 1 0 4140 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _2613_
timestamp 18001
transform -1 0 14812 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2614_
timestamp 18001
transform -1 0 4784 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2615_
timestamp 18001
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2616_
timestamp 18001
transform 1 0 4140 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2617_
timestamp 18001
transform -1 0 10304 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2618_
timestamp 18001
transform 1 0 9844 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2619_
timestamp 18001
transform -1 0 10028 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _2620_
timestamp 18001
transform 1 0 9108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2621_
timestamp 18001
transform -1 0 5428 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2622_
timestamp 18001
transform 1 0 3956 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2623_
timestamp 18001
transform 1 0 5520 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2624_
timestamp 18001
transform 1 0 5612 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _2625_
timestamp 18001
transform 1 0 6164 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _2626_
timestamp 18001
transform -1 0 6808 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2627_
timestamp 18001
transform 1 0 8188 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2628_
timestamp 18001
transform 1 0 7820 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2629_
timestamp 18001
transform 1 0 8096 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _2630_
timestamp 18001
transform 1 0 5428 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2631_
timestamp 18001
transform 1 0 5796 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o22ai_1  _2632_
timestamp 18001
transform 1 0 6992 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2633_
timestamp 18001
transform 1 0 7176 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2634_
timestamp 18001
transform 1 0 6256 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2635_
timestamp 18001
transform 1 0 4048 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2636_
timestamp 18001
transform -1 0 5520 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2637_
timestamp 18001
transform 1 0 4784 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2638_
timestamp 18001
transform -1 0 9200 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2639_
timestamp 18001
transform 1 0 8464 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _2640_
timestamp 18001
transform 1 0 8096 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2641_
timestamp 18001
transform 1 0 8004 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _2642_
timestamp 18001
transform -1 0 7544 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2643_
timestamp 18001
transform 1 0 7268 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2644_
timestamp 18001
transform 1 0 7912 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _2645_
timestamp 18001
transform -1 0 7268 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2646_
timestamp 18001
transform 1 0 6440 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2647_
timestamp 18001
transform 1 0 5152 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _2648_
timestamp 18001
transform 1 0 8372 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2649_
timestamp 18001
transform -1 0 10304 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2650_
timestamp 18001
transform -1 0 10304 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2651_
timestamp 18001
transform -1 0 10948 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2652_
timestamp 18001
transform 1 0 9568 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2653_
timestamp 18001
transform 1 0 8924 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2654_
timestamp 18001
transform -1 0 8004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _2655_
timestamp 18001
transform 1 0 7544 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2656_
timestamp 18001
transform -1 0 7544 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2657_
timestamp 18001
transform 1 0 6532 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _2658_
timestamp 18001
transform 1 0 7176 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2659_
timestamp 18001
transform -1 0 6992 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2660_
timestamp 18001
transform 1 0 12696 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2661_
timestamp 18001
transform 1 0 12420 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2662_
timestamp 18001
transform 1 0 12236 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2663_
timestamp 18001
transform -1 0 12972 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2664_
timestamp 18001
transform 1 0 12420 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2665_
timestamp 18001
transform 1 0 12972 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2666_
timestamp 18001
transform -1 0 10948 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_1  _2667_
timestamp 18001
transform -1 0 8556 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2668_
timestamp 18001
transform 1 0 9476 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2669_
timestamp 18001
transform 1 0 25576 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_4  _2670_
timestamp 18001
transform 1 0 24748 0 1 16320
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _2671_
timestamp 18001
transform 1 0 11684 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2672_
timestamp 18001
transform 1 0 7636 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2673_
timestamp 18001
transform 1 0 4324 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2674_
timestamp 18001
transform 1 0 3496 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2675_
timestamp 18001
transform 1 0 6348 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2676_
timestamp 18001
transform 1 0 3772 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2677_
timestamp 18001
transform 1 0 2668 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2678_
timestamp 18001
transform 1 0 9476 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _2679_
timestamp 18001
transform -1 0 18768 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _2680_
timestamp 18001
transform 1 0 17940 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _2681_
timestamp 18001
transform -1 0 30176 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2682_
timestamp 18001
transform -1 0 30544 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _2683_
timestamp 18001
transform 1 0 19320 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2684_
timestamp 18001
transform 1 0 16744 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _2685_
timestamp 18001
transform 1 0 31740 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2686_
timestamp 18001
transform 1 0 38456 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2687_
timestamp 18001
transform -1 0 32568 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2688_
timestamp 18001
transform -1 0 28796 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2689_
timestamp 18001
transform -1 0 38180 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2690_
timestamp 18001
transform -1 0 30268 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2691_
timestamp 18001
transform 1 0 38180 0 -1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2692_
timestamp 18001
transform 1 0 38180 0 -1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2693_
timestamp 18001
transform 1 0 32108 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2694_
timestamp 18001
transform 1 0 29900 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2695_
timestamp 18001
transform -1 0 36432 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2696_
timestamp 18001
transform -1 0 29256 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2697_
timestamp 18001
transform -1 0 36800 0 1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _2698_
timestamp 18001
transform 1 0 28796 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2699_
timestamp 18001
transform 1 0 24656 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2700_
timestamp 18001
transform 1 0 26956 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2701_
timestamp 18001
transform -1 0 31372 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2702_
timestamp 18001
transform -1 0 31280 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2703_
timestamp 18001
transform 1 0 24748 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2704_
timestamp 18001
transform -1 0 28796 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2705_
timestamp 18001
transform -1 0 21160 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2706_
timestamp 18001
transform 1 0 38272 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2707_
timestamp 18001
transform -1 0 39744 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2708_
timestamp 18001
transform -1 0 38180 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2709_
timestamp 18001
transform 1 0 38456 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2710_
timestamp 18001
transform 1 0 38180 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2711_
timestamp 18001
transform 1 0 36708 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2712_
timestamp 18001
transform 1 0 16008 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2713_
timestamp 18001
transform 1 0 12696 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2714_
timestamp 18001
transform -1 0 19688 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2715_
timestamp 18001
transform -1 0 15180 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2716_
timestamp 18001
transform 1 0 15088 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2717_
timestamp 18001
transform 1 0 19320 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_2  _2718_
timestamp 18001
transform 1 0 28152 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2719_
timestamp 18001
transform 1 0 17296 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2720_
timestamp 18001
transform 1 0 16652 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2721_
timestamp 18001
transform 1 0 19688 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2722_
timestamp 18001
transform 1 0 19228 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2723_
timestamp 18001
transform -1 0 23000 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2724_
timestamp 18001
transform 1 0 18032 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2725_
timestamp 18001
transform 1 0 19872 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2726_
timestamp 18001
transform 1 0 15548 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2727_
timestamp 18001
transform 1 0 17112 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2728_
timestamp 18001
transform 1 0 15272 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2729_
timestamp 18001
transform 1 0 13800 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2730_
timestamp 18001
transform 1 0 11776 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2731_
timestamp 18001
transform 1 0 10396 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2732_
timestamp 18001
transform 1 0 11960 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2733_
timestamp 18001
transform 1 0 11500 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2734_
timestamp 18001
transform 1 0 10672 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2735_
timestamp 18001
transform 1 0 13616 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2736_
timestamp 18001
transform 1 0 12972 0 -1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2737_
timestamp 18001
transform 1 0 13432 0 -1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2738_
timestamp 18001
transform 1 0 14996 0 1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2739_
timestamp 18001
transform -1 0 20148 0 -1 39168
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2740_
timestamp 18001
transform 1 0 19780 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2741_
timestamp 18001
transform 1 0 19596 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2742_
timestamp 18001
transform 1 0 19596 0 -1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2743_
timestamp 18001
transform 1 0 17664 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2744_
timestamp 18001
transform 1 0 12144 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2745_
timestamp 18001
transform 1 0 7268 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2746_
timestamp 18001
transform 1 0 3772 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2747_
timestamp 18001
transform 1 0 1564 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2748_
timestamp 18001
transform 1 0 3680 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2749_
timestamp 18001
transform 1 0 1564 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2750_
timestamp 18001
transform 1 0 1380 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2751_
timestamp 18001
transform -1 0 10764 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2752_
timestamp 18001
transform 1 0 10948 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2753_
timestamp 18001
transform 1 0 6808 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2754_
timestamp 18001
transform 1 0 3036 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2755_
timestamp 18001
transform 1 0 1472 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2756_
timestamp 18001
transform 1 0 3496 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2757_
timestamp 18001
transform 1 0 1840 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2758_
timestamp 18001
transform 1 0 1472 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2759_
timestamp 18001
transform 1 0 8556 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2760_
timestamp 18001
transform 1 0 22172 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2761_
timestamp 18001
transform 1 0 24748 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2762_
timestamp 18001
transform -1 0 28796 0 1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2763_
timestamp 18001
transform 1 0 22356 0 -1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2764_
timestamp 18001
transform 1 0 24564 0 1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2765_
timestamp 18001
transform 1 0 22632 0 -1 39168
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2766_
timestamp 18001
transform 1 0 23000 0 -1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2767_
timestamp 18001
transform 1 0 25116 0 1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2768_
timestamp 18001
transform 1 0 23552 0 -1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2769_
timestamp 18001
transform 1 0 14444 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2770_
timestamp 18001
transform 1 0 11960 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2771_
timestamp 18001
transform 1 0 6900 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2772_
timestamp 18001
transform 1 0 3864 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2773_
timestamp 18001
transform -1 0 5980 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2774_
timestamp 18001
transform 1 0 6348 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2775_
timestamp 18001
transform 1 0 8280 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2776_
timestamp 18001
transform 1 0 10304 0 1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2777_
timestamp 18001
transform 1 0 12512 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2778_
timestamp 18001
transform 1 0 6808 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2779_
timestamp 18001
transform 1 0 5520 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2780_
timestamp 18001
transform 1 0 2484 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2781_
timestamp 18001
transform 1 0 4416 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2782_
timestamp 18001
transform 1 0 3772 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2783_
timestamp 18001
transform 1 0 3772 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2784_
timestamp 18001
transform 1 0 6992 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2785_
timestamp 18001
transform -1 0 3956 0 -1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2786_
timestamp 18001
transform -1 0 5336 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2787_
timestamp 18001
transform -1 0 3680 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2788_
timestamp 18001
transform -1 0 3588 0 1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2789_
timestamp 18001
transform -1 0 4416 0 -1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2790_
timestamp 18001
transform 1 0 4140 0 -1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2791_
timestamp 18001
transform -1 0 3496 0 1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2792_
timestamp 18001
transform -1 0 4600 0 -1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2793_
timestamp 18001
transform -1 0 15548 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2794_
timestamp 18001
transform 1 0 2116 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2795_
timestamp 18001
transform 1 0 4784 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2796_
timestamp 18001
transform 1 0 3496 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2797_
timestamp 18001
transform 1 0 2944 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2798_
timestamp 18001
transform -1 0 6072 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2799_
timestamp 18001
transform 1 0 3956 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2800_
timestamp 18001
transform 1 0 9200 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2801_
timestamp 18001
transform 1 0 22448 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2802_
timestamp 18001
transform -1 0 26220 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2803_
timestamp 18001
transform 1 0 10856 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2804_
timestamp 18001
transform 1 0 6900 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2805_
timestamp 18001
transform 1 0 3772 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2806_
timestamp 18001
transform 1 0 1656 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2807_
timestamp 18001
transform 1 0 5152 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2808_
timestamp 18001
transform 1 0 2484 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2809_
timestamp 18001
transform 1 0 1564 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2810_
timestamp 18001
transform 1 0 8740 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2811_
timestamp 18001
transform 1 0 17204 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2812_
timestamp 18001
transform 1 0 29716 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2813_
timestamp 18001
transform 1 0 14628 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _2814_
timestamp 18001
transform -1 0 2116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 18001
transform -1 0 18308 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 18001
transform -1 0 23092 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 18001
transform -1 0 20332 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 18001
transform -1 0 39376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 18001
transform 1 0 20792 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk
timestamp 18001
transform 1 0 8924 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 18001
transform 1 0 6072 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 18001
transform -1 0 16560 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 18001
transform 1 0 14720 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 18001
transform 1 0 4324 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 18001
transform -1 0 4600 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 18001
transform 1 0 6348 0 -1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 18001
transform -1 0 8648 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 18001
transform -1 0 25484 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 18001
transform -1 0 24104 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 18001
transform 1 0 32476 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 18001
transform -1 0 32936 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 18001
transform 1 0 21804 0 -1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 18001
transform -1 0 23828 0 -1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 18001
transform 1 0 32844 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 18001
transform -1 0 31188 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_6  clkload0
timestamp 18001
transform 1 0 8188 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload1
timestamp 18001
transform -1 0 6992 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_8  clkload2
timestamp 18001
transform 1 0 15732 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_6  clkload3
timestamp 18001
transform 1 0 14076 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_4  clkload4
timestamp 18001
transform 1 0 2392 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__bufinv_16  clkload5
timestamp 18001
transform 1 0 5520 0 1 31552
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_4  clkload6
timestamp 18001
transform 1 0 8648 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__inv_6  clkload7
timestamp 18001
transform 1 0 24472 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  clkload8
timestamp 18001
transform 1 0 23092 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  clkload9
timestamp 18001
transform 1 0 32476 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__inv_6  clkload10
timestamp 18001
transform 1 0 31280 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload11
timestamp 18001
transform 1 0 21620 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload12
timestamp 18001
transform 1 0 22816 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_4  clkload13
timestamp 18001
transform 1 0 33672 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__inv_6  clkload14
timestamp 18001
transform 1 0 30176 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  fanout19
timestamp 18001
transform -1 0 11960 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout20
timestamp 18001
transform 1 0 18032 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout21
timestamp 18001
transform -1 0 38916 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout22
timestamp 18001
transform -1 0 12972 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout23
timestamp 18001
transform -1 0 9292 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout24
timestamp 18001
transform 1 0 11592 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout25
timestamp 18001
transform -1 0 23092 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  fanout26
timestamp 18001
transform -1 0 21528 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout27
timestamp 18001
transform -1 0 23092 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout28
timestamp 18001
transform 1 0 13156 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 18001
transform 1 0 39100 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout30
timestamp 18001
transform 1 0 10948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout31
timestamp 18001
transform -1 0 11040 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout32
timestamp 18001
transform -1 0 10856 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout33
timestamp 18001
transform 1 0 14076 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout34
timestamp 18001
transform -1 0 35788 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout35
timestamp 18001
transform -1 0 32752 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp 18001
transform -1 0 31924 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout37
timestamp 18001
transform 1 0 35696 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout38
timestamp 18001
transform -1 0 32568 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout39
timestamp 18001
transform -1 0 31004 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout40
timestamp 18001
transform 1 0 35512 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout41
timestamp 18001
transform 1 0 32292 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout42
timestamp 18001
transform 1 0 34224 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout43
timestamp 18001
transform 1 0 30636 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout44
timestamp 18001
transform 1 0 30728 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout45
timestamp 18001
transform -1 0 14720 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout46
timestamp 18001
transform -1 0 19596 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout47
timestamp 18001
transform -1 0 19964 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout48
timestamp 18001
transform -1 0 15732 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout49
timestamp 18001
transform 1 0 24932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout50
timestamp 18001
transform -1 0 24104 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout51
timestamp 18001
transform -1 0 32568 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout52
timestamp 18001
transform 1 0 25760 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout53
timestamp 18001
transform -1 0 21252 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout54
timestamp 18001
transform -1 0 29992 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout55
timestamp 18001
transform -1 0 24748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout56
timestamp 18001
transform 1 0 24748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout57
timestamp 18001
transform 1 0 20792 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout58
timestamp 18001
transform 1 0 20884 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout59
timestamp 18001
transform -1 0 17204 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout60
timestamp 18001
transform -1 0 21528 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout61
timestamp 18001
transform 1 0 33672 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout62
timestamp 18001
transform 1 0 34040 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout63
timestamp 18001
transform 1 0 35788 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout64
timestamp 18001
transform 1 0 31740 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout65
timestamp 18001
transform 1 0 31096 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout66
timestamp 18001
transform 1 0 31740 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout67
timestamp 18001
transform -1 0 25760 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout68
timestamp 18001
transform -1 0 30820 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout69
timestamp 18001
transform -1 0 32016 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout70
timestamp 18001
transform 1 0 22172 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout71
timestamp 18001
transform -1 0 27324 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout72
timestamp 18001
transform -1 0 27692 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout73
timestamp 18001
transform 1 0 24380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout74
timestamp 18001
transform -1 0 23368 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout75
timestamp 18001
transform 1 0 33488 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout76
timestamp 18001
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout77
timestamp 18001
transform -1 0 24288 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout78
timestamp 18001
transform 1 0 34868 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout79
timestamp 18001
transform -1 0 32016 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout80
timestamp 18001
transform 1 0 33488 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout81
timestamp 18001
transform 1 0 33856 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout82
timestamp 18001
transform -1 0 32016 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout83
timestamp 18001
transform -1 0 29348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout84
timestamp 18001
transform -1 0 29900 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout85
timestamp 18001
transform 1 0 37720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout86
timestamp 18001
transform -1 0 30912 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout87
timestamp 18001
transform -1 0 24288 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout88
timestamp 18001
transform 1 0 24104 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout89
timestamp 18001
transform -1 0 35788 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout90
timestamp 18001
transform 1 0 34960 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout91
timestamp 18001
transform 1 0 35512 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout92
timestamp 18001
transform -1 0 29440 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout93
timestamp 18001
transform -1 0 32660 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout94
timestamp 18001
transform -1 0 37904 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout95
timestamp 18001
transform -1 0 28888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout96
timestamp 18001
transform -1 0 32384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout97
timestamp 18001
transform 1 0 36340 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout98
timestamp 18001
transform 1 0 27692 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout99
timestamp 18001
transform -1 0 31188 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout100
timestamp 18001
transform -1 0 38640 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout101
timestamp 18001
transform 1 0 37904 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout102
timestamp 18001
transform -1 0 29716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout103
timestamp 18001
transform -1 0 38824 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout104
timestamp 18001
transform -1 0 38456 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout105
timestamp 18001
transform 1 0 28520 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout106
timestamp 18001
transform 1 0 28520 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout107
timestamp 18001
transform -1 0 26864 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout108
timestamp 18001
transform 1 0 30176 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout109
timestamp 18001
transform -1 0 28980 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout110
timestamp 18001
transform 1 0 29440 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout111
timestamp 18001
transform 1 0 28704 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout112
timestamp 18001
transform 1 0 29532 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  fanout113
timestamp 18001
transform -1 0 29072 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  fanout114
timestamp 18001
transform -1 0 28520 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout115
timestamp 18001
transform 1 0 28796 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout116
timestamp 18001
transform -1 0 28152 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout117
timestamp 18001
transform 1 0 20608 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout118
timestamp 18001
transform -1 0 23552 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout119
timestamp 18001
transform 1 0 23828 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout120
timestamp 18001
transform -1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout121
timestamp 18001
transform -1 0 29440 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout122
timestamp 18001
transform 1 0 29808 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout123
timestamp 18001
transform -1 0 21712 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout124
timestamp 18001
transform -1 0 24564 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout125
timestamp 18001
transform -1 0 31372 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout126
timestamp 18001
transform -1 0 29164 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout127
timestamp 18001
transform 1 0 30360 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout128
timestamp 18001
transform 1 0 28336 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout129
timestamp 18001
transform -1 0 4324 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout130
timestamp 18001
transform -1 0 13892 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout131
timestamp 18001
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout132
timestamp 18001
transform 1 0 20148 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout133
timestamp 18001
transform 1 0 20700 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout134
timestamp 18001
transform -1 0 4692 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout135
timestamp 18001
transform 1 0 9660 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout136
timestamp 18001
transform -1 0 4968 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout137
timestamp 18001
transform -1 0 8648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout138
timestamp 18001
transform 1 0 21160 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout139
timestamp 18001
transform -1 0 13984 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout140
timestamp 18001
transform 1 0 20332 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout141
timestamp 18001
transform 1 0 30084 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout142
timestamp 18001
transform -1 0 40204 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout143
timestamp 18001
transform -1 0 30820 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout144
timestamp 18001
transform -1 0 39744 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout145
timestamp 18001
transform -1 0 40296 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout146
timestamp 18001
transform -1 0 38548 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout147
timestamp 18001
transform -1 0 38916 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout148
timestamp 18001
transform -1 0 38088 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636986456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636986456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 18001
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636986456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1636986456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 18001
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636986456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1636986456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 18001
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1636986456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_97
timestamp 18001
transform 1 0 10028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_105
timestamp 18001
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 18001
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_141
timestamp 18001
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_147
timestamp 18001
transform 1 0 14628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_158
timestamp 18001
transform 1 0 15640 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_169
timestamp 18001
transform 1 0 16652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_194
timestamp 18001
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_200
timestamp 18001
transform 1 0 19504 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_204
timestamp 18001
transform 1 0 19872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_213
timestamp 18001
transform 1 0 20700 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1636986456
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_237
timestamp 18001
transform 1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_246
timestamp 18001
transform 1 0 23736 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1636986456
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1636986456
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 18001
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1636986456
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1636986456
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 18001
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1636986456
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1636986456
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 18001
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1636986456
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1636986456
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 18001
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 1636986456
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_377
timestamp 1636986456
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 18001
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_393
timestamp 1636986456
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_405
timestamp 1636986456
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_417
timestamp 18001
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_421
timestamp 18001
transform 1 0 39836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_425
timestamp 18001
transform 1 0 40204 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636986456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636986456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636986456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1636986456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 18001
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 18001
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1636986456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1636986456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1636986456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1636986456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 18001
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 18001
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_113
timestamp 18001
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 18001
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 18001
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_178
timestamp 18001
transform 1 0 17480 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_247
timestamp 18001
transform 1 0 23828 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_269
timestamp 18001
transform 1 0 25852 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_277
timestamp 18001
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1636986456
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1636986456
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1636986456
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1636986456
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 18001
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 18001
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1636986456
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1636986456
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1636986456
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1636986456
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 18001
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 18001
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 1636986456
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_405
timestamp 1636986456
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_417
timestamp 18001
transform 1 0 39468 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_425
timestamp 18001
transform 1 0 40204 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636986456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636986456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 18001
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1636986456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1636986456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1636986456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1636986456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 18001
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 18001
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1636986456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_97
timestamp 18001
transform 1 0 10028 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_103
timestamp 18001
transform 1 0 10580 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 18001
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_141
timestamp 18001
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_153
timestamp 18001
transform 1 0 15180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_185
timestamp 18001
transform 1 0 18124 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_193
timestamp 18001
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_205
timestamp 1636986456
transform 1 0 19964 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_217
timestamp 18001
transform 1 0 21068 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_231
timestamp 18001
transform 1 0 22356 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_281
timestamp 1636986456
transform 1 0 26956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_293
timestamp 1636986456
transform 1 0 28060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_305
timestamp 18001
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1636986456
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1636986456
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1636986456
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1636986456
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 18001
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 18001
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1636986456
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1636986456
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1636986456
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 1636986456
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 18001
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 18001
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_421
timestamp 18001
transform 1 0 39836 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636986456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636986456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1636986456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1636986456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 18001
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 18001
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1636986456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1636986456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1636986456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1636986456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 18001
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 18001
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_131
timestamp 18001
transform 1 0 13156 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_149
timestamp 18001
transform 1 0 14812 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_161
timestamp 18001
transform 1 0 15916 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_172
timestamp 18001
transform 1 0 16928 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_182
timestamp 18001
transform 1 0 17848 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_186
timestamp 18001
transform 1 0 18216 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_213
timestamp 18001
transform 1 0 20700 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_225
timestamp 18001
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_235
timestamp 18001
transform 1 0 22724 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_244
timestamp 1636986456
transform 1 0 23552 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_256
timestamp 1636986456
transform 1 0 24656 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_268
timestamp 1636986456
transform 1 0 25760 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1636986456
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_293
timestamp 18001
transform 1 0 28060 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_315
timestamp 1636986456
transform 1 0 30084 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_327
timestamp 18001
transform 1 0 31188 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 18001
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1636986456
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1636986456
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1636986456
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1636986456
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 18001
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 18001
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1636986456
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1636986456
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_417
timestamp 18001
transform 1 0 39468 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_425
timestamp 18001
transform 1 0 40204 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1636986456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1636986456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 18001
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1636986456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1636986456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1636986456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1636986456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 18001
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 18001
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1636986456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1636986456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_109
timestamp 18001
transform 1 0 11132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_113
timestamp 18001
transform 1 0 11500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 18001
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_141
timestamp 18001
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_152
timestamp 18001
transform 1 0 15088 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_174
timestamp 18001
transform 1 0 17112 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_238
timestamp 1636986456
transform 1 0 23000 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_250
timestamp 18001
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_253
timestamp 18001
transform 1 0 24380 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_280
timestamp 1636986456
transform 1 0 26864 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_292
timestamp 1636986456
transform 1 0 27968 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_304
timestamp 18001
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1636986456
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1636986456
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1636986456
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1636986456
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 18001
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 18001
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1636986456
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1636986456
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1636986456
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1636986456
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 18001
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 18001
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_421
timestamp 18001
transform 1 0 39836 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_425
timestamp 18001
transform 1 0 40204 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1636986456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1636986456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1636986456
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1636986456
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 18001
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 18001
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1636986456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1636986456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1636986456
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1636986456
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 18001
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 18001
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_113
timestamp 18001
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_164
timestamp 18001
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_196
timestamp 18001
transform 1 0 19136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_206
timestamp 18001
transform 1 0 20056 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_217
timestamp 18001
transform 1 0 21068 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_245
timestamp 18001
transform 1 0 23644 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_253
timestamp 18001
transform 1 0 24380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 18001
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_306
timestamp 18001
transform 1 0 29256 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_314
timestamp 18001
transform 1 0 29992 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_321
timestamp 1636986456
transform 1 0 30636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_333
timestamp 18001
transform 1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1636986456
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1636986456
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1636986456
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1636986456
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 18001
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 18001
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1636986456
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1636986456
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_417
timestamp 18001
transform 1 0 39468 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_425
timestamp 18001
transform 1 0 40204 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1636986456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1636986456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 18001
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1636986456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1636986456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1636986456
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1636986456
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 18001
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 18001
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1636986456
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_97
timestamp 18001
transform 1 0 10028 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1636986456
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 18001
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 18001
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1636986456
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1636986456
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_165
timestamp 18001
transform 1 0 16284 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_182
timestamp 18001
transform 1 0 17848 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_191
timestamp 18001
transform 1 0 18676 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_197
timestamp 18001
transform 1 0 19228 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_207
timestamp 18001
transform 1 0 20148 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_214
timestamp 18001
transform 1 0 20792 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_226
timestamp 18001
transform 1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_253
timestamp 18001
transform 1 0 24380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_272
timestamp 18001
transform 1 0 26128 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_280
timestamp 18001
transform 1 0 26864 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_329
timestamp 1636986456
transform 1 0 31372 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_341
timestamp 1636986456
transform 1 0 32476 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_353
timestamp 18001
transform 1 0 33580 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_361
timestamp 18001
transform 1 0 34316 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1636986456
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1636986456
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1636986456
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1636986456
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 18001
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 18001
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_421
timestamp 18001
transform 1 0 39836 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_425
timestamp 18001
transform 1 0 40204 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1636986456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1636986456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1636986456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1636986456
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 18001
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 18001
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1636986456
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1636986456
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1636986456
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1636986456
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 18001
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 18001
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_130
timestamp 1636986456
transform 1 0 13064 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_142
timestamp 18001
transform 1 0 14168 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_146
timestamp 18001
transform 1 0 14536 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1636986456
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_222
timestamp 18001
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_225
timestamp 18001
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_229
timestamp 18001
transform 1 0 22172 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1636986456
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_249
timestamp 18001
transform 1 0 24012 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_257
timestamp 18001
transform 1 0 24748 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_263
timestamp 1636986456
transform 1 0 25300 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_275
timestamp 18001
transform 1 0 26404 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_294
timestamp 1636986456
transform 1 0 28152 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_306
timestamp 18001
transform 1 0 29256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_328
timestamp 18001
transform 1 0 31280 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1636986456
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1636986456
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1636986456
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1636986456
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 18001
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 18001
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1636986456
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1636986456
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_417
timestamp 18001
transform 1 0 39468 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_425
timestamp 18001
transform 1 0 40204 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1636986456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1636986456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 18001
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1636986456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1636986456
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1636986456
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1636986456
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 18001
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 18001
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1636986456
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1636986456
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_109
timestamp 18001
transform 1 0 11132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_125
timestamp 18001
transform 1 0 12604 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_131
timestamp 18001
transform 1 0 13156 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 18001
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_151
timestamp 18001
transform 1 0 14996 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_155
timestamp 18001
transform 1 0 15364 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_179
timestamp 1636986456
transform 1 0 17572 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_191
timestamp 18001
transform 1 0 18676 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 18001
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1636986456
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_209
timestamp 18001
transform 1 0 20332 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_213
timestamp 18001
transform 1 0 20700 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_220
timestamp 1636986456
transform 1 0 21344 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_232
timestamp 1636986456
transform 1 0 22448 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_244
timestamp 18001
transform 1 0 23552 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1636986456
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1636986456
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1636986456
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1636986456
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 18001
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 18001
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_320
timestamp 1636986456
transform 1 0 30544 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_332
timestamp 1636986456
transform 1 0 31648 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_344
timestamp 18001
transform 1 0 32752 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_352
timestamp 18001
transform 1 0 33488 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_361
timestamp 18001
transform 1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1636986456
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_377
timestamp 18001
transform 1 0 35788 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_403
timestamp 1636986456
transform 1 0 38180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_415
timestamp 18001
transform 1 0 39284 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 18001
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_421
timestamp 18001
transform 1 0 39836 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_425
timestamp 18001
transform 1 0 40204 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1636986456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1636986456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1636986456
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1636986456
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 18001
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 18001
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1636986456
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_69
timestamp 18001
transform 1 0 7452 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_80
timestamp 18001
transform 1 0 8464 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_108
timestamp 18001
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_113
timestamp 18001
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_117
timestamp 18001
transform 1 0 11868 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_121
timestamp 18001
transform 1 0 12236 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_156
timestamp 18001
transform 1 0 15456 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_179
timestamp 18001
transform 1 0 17572 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1636986456
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_205
timestamp 18001
transform 1 0 19964 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_211
timestamp 18001
transform 1 0 20516 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_225
timestamp 18001
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_232
timestamp 1636986456
transform 1 0 22448 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_244
timestamp 18001
transform 1 0 23552 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_252
timestamp 18001
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_267
timestamp 18001
transform 1 0 25668 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1636986456
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_305
timestamp 18001
transform 1 0 29164 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_312
timestamp 18001
transform 1 0 29808 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_320
timestamp 18001
transform 1 0 30544 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_332
timestamp 18001
transform 1 0 31648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_345
timestamp 18001
transform 1 0 32844 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_353
timestamp 18001
transform 1 0 33580 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_364
timestamp 18001
transform 1 0 34592 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_379
timestamp 1636986456
transform 1 0 35972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 18001
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_396
timestamp 18001
transform 1 0 37536 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_424
timestamp 18001
transform 1 0 40112 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1636986456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1636986456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 18001
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1636986456
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_41
timestamp 18001
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_53
timestamp 18001
transform 1 0 5980 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_66
timestamp 18001
transform 1 0 7176 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_81
timestamp 18001
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_85
timestamp 18001
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_98
timestamp 18001
transform 1 0 10120 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_104
timestamp 18001
transform 1 0 10672 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_111
timestamp 1636986456
transform 1 0 11316 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_123
timestamp 1636986456
transform 1 0 12420 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_135
timestamp 18001
transform 1 0 13524 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_147
timestamp 18001
transform 1 0 14628 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_185
timestamp 18001
transform 1 0 18124 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_194
timestamp 18001
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_200
timestamp 18001
transform 1 0 19504 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_204
timestamp 18001
transform 1 0 19872 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_212
timestamp 18001
transform 1 0 20608 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_234
timestamp 18001
transform 1 0 22632 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_243
timestamp 18001
transform 1 0 23460 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_253
timestamp 18001
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_275
timestamp 18001
transform 1 0 26404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_285
timestamp 18001
transform 1 0 27324 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_309
timestamp 18001
transform 1 0 29532 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_339
timestamp 18001
transform 1 0 32292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_360
timestamp 18001
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_378
timestamp 18001
transform 1 0 35880 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_382
timestamp 18001
transform 1 0 36248 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_410
timestamp 18001
transform 1 0 38824 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_418
timestamp 18001
transform 1 0 39560 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_425
timestamp 18001
transform 1 0 40204 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1636986456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1636986456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_27
timestamp 18001
transform 1 0 3588 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_33
timestamp 18001
transform 1 0 4140 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 18001
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_57
timestamp 18001
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_65
timestamp 18001
transform 1 0 7084 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_87
timestamp 1636986456
transform 1 0 9108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_99
timestamp 18001
transform 1 0 10212 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_110
timestamp 18001
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_126
timestamp 18001
transform 1 0 12696 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 18001
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 18001
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_169
timestamp 18001
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_184
timestamp 18001
transform 1 0 18032 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_196
timestamp 18001
transform 1 0 19136 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_215
timestamp 18001
transform 1 0 20884 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_222
timestamp 18001
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_230
timestamp 18001
transform 1 0 22264 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_254
timestamp 18001
transform 1 0 24472 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 18001
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_322
timestamp 1636986456
transform 1 0 30728 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_334
timestamp 18001
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_343
timestamp 18001
transform 1 0 32660 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_349
timestamp 18001
transform 1 0 33212 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_356
timestamp 18001
transform 1 0 33856 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_368
timestamp 18001
transform 1 0 34960 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_376
timestamp 18001
transform 1 0 35696 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_388
timestamp 18001
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_393
timestamp 18001
transform 1 0 37260 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_397
timestamp 18001
transform 1 0 37628 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_402
timestamp 18001
transform 1 0 38088 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1636986456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1636986456
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 18001
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1636986456
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1636986456
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_53
timestamp 18001
transform 1 0 5980 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_61
timestamp 18001
transform 1 0 6716 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_70
timestamp 18001
transform 1 0 7544 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_75
timestamp 18001
transform 1 0 8004 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_80
timestamp 18001
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1636986456
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_97
timestamp 18001
transform 1 0 10028 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_128
timestamp 1636986456
transform 1 0 12880 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_159
timestamp 1636986456
transform 1 0 15732 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_171
timestamp 18001
transform 1 0 16836 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_184
timestamp 1636986456
transform 1 0 18032 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1636986456
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_219
timestamp 18001
transform 1 0 21252 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_227
timestamp 18001
transform 1 0 21988 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_235
timestamp 1636986456
transform 1 0 22724 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_247
timestamp 18001
transform 1 0 23828 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_268
timestamp 18001
transform 1 0 25760 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_286
timestamp 18001
transform 1 0 27416 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_291
timestamp 18001
transform 1 0 27876 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_313
timestamp 18001
transform 1 0 29900 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_324
timestamp 18001
transform 1 0 30912 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_331
timestamp 1636986456
transform 1 0 31556 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_343
timestamp 18001
transform 1 0 32660 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_354
timestamp 18001
transform 1 0 33672 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_362
timestamp 18001
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_365
timestamp 18001
transform 1 0 34684 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1636986456
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_389
timestamp 18001
transform 1 0 36892 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_408
timestamp 1636986456
transform 1 0 38640 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_421
timestamp 18001
transform 1 0 39836 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_425
timestamp 18001
transform 1 0 40204 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1636986456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1636986456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1636986456
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1636986456
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 18001
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 18001
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_69
timestamp 18001
transform 1 0 7452 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_75
timestamp 18001
transform 1 0 8004 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_82
timestamp 18001
transform 1 0 8648 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_95
timestamp 18001
transform 1 0 9844 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_103
timestamp 18001
transform 1 0 10580 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_119
timestamp 18001
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_136
timestamp 18001
transform 1 0 13616 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_142
timestamp 18001
transform 1 0 14168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_151
timestamp 18001
transform 1 0 14996 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_159
timestamp 18001
transform 1 0 15732 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_165
timestamp 18001
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1636986456
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_181
timestamp 18001
transform 1 0 17756 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_189
timestamp 1636986456
transform 1 0 18492 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_201
timestamp 18001
transform 1 0 19596 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_209
timestamp 18001
transform 1 0 20332 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 18001
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 18001
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_225
timestamp 18001
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_239
timestamp 18001
transform 1 0 23092 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_247
timestamp 18001
transform 1 0 23828 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_254
timestamp 18001
transform 1 0 24472 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_258
timestamp 18001
transform 1 0 24840 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_264
timestamp 1636986456
transform 1 0 25392 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_276
timestamp 18001
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_293
timestamp 18001
transform 1 0 28060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_297
timestamp 18001
transform 1 0 28428 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_302
timestamp 18001
transform 1 0 28888 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_307
timestamp 18001
transform 1 0 29348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_311
timestamp 18001
transform 1 0 29716 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_330
timestamp 18001
transform 1 0 31464 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_347
timestamp 1636986456
transform 1 0 33028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_359
timestamp 18001
transform 1 0 34132 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_368
timestamp 18001
transform 1 0 34960 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 18001
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_393
timestamp 18001
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_410
timestamp 1636986456
transform 1 0 38824 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_422
timestamp 18001
transform 1 0 39928 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1636986456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1636986456
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 18001
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_29
timestamp 18001
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_51
timestamp 18001
transform 1 0 5796 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_74
timestamp 18001
transform 1 0 7912 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_100
timestamp 18001
transform 1 0 10304 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_108
timestamp 18001
transform 1 0 11040 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_114
timestamp 18001
transform 1 0 11592 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_120
timestamp 18001
transform 1 0 12144 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_129
timestamp 18001
transform 1 0 12972 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_137
timestamp 18001
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_141
timestamp 18001
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_151
timestamp 18001
transform 1 0 14996 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_184
timestamp 18001
transform 1 0 18032 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_208
timestamp 1636986456
transform 1 0 20240 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_220
timestamp 1636986456
transform 1 0 21344 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_232
timestamp 1636986456
transform 1 0 22448 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_244
timestamp 18001
transform 1 0 23552 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_253
timestamp 18001
transform 1 0 24380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_279
timestamp 18001
transform 1 0 26772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_287
timestamp 18001
transform 1 0 27508 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_309
timestamp 18001
transform 1 0 29532 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_315
timestamp 18001
transform 1 0 30084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_327
timestamp 18001
transform 1 0 31188 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_335
timestamp 18001
transform 1 0 31924 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_347
timestamp 1636986456
transform 1 0 33028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_359
timestamp 18001
transform 1 0 34132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 18001
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_365
timestamp 18001
transform 1 0 34684 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_373
timestamp 18001
transform 1 0 35420 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_378
timestamp 18001
transform 1 0 35880 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_386
timestamp 18001
transform 1 0 36616 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_393
timestamp 18001
transform 1 0 37260 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_421
timestamp 18001
transform 1 0 39836 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_425
timestamp 18001
transform 1 0 40204 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1636986456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1636986456
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1636986456
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1636986456
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 18001
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 18001
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_78
timestamp 18001
transform 1 0 8280 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_88
timestamp 18001
transform 1 0 9200 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_100
timestamp 1636986456
transform 1 0 10304 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_113
timestamp 18001
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_121
timestamp 18001
transform 1 0 12236 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_130
timestamp 1636986456
transform 1 0 13064 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_142
timestamp 18001
transform 1 0 14168 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_153
timestamp 1636986456
transform 1 0 15180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_165
timestamp 18001
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_169
timestamp 18001
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_175
timestamp 1636986456
transform 1 0 17204 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_187
timestamp 1636986456
transform 1 0 18308 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_199
timestamp 1636986456
transform 1 0 19412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_211
timestamp 18001
transform 1 0 20516 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_215
timestamp 18001
transform 1 0 20884 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_234
timestamp 18001
transform 1 0 22632 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_244
timestamp 18001
transform 1 0 23552 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_265
timestamp 18001
transform 1 0 25484 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_274
timestamp 18001
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_281
timestamp 18001
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_297
timestamp 1636986456
transform 1 0 28428 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_309
timestamp 18001
transform 1 0 29532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_319
timestamp 18001
transform 1 0 30452 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_352
timestamp 1636986456
transform 1 0 33488 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_364
timestamp 1636986456
transform 1 0 34592 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_376
timestamp 1636986456
transform 1 0 35696 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_388
timestamp 18001
transform 1 0 36800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_399
timestamp 18001
transform 1 0 37812 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_403
timestamp 18001
transform 1 0 38180 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_409
timestamp 18001
transform 1 0 38732 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_415
timestamp 18001
transform 1 0 39284 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_423
timestamp 18001
transform 1 0 40020 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_3
timestamp 18001
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_11
timestamp 1636986456
transform 1 0 2116 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_23
timestamp 18001
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 18001
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1636986456
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1636986456
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1636986456
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_65
timestamp 18001
transform 1 0 7084 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_88
timestamp 18001
transform 1 0 9200 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_110
timestamp 18001
transform 1 0 11224 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_119
timestamp 18001
transform 1 0 12052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_132
timestamp 18001
transform 1 0 13248 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_144
timestamp 18001
transform 1 0 14352 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_152
timestamp 18001
transform 1 0 15088 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_159
timestamp 1636986456
transform 1 0 15732 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_171
timestamp 18001
transform 1 0 16836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_190
timestamp 18001
transform 1 0 18584 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_197
timestamp 18001
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_201
timestamp 18001
transform 1 0 19596 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_207
timestamp 18001
transform 1 0 20148 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_214
timestamp 18001
transform 1 0 20792 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_218
timestamp 18001
transform 1 0 21160 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_227
timestamp 18001
transform 1 0 21988 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_238
timestamp 18001
transform 1 0 23000 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_248
timestamp 18001
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_258
timestamp 18001
transform 1 0 24840 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_266
timestamp 18001
transform 1 0 25576 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_274
timestamp 18001
transform 1 0 26312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_278
timestamp 18001
transform 1 0 26680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_283
timestamp 18001
transform 1 0 27140 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_296
timestamp 18001
transform 1 0 28336 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_301
timestamp 18001
transform 1 0 28796 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_323
timestamp 18001
transform 1 0 30820 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_327
timestamp 18001
transform 1 0 31188 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_353
timestamp 18001
transform 1 0 33580 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_362
timestamp 18001
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_372
timestamp 18001
transform 1 0 35328 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_380
timestamp 18001
transform 1 0 36064 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_396
timestamp 1636986456
transform 1 0 37536 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_408
timestamp 1636986456
transform 1 0 38640 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_421
timestamp 18001
transform 1 0 39836 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_425
timestamp 18001
transform 1 0 40204 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1636986456
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_15
timestamp 18001
transform 1 0 2484 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_23
timestamp 18001
transform 1 0 3220 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_46
timestamp 18001
transform 1 0 5336 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 18001
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_62
timestamp 1636986456
transform 1 0 6808 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_74
timestamp 18001
transform 1 0 7912 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_88
timestamp 18001
transform 1 0 9200 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_102
timestamp 18001
transform 1 0 10488 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_110
timestamp 18001
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1636986456
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_125
timestamp 18001
transform 1 0 12604 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_135
timestamp 18001
transform 1 0 13524 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_162
timestamp 18001
transform 1 0 16008 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_169
timestamp 18001
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_177
timestamp 1636986456
transform 1 0 17388 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_189
timestamp 1636986456
transform 1 0 18492 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_201
timestamp 18001
transform 1 0 19596 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_218
timestamp 18001
transform 1 0 21160 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1636986456
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_237
timestamp 18001
transform 1 0 22908 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_273
timestamp 18001
transform 1 0 26220 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 18001
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1636986456
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_293
timestamp 18001
transform 1 0 28060 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_300
timestamp 1636986456
transform 1 0 28704 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_312
timestamp 1636986456
transform 1 0 29808 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_324
timestamp 18001
transform 1 0 30912 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_337
timestamp 18001
transform 1 0 32108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_358
timestamp 18001
transform 1 0 34040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_362
timestamp 18001
transform 1 0 34408 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_371
timestamp 1636986456
transform 1 0 35236 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_383
timestamp 18001
transform 1 0 36340 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_393
timestamp 18001
transform 1 0 37260 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_413
timestamp 1636986456
transform 1 0 39100 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_425
timestamp 18001
transform 1 0 40204 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1636986456
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1636986456
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 18001
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_41
timestamp 18001
transform 1 0 4876 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_73
timestamp 18001
transform 1 0 7820 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_81
timestamp 18001
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1636986456
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1636986456
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1636986456
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_121
timestamp 18001
transform 1 0 12236 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_132
timestamp 18001
transform 1 0 13248 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_156
timestamp 1636986456
transform 1 0 15456 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_168
timestamp 18001
transform 1 0 16560 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_188
timestamp 18001
transform 1 0 18400 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 18001
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_216
timestamp 1636986456
transform 1 0 20976 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_228
timestamp 1636986456
transform 1 0 22080 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_240
timestamp 1636986456
transform 1 0 23184 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1636986456
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_265
timestamp 18001
transform 1 0 25484 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_274
timestamp 1636986456
transform 1 0 26312 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_286
timestamp 18001
transform 1 0 27416 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_295
timestamp 1636986456
transform 1 0 28244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 18001
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_309
timestamp 18001
transform 1 0 29532 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_316
timestamp 18001
transform 1 0 30176 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_324
timestamp 1636986456
transform 1 0 30912 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_336
timestamp 18001
transform 1 0 32016 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_340
timestamp 18001
transform 1 0 32384 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_350
timestamp 18001
transform 1 0 33304 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_356
timestamp 18001
transform 1 0 33856 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_377
timestamp 1636986456
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_389
timestamp 1636986456
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_401
timestamp 18001
transform 1 0 37996 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_408
timestamp 1636986456
transform 1 0 38640 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_421
timestamp 18001
transform 1 0 39836 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_425
timestamp 18001
transform 1 0 40204 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_3
timestamp 18001
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_31
timestamp 18001
transform 1 0 3956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_40
timestamp 18001
transform 1 0 4784 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 18001
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_57
timestamp 18001
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_82
timestamp 1636986456
transform 1 0 8648 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_94
timestamp 18001
transform 1 0 9752 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_102
timestamp 18001
transform 1 0 10488 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 18001
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_119
timestamp 18001
transform 1 0 12052 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_123
timestamp 18001
transform 1 0 12420 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_133
timestamp 18001
transform 1 0 13340 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 1636986456
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 18001
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 18001
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_185
timestamp 18001
transform 1 0 18124 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_195
timestamp 1636986456
transform 1 0 19044 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_207
timestamp 18001
transform 1 0 20148 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_215
timestamp 18001
transform 1 0 20884 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 18001
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_267
timestamp 1636986456
transform 1 0 25668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 18001
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_289
timestamp 18001
transform 1 0 27692 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_306
timestamp 18001
transform 1 0 29256 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_310
timestamp 18001
transform 1 0 29624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 18001
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 18001
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_344
timestamp 1636986456
transform 1 0 32752 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_356
timestamp 18001
transform 1 0 33856 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_364
timestamp 18001
transform 1 0 34592 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_374
timestamp 1636986456
transform 1 0 35512 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_386
timestamp 18001
transform 1 0 36616 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_393
timestamp 1636986456
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_405
timestamp 18001
transform 1 0 38364 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_414
timestamp 1636986456
transform 1 0 39192 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1636986456
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_15
timestamp 18001
transform 1 0 2484 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_23
timestamp 18001
transform 1 0 3220 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_48
timestamp 1636986456
transform 1 0 5520 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_60
timestamp 18001
transform 1 0 6624 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_81
timestamp 18001
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_85
timestamp 18001
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_126
timestamp 18001
transform 1 0 12696 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_136
timestamp 18001
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_156
timestamp 18001
transform 1 0 15456 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_160
timestamp 18001
transform 1 0 15824 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_185
timestamp 18001
transform 1 0 18124 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_193
timestamp 18001
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_210
timestamp 18001
transform 1 0 20424 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_214
timestamp 18001
transform 1 0 20792 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_223
timestamp 18001
transform 1 0 21620 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_227
timestamp 18001
transform 1 0 21988 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_241
timestamp 18001
transform 1 0 23276 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_249
timestamp 18001
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1636986456
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_265
timestamp 18001
transform 1 0 25484 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_286
timestamp 1636986456
transform 1 0 27416 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_298
timestamp 18001
transform 1 0 28520 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_306
timestamp 18001
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_309
timestamp 18001
transform 1 0 29532 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_318
timestamp 1636986456
transform 1 0 30360 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_330
timestamp 18001
transform 1 0 31464 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_352
timestamp 1636986456
transform 1 0 33488 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_371
timestamp 1636986456
transform 1 0 35236 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_383
timestamp 1636986456
transform 1 0 36340 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_395
timestamp 1636986456
transform 1 0 37444 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_418
timestamp 18001
transform 1 0 39560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_421
timestamp 18001
transform 1 0 39836 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_425
timestamp 18001
transform 1 0 40204 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1636986456
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1636986456
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_27
timestamp 18001
transform 1 0 3588 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_40
timestamp 1636986456
transform 1 0 4784 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_52
timestamp 18001
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1636986456
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1636986456
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_81
timestamp 18001
transform 1 0 8556 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_87
timestamp 18001
transform 1 0 9108 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_94
timestamp 18001
transform 1 0 9752 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_98
timestamp 18001
transform 1 0 10120 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_107
timestamp 18001
transform 1 0 10948 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 18001
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_113
timestamp 18001
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_119
timestamp 18001
transform 1 0 12052 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_142
timestamp 1636986456
transform 1 0 14168 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_154
timestamp 18001
transform 1 0 15272 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 18001
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1636986456
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 1636986456
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_193
timestamp 18001
transform 1 0 18860 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_204
timestamp 1636986456
transform 1 0 19872 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_216
timestamp 18001
transform 1 0 20976 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1636986456
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_237
timestamp 18001
transform 1 0 22908 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_257
timestamp 18001
transform 1 0 24748 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_265
timestamp 18001
transform 1 0 25484 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_270
timestamp 18001
transform 1 0 25944 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_284
timestamp 18001
transform 1 0 27232 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_298
timestamp 18001
transform 1 0 28520 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_303
timestamp 1636986456
transform 1 0 28980 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_315
timestamp 18001
transform 1 0 30084 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_324
timestamp 1636986456
transform 1 0 30912 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_337
timestamp 18001
transform 1 0 32108 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_341
timestamp 18001
transform 1 0 32476 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_348
timestamp 1636986456
transform 1 0 33120 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_360
timestamp 1636986456
transform 1 0 34224 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_372
timestamp 1636986456
transform 1 0 35328 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_384
timestamp 18001
transform 1 0 36432 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_399
timestamp 18001
transform 1 0 37812 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_411
timestamp 1636986456
transform 1 0 38916 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_423
timestamp 18001
transform 1 0 40020 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1636986456
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1636986456
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 18001
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_29
timestamp 18001
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_43
timestamp 18001
transform 1 0 5060 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_51
timestamp 18001
transform 1 0 5796 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_63
timestamp 18001
transform 1 0 6900 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_74
timestamp 18001
transform 1 0 7912 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_85
timestamp 18001
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_103
timestamp 1636986456
transform 1 0 10580 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_115
timestamp 18001
transform 1 0 11684 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_123
timestamp 18001
transform 1 0 12420 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_127
timestamp 1636986456
transform 1 0 12788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 18001
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_141
timestamp 18001
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_152
timestamp 18001
transform 1 0 15088 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_167
timestamp 18001
transform 1 0 16468 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_171
timestamp 18001
transform 1 0 16836 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_178
timestamp 18001
transform 1 0 17480 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_186
timestamp 18001
transform 1 0 18216 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_197
timestamp 18001
transform 1 0 19228 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_219
timestamp 18001
transform 1 0 21252 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_242
timestamp 18001
transform 1 0 23368 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_250
timestamp 18001
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_253
timestamp 18001
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_259
timestamp 18001
transform 1 0 24932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_263
timestamp 18001
transform 1 0 25300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_272
timestamp 18001
transform 1 0 26128 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_279
timestamp 1636986456
transform 1 0 26772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_305
timestamp 18001
transform 1 0 29164 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_309
timestamp 18001
transform 1 0 29532 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_321
timestamp 1636986456
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_333
timestamp 1636986456
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_345
timestamp 1636986456
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_357
timestamp 18001
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 18001
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_365
timestamp 1636986456
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_377
timestamp 18001
transform 1 0 35788 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_394
timestamp 1636986456
transform 1 0 37352 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_406
timestamp 1636986456
transform 1 0 38456 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_418
timestamp 18001
transform 1 0 39560 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_421
timestamp 18001
transform 1 0 39836 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_425
timestamp 18001
transform 1 0 40204 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1636986456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1636986456
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_27
timestamp 18001
transform 1 0 3588 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_31
timestamp 18001
transform 1 0 3956 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_39
timestamp 18001
transform 1 0 4692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_43
timestamp 18001
transform 1 0 5060 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_47
timestamp 18001
transform 1 0 5428 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp 18001
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_83
timestamp 18001
transform 1 0 8740 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_106
timestamp 18001
transform 1 0 10856 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_113
timestamp 18001
transform 1 0 11500 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_121
timestamp 18001
transform 1 0 12236 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_143
timestamp 18001
transform 1 0 14260 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_147
timestamp 18001
transform 1 0 14628 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_166
timestamp 18001
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_183
timestamp 1636986456
transform 1 0 17940 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_195
timestamp 18001
transform 1 0 19044 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_199
timestamp 18001
transform 1 0 19412 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_212
timestamp 1636986456
transform 1 0 20608 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_225
timestamp 18001
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1636986456
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_249
timestamp 18001
transform 1 0 24012 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_262
timestamp 1636986456
transform 1 0 25208 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_274
timestamp 18001
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1636986456
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1636986456
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 1636986456
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 1636986456
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_329
timestamp 18001
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 18001
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 1636986456
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_349
timestamp 18001
transform 1 0 33212 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_355
timestamp 18001
transform 1 0 33764 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_363
timestamp 1636986456
transform 1 0 34500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_375
timestamp 18001
transform 1 0 35604 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_381
timestamp 18001
transform 1 0 36156 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_389
timestamp 18001
transform 1 0 36892 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_393
timestamp 1636986456
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_405
timestamp 18001
transform 1 0 38364 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_413
timestamp 1636986456
transform 1 0 39100 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_425
timestamp 18001
transform 1 0 40204 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1636986456
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1636986456
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 18001
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_29
timestamp 18001
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_37
timestamp 18001
transform 1 0 4508 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_59
timestamp 18001
transform 1 0 6532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_65
timestamp 18001
transform 1 0 7084 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_76
timestamp 18001
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_85
timestamp 18001
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_93
timestamp 18001
transform 1 0 9660 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_105
timestamp 18001
transform 1 0 10764 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_119
timestamp 1636986456
transform 1 0 12052 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_135
timestamp 18001
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 18001
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1636986456
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1636986456
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_165
timestamp 18001
transform 1 0 16284 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_178
timestamp 18001
transform 1 0 17480 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_182
timestamp 18001
transform 1 0 17848 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 18001
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 18001
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_197
timestamp 18001
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_205
timestamp 18001
transform 1 0 19964 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_213
timestamp 1636986456
transform 1 0 20700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_225
timestamp 18001
transform 1 0 21804 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_234
timestamp 1636986456
transform 1 0 22632 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_246
timestamp 18001
transform 1 0 23736 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_270
timestamp 1636986456
transform 1 0 25944 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_282
timestamp 1636986456
transform 1 0 27048 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_294
timestamp 18001
transform 1 0 28152 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 18001
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_309
timestamp 18001
transform 1 0 29532 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_322
timestamp 18001
transform 1 0 30728 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_338
timestamp 18001
transform 1 0 32200 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_348
timestamp 1636986456
transform 1 0 33120 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_360
timestamp 18001
transform 1 0 34224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_365
timestamp 18001
transform 1 0 34684 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_373
timestamp 1636986456
transform 1 0 35420 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_385
timestamp 1636986456
transform 1 0 36524 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_397
timestamp 18001
transform 1 0 37628 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_403
timestamp 18001
transform 1 0 38180 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_416
timestamp 18001
transform 1 0 39376 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_421
timestamp 18001
transform 1 0 39836 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_425
timestamp 18001
transform 1 0 40204 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1636986456
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_15
timestamp 18001
transform 1 0 2484 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_19
timestamp 18001
transform 1 0 2852 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_49
timestamp 18001
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 18001
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1636986456
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_72
timestamp 18001
transform 1 0 7728 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_83
timestamp 18001
transform 1 0 8740 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_89
timestamp 18001
transform 1 0 9292 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_93
timestamp 18001
transform 1 0 9660 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_101
timestamp 18001
transform 1 0 10396 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 18001
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_127
timestamp 18001
transform 1 0 12788 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_143
timestamp 18001
transform 1 0 14260 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_154
timestamp 18001
transform 1 0 15272 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 18001
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1636986456
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1636986456
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1636986456
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1636986456
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 18001
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 18001
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1636986456
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1636986456
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_249
timestamp 18001
transform 1 0 24012 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_256
timestamp 1636986456
transform 1 0 24656 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_268
timestamp 1636986456
transform 1 0 25760 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_287
timestamp 18001
transform 1 0 27508 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_297
timestamp 1636986456
transform 1 0 28428 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_309
timestamp 18001
transform 1 0 29532 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_313
timestamp 18001
transform 1 0 29900 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_321
timestamp 18001
transform 1 0 30636 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_333
timestamp 18001
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 1636986456
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_349
timestamp 18001
transform 1 0 33212 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_357
timestamp 18001
transform 1 0 33948 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_373
timestamp 1636986456
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_393
timestamp 1636986456
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_405
timestamp 1636986456
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_417
timestamp 18001
transform 1 0 39468 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_425
timestamp 18001
transform 1 0 40204 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1636986456
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1636986456
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 18001
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_29
timestamp 18001
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_37
timestamp 18001
transform 1 0 4508 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_60
timestamp 18001
transform 1 0 6624 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_70
timestamp 18001
transform 1 0 7544 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_81
timestamp 18001
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_94
timestamp 18001
transform 1 0 9752 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_152
timestamp 1636986456
transform 1 0 15088 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_164
timestamp 18001
transform 1 0 16192 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_175
timestamp 1636986456
transform 1 0 17204 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_187
timestamp 18001
transform 1 0 18308 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 18001
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1636986456
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_209
timestamp 18001
transform 1 0 20332 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_224
timestamp 18001
transform 1 0 21712 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_241
timestamp 18001
transform 1 0 23276 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_249
timestamp 18001
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_253
timestamp 18001
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_280
timestamp 1636986456
transform 1 0 26864 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_292
timestamp 18001
transform 1 0 27968 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_302
timestamp 18001
transform 1 0 28888 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1636986456
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_321
timestamp 1636986456
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_333
timestamp 1636986456
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_345
timestamp 1636986456
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_357
timestamp 18001
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_363
timestamp 18001
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_365
timestamp 1636986456
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_377
timestamp 18001
transform 1 0 35788 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_383
timestamp 18001
transform 1 0 36340 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_392
timestamp 1636986456
transform 1 0 37168 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_404
timestamp 18001
transform 1 0 38272 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_410
timestamp 18001
transform 1 0 38824 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_418
timestamp 18001
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_421
timestamp 18001
transform 1 0 39836 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_425
timestamp 18001
transform 1 0 40204 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1636986456
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_35
timestamp 1636986456
transform 1 0 4324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_47
timestamp 18001
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 18001
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_57
timestamp 18001
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_73
timestamp 18001
transform 1 0 7820 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_77
timestamp 1636986456
transform 1 0 8188 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_89
timestamp 18001
transform 1 0 9292 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_96
timestamp 18001
transform 1 0 9936 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 18001
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_113
timestamp 18001
transform 1 0 11500 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_119
timestamp 1636986456
transform 1 0 12052 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_131
timestamp 18001
transform 1 0 13156 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_135
timestamp 18001
transform 1 0 13524 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_141
timestamp 1636986456
transform 1 0 14076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_153
timestamp 1636986456
transform 1 0 15180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_165
timestamp 18001
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_169
timestamp 18001
transform 1 0 16652 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_177
timestamp 18001
transform 1 0 17388 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_185
timestamp 18001
transform 1 0 18124 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_198
timestamp 18001
transform 1 0 19320 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_206
timestamp 1636986456
transform 1 0 20056 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_218
timestamp 18001
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1636986456
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_237
timestamp 18001
transform 1 0 22908 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_245
timestamp 18001
transform 1 0 23644 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_260
timestamp 1636986456
transform 1 0 25024 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_272
timestamp 18001
transform 1 0 26128 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_293
timestamp 18001
transform 1 0 28060 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_304
timestamp 18001
transform 1 0 29072 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_312
timestamp 18001
transform 1 0 29808 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_319
timestamp 1636986456
transform 1 0 30452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_331
timestamp 18001
transform 1 0 31556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 18001
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 1636986456
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_349
timestamp 18001
transform 1 0 33212 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_353
timestamp 18001
transform 1 0 33580 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_357
timestamp 1636986456
transform 1 0 33948 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_383
timestamp 18001
transform 1 0 36340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 18001
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_393
timestamp 18001
transform 1 0 37260 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_399
timestamp 18001
transform 1 0 37812 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_406
timestamp 1636986456
transform 1 0 38456 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_418
timestamp 18001
transform 1 0 39560 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1636986456
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1636986456
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 18001
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_46
timestamp 1636986456
transform 1 0 5336 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_58
timestamp 18001
transform 1 0 6440 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_69
timestamp 1636986456
transform 1 0 7452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_85
timestamp 18001
transform 1 0 8924 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_91
timestamp 18001
transform 1 0 9476 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_96
timestamp 18001
transform 1 0 9936 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_104
timestamp 18001
transform 1 0 10672 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_110
timestamp 1636986456
transform 1 0 11224 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_122
timestamp 18001
transform 1 0 12328 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_126
timestamp 18001
transform 1 0 12696 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_136
timestamp 18001
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1636986456
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1636986456
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_165
timestamp 18001
transform 1 0 16284 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_174
timestamp 18001
transform 1 0 17112 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_182
timestamp 18001
transform 1 0 17848 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_190
timestamp 18001
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1636986456
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1636986456
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_221
timestamp 18001
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_244
timestamp 18001
transform 1 0 23552 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_253
timestamp 18001
transform 1 0 24380 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_260
timestamp 1636986456
transform 1 0 25024 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_272
timestamp 18001
transform 1 0 26128 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_279
timestamp 1636986456
transform 1 0 26772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_291
timestamp 18001
transform 1 0 27876 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_295
timestamp 18001
transform 1 0 28244 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_303
timestamp 18001
transform 1 0 28980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 18001
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1636986456
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_321
timestamp 18001
transform 1 0 30636 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_325
timestamp 18001
transform 1 0 31004 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_342
timestamp 18001
transform 1 0 32568 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_349
timestamp 18001
transform 1 0 33212 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 18001
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 1636986456
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_377
timestamp 18001
transform 1 0 35788 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_388
timestamp 1636986456
transform 1 0 36800 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_400
timestamp 18001
transform 1 0 37904 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_409
timestamp 18001
transform 1 0 38732 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_417
timestamp 18001
transform 1 0 39468 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_421
timestamp 18001
transform 1 0 39836 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_425
timestamp 18001
transform 1 0 40204 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1636986456
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_15
timestamp 18001
transform 1 0 2484 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_26
timestamp 18001
transform 1 0 3496 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_49
timestamp 18001
transform 1 0 5612 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 18001
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_74
timestamp 1636986456
transform 1 0 7912 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_86
timestamp 1636986456
transform 1 0 9016 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_98
timestamp 1636986456
transform 1 0 10120 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_110
timestamp 18001
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_113
timestamp 18001
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_144
timestamp 18001
transform 1 0 14352 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_152
timestamp 18001
transform 1 0 15088 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_175
timestamp 1636986456
transform 1 0 17204 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_187
timestamp 1636986456
transform 1 0 18308 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_199
timestamp 1636986456
transform 1 0 19412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_211
timestamp 1636986456
transform 1 0 20516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 18001
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_225
timestamp 18001
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_235
timestamp 1636986456
transform 1 0 22724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_247
timestamp 18001
transform 1 0 23828 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_258
timestamp 1636986456
transform 1 0 24840 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_270
timestamp 18001
transform 1 0 25944 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_286
timestamp 18001
transform 1 0 27416 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_294
timestamp 1636986456
transform 1 0 28152 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_306
timestamp 18001
transform 1 0 29256 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_314
timestamp 18001
transform 1 0 29992 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_323
timestamp 1636986456
transform 1 0 30820 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 18001
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_342
timestamp 1636986456
transform 1 0 32568 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_354
timestamp 1636986456
transform 1 0 33672 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_366
timestamp 1636986456
transform 1 0 34776 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_378
timestamp 1636986456
transform 1 0 35880 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_390
timestamp 18001
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_393
timestamp 18001
transform 1 0 37260 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_401
timestamp 18001
transform 1 0 37996 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_412
timestamp 18001
transform 1 0 39008 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_3
timestamp 18001
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_25
timestamp 18001
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_29
timestamp 18001
transform 1 0 3772 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_64
timestamp 18001
transform 1 0 6992 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_70
timestamp 18001
transform 1 0 7544 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_80
timestamp 18001
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_85
timestamp 18001
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_100
timestamp 18001
transform 1 0 10304 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_134
timestamp 18001
transform 1 0 13432 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1636986456
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_153
timestamp 18001
transform 1 0 15180 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_162
timestamp 1636986456
transform 1 0 16008 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_174
timestamp 1636986456
transform 1 0 17112 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_186
timestamp 18001
transform 1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 18001
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1636986456
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_220
timestamp 18001
transform 1 0 21344 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_231
timestamp 1636986456
transform 1 0 22356 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_243
timestamp 18001
transform 1 0 23460 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 18001
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_264
timestamp 18001
transform 1 0 25392 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_273
timestamp 18001
transform 1 0 26220 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_279
timestamp 18001
transform 1 0 26772 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_285
timestamp 18001
transform 1 0 27324 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_291
timestamp 18001
transform 1 0 27876 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_320
timestamp 18001
transform 1 0 30544 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_324
timestamp 18001
transform 1 0 30912 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_337
timestamp 1636986456
transform 1 0 32108 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_349
timestamp 1636986456
transform 1 0 33212 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_361
timestamp 18001
transform 1 0 34316 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_370
timestamp 18001
transform 1 0 35144 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_374
timestamp 18001
transform 1 0 35512 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_382
timestamp 1636986456
transform 1 0 36248 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_394
timestamp 1636986456
transform 1 0 37352 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_406
timestamp 18001
transform 1 0 38456 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_416
timestamp 18001
transform 1 0 39376 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_421
timestamp 18001
transform 1 0 39836 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_425
timestamp 18001
transform 1 0 40204 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_3
timestamp 18001
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_43
timestamp 18001
transform 1 0 5060 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_52
timestamp 18001
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 18001
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1636986456
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_125
timestamp 18001
transform 1 0 12604 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_133
timestamp 18001
transform 1 0 13340 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_141
timestamp 18001
transform 1 0 14076 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_149
timestamp 18001
transform 1 0 14812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_162
timestamp 18001
transform 1 0 16008 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 18001
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_169
timestamp 18001
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_184
timestamp 18001
transform 1 0 18032 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_190
timestamp 1636986456
transform 1 0 18584 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_202
timestamp 1636986456
transform 1 0 19688 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_214
timestamp 18001
transform 1 0 20792 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_222
timestamp 18001
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_229
timestamp 1636986456
transform 1 0 22172 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_241
timestamp 18001
transform 1 0 23276 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_251
timestamp 1636986456
transform 1 0 24196 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_263
timestamp 1636986456
transform 1 0 25300 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_275
timestamp 18001
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 18001
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_281
timestamp 18001
transform 1 0 26956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_285
timestamp 18001
transform 1 0 27324 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_291
timestamp 18001
transform 1 0 27876 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_299
timestamp 18001
transform 1 0 28612 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_322
timestamp 18001
transform 1 0 30728 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_326
timestamp 18001
transform 1 0 31096 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_332
timestamp 18001
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_337
timestamp 1636986456
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_349
timestamp 18001
transform 1 0 33212 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_372
timestamp 18001
transform 1 0 35328 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_380
timestamp 18001
transform 1 0 36064 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_388
timestamp 18001
transform 1 0 36800 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_393
timestamp 1636986456
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_413
timestamp 1636986456
transform 1 0 39100 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_425
timestamp 18001
transform 1 0 40204 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1636986456
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1636986456
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 18001
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_45
timestamp 18001
transform 1 0 5244 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_68
timestamp 18001
transform 1 0 7360 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_85
timestamp 18001
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_105
timestamp 1636986456
transform 1 0 10764 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_117
timestamp 18001
transform 1 0 11868 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_133
timestamp 18001
transform 1 0 13340 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_160
timestamp 1636986456
transform 1 0 15824 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_172
timestamp 1636986456
transform 1 0 16928 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_184
timestamp 1636986456
transform 1 0 18032 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_197
timestamp 18001
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_205
timestamp 18001
transform 1 0 19964 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_227
timestamp 18001
transform 1 0 21988 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_235
timestamp 18001
transform 1 0 22724 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_242
timestamp 18001
transform 1 0 23368 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_247
timestamp 18001
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 18001
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_266
timestamp 18001
transform 1 0 25576 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_270
timestamp 18001
transform 1 0 25944 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_277
timestamp 18001
transform 1 0 26588 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_296
timestamp 18001
transform 1 0 28336 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_309
timestamp 18001
transform 1 0 29532 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_322
timestamp 18001
transform 1 0 30728 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_333
timestamp 1636986456
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_345
timestamp 1636986456
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_357
timestamp 18001
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_363
timestamp 18001
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_365
timestamp 1636986456
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_377
timestamp 18001
transform 1 0 35788 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_385
timestamp 18001
transform 1 0 36524 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_396
timestamp 18001
transform 1 0 37536 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_404
timestamp 18001
transform 1 0 38272 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_416
timestamp 18001
transform 1 0 39376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_421
timestamp 18001
transform 1 0 39836 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_425
timestamp 18001
transform 1 0 40204 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1636986456
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_15
timestamp 18001
transform 1 0 2484 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 18001
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_63
timestamp 1636986456
transform 1 0 6900 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_75
timestamp 18001
transform 1 0 8004 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 18001
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_113
timestamp 18001
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_125
timestamp 18001
transform 1 0 12604 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1636986456
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_181
timestamp 18001
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_185
timestamp 18001
transform 1 0 18124 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_191
timestamp 1636986456
transform 1 0 18676 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_203
timestamp 18001
transform 1 0 19780 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_216
timestamp 18001
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_225
timestamp 18001
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_233
timestamp 18001
transform 1 0 22540 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_241
timestamp 1636986456
transform 1 0 23276 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_253
timestamp 18001
transform 1 0 24380 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_281
timestamp 18001
transform 1 0 26956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_298
timestamp 18001
transform 1 0 28520 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_306
timestamp 18001
transform 1 0 29256 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_317
timestamp 18001
transform 1 0 30268 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_325
timestamp 18001
transform 1 0 31004 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_335
timestamp 18001
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_337
timestamp 18001
transform 1 0 32108 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_348
timestamp 18001
transform 1 0 33120 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_354
timestamp 18001
transform 1 0 33672 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_360
timestamp 1636986456
transform 1 0 34224 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_372
timestamp 1636986456
transform 1 0 35328 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_384
timestamp 18001
transform 1 0 36432 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_393
timestamp 18001
transform 1 0 37260 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_401
timestamp 18001
transform 1 0 37996 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_410
timestamp 1636986456
transform 1 0 38824 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_422
timestamp 18001
transform 1 0 39928 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_3
timestamp 18001
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_7
timestamp 18001
transform 1 0 1748 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_29
timestamp 18001
transform 1 0 3772 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_35
timestamp 18001
transform 1 0 4324 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_67
timestamp 18001
transform 1 0 7268 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_80
timestamp 18001
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1636986456
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_97
timestamp 18001
transform 1 0 10028 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_141
timestamp 18001
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_151
timestamp 1636986456
transform 1 0 14996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_163
timestamp 18001
transform 1 0 16100 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_171
timestamp 18001
transform 1 0 16836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_177
timestamp 18001
transform 1 0 17388 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_185
timestamp 18001
transform 1 0 18124 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_192
timestamp 18001
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_211
timestamp 18001
transform 1 0 20516 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_234
timestamp 18001
transform 1 0 22632 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_240
timestamp 18001
transform 1 0 23184 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_248
timestamp 18001
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1636986456
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_265
timestamp 18001
transform 1 0 25484 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_278
timestamp 1636986456
transform 1 0 26680 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_290
timestamp 18001
transform 1 0 27784 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_298
timestamp 18001
transform 1 0 28520 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 18001
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_309
timestamp 18001
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_317
timestamp 18001
transform 1 0 30268 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_325
timestamp 18001
transform 1 0 31004 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_342
timestamp 18001
transform 1 0 32568 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_350
timestamp 18001
transform 1 0 33304 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_360
timestamp 18001
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_365
timestamp 18001
transform 1 0 34684 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_373
timestamp 18001
transform 1 0 35420 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_380
timestamp 18001
transform 1 0 36064 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_384
timestamp 18001
transform 1 0 36432 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_391
timestamp 1636986456
transform 1 0 37076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_403
timestamp 18001
transform 1 0 38180 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_411
timestamp 18001
transform 1 0 38916 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_419
timestamp 18001
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_421
timestamp 18001
transform 1 0 39836 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_425
timestamp 18001
transform 1 0 40204 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_3
timestamp 18001
transform 1 0 1380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_24
timestamp 18001
transform 1 0 3312 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_57
timestamp 18001
transform 1 0 6348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_61
timestamp 18001
transform 1 0 6716 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_99
timestamp 1636986456
transform 1 0 10212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 18001
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1636986456
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_125
timestamp 18001
transform 1 0 12604 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_132
timestamp 18001
transform 1 0 13248 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_140
timestamp 18001
transform 1 0 13984 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_147
timestamp 1636986456
transform 1 0 14628 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_159
timestamp 18001
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 18001
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_175
timestamp 1636986456
transform 1 0 17204 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_187
timestamp 1636986456
transform 1 0 18308 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_199
timestamp 1636986456
transform 1 0 19412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_211
timestamp 18001
transform 1 0 20516 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_222
timestamp 18001
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1636986456
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_237
timestamp 18001
transform 1 0 22908 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_245
timestamp 18001
transform 1 0 23644 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_250
timestamp 1636986456
transform 1 0 24104 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_262
timestamp 1636986456
transform 1 0 25208 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_274
timestamp 18001
transform 1 0 26312 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_281
timestamp 18001
transform 1 0 26956 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_298
timestamp 1636986456
transform 1 0 28520 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_310
timestamp 1636986456
transform 1 0 29624 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_322
timestamp 18001
transform 1 0 30728 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_330
timestamp 18001
transform 1 0 31464 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_335
timestamp 18001
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 1636986456
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_349
timestamp 18001
transform 1 0 33212 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_360
timestamp 18001
transform 1 0 34224 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_370
timestamp 18001
transform 1 0 35144 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_388
timestamp 18001
transform 1 0 36800 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_393
timestamp 1636986456
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_405
timestamp 1636986456
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_417
timestamp 18001
transform 1 0 39468 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_425
timestamp 18001
transform 1 0 40204 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_3
timestamp 18001
transform 1 0 1380 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_24
timestamp 18001
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_29
timestamp 18001
transform 1 0 3772 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_69
timestamp 18001
transform 1 0 7452 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_75
timestamp 18001
transform 1 0 8004 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 18001
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_115
timestamp 18001
transform 1 0 11684 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_121
timestamp 18001
transform 1 0 12236 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_141
timestamp 18001
transform 1 0 14076 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_155
timestamp 1636986456
transform 1 0 15364 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_167
timestamp 18001
transform 1 0 16468 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_187
timestamp 18001
transform 1 0 18308 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 18001
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_197
timestamp 18001
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_201
timestamp 18001
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_215
timestamp 18001
transform 1 0 20884 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_223
timestamp 18001
transform 1 0 21620 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_227
timestamp 18001
transform 1 0 21988 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_250
timestamp 18001
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_274
timestamp 18001
transform 1 0 26312 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_288
timestamp 1636986456
transform 1 0 27600 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_300
timestamp 18001
transform 1 0 28704 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_309
timestamp 18001
transform 1 0 29532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_323
timestamp 18001
transform 1 0 30820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_331
timestamp 18001
transform 1 0 31556 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_339
timestamp 1636986456
transform 1 0 32292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_351
timestamp 1636986456
transform 1 0 33396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 18001
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_365
timestamp 1636986456
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_377
timestamp 1636986456
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_389
timestamp 18001
transform 1 0 36892 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_397
timestamp 18001
transform 1 0 37628 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_417
timestamp 18001
transform 1 0 39468 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_421
timestamp 18001
transform 1 0 39836 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_425
timestamp 18001
transform 1 0 40204 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_3
timestamp 18001
transform 1 0 1380 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_11
timestamp 18001
transform 1 0 2116 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1636986456
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_69
timestamp 18001
transform 1 0 7452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_77
timestamp 18001
transform 1 0 8188 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_86
timestamp 18001
transform 1 0 9016 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_98
timestamp 18001
transform 1 0 10120 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_110
timestamp 18001
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_113
timestamp 18001
transform 1 0 11500 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_126
timestamp 1636986456
transform 1 0 12696 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_143
timestamp 1636986456
transform 1 0 14260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_155
timestamp 1636986456
transform 1 0 15364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 18001
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 1636986456
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 1636986456
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 1636986456
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_205
timestamp 18001
transform 1 0 19964 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_222
timestamp 18001
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 1636986456
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 1636986456
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_255
timestamp 18001
transform 1 0 24564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_263
timestamp 18001
transform 1 0 25300 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_281
timestamp 18001
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_307
timestamp 18001
transform 1 0 29348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_324
timestamp 18001
transform 1 0 30912 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_328
timestamp 18001
transform 1 0 31280 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_351
timestamp 1636986456
transform 1 0 33396 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_363
timestamp 1636986456
transform 1 0 34500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_375
timestamp 18001
transform 1 0 35604 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_385
timestamp 18001
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_391
timestamp 18001
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_393
timestamp 18001
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_406
timestamp 1636986456
transform 1 0 38456 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_418
timestamp 18001
transform 1 0 39560 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_3
timestamp 18001
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_11
timestamp 18001
transform 1 0 2116 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_29
timestamp 18001
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_70
timestamp 1636986456
transform 1 0 7544 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_82
timestamp 18001
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_88
timestamp 18001
transform 1 0 9200 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_92
timestamp 18001
transform 1 0 9568 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_122
timestamp 18001
transform 1 0 12328 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_134
timestamp 18001
transform 1 0 13432 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_150
timestamp 1636986456
transform 1 0 14904 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_162
timestamp 18001
transform 1 0 16008 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_175
timestamp 18001
transform 1 0 17204 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_193
timestamp 18001
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1636986456
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 1636986456
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_221
timestamp 18001
transform 1 0 21436 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_229
timestamp 18001
transform 1 0 22172 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_233
timestamp 1636986456
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_245
timestamp 18001
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 18001
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1636986456
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_265
timestamp 1636986456
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_277
timestamp 1636986456
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_289
timestamp 1636986456
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_301
timestamp 18001
transform 1 0 28796 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 18001
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_309
timestamp 18001
transform 1 0 29532 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_320
timestamp 18001
transform 1 0 30544 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_326
timestamp 18001
transform 1 0 31096 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_334
timestamp 18001
transform 1 0 31832 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_342
timestamp 18001
transform 1 0 32568 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_353
timestamp 18001
transform 1 0 33580 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_361
timestamp 18001
transform 1 0 34316 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_365
timestamp 1636986456
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_377
timestamp 18001
transform 1 0 35788 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_388
timestamp 1636986456
transform 1 0 36800 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_400
timestamp 18001
transform 1 0 37904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_410
timestamp 18001
transform 1 0 38824 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_421
timestamp 18001
transform 1 0 39836 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_425
timestamp 18001
transform 1 0 40204 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1636986456
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_24
timestamp 18001
transform 1 0 3312 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_47
timestamp 18001
transform 1 0 5428 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_64
timestamp 18001
transform 1 0 6992 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_72
timestamp 18001
transform 1 0 7728 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_88
timestamp 1636986456
transform 1 0 9200 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_100
timestamp 18001
transform 1 0 10304 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_113
timestamp 18001
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_119
timestamp 18001
transform 1 0 12052 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_148
timestamp 18001
transform 1 0 14720 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_162
timestamp 18001
transform 1 0 16008 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_169
timestamp 18001
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_201
timestamp 18001
transform 1 0 19596 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_208
timestamp 18001
transform 1 0 20240 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_215
timestamp 18001
transform 1 0 20884 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 18001
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_225
timestamp 18001
transform 1 0 21804 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_245
timestamp 18001
transform 1 0 23644 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_252
timestamp 1636986456
transform 1 0 24288 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_264
timestamp 1636986456
transform 1 0 25392 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_276
timestamp 18001
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_286
timestamp 18001
transform 1 0 27416 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_290
timestamp 18001
transform 1 0 27784 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_311
timestamp 1636986456
transform 1 0 29716 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_323
timestamp 18001
transform 1 0 30820 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_328
timestamp 18001
transform 1 0 31280 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_337
timestamp 18001
transform 1 0 32108 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_345
timestamp 18001
transform 1 0 32844 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_353
timestamp 18001
transform 1 0 33580 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_370
timestamp 1636986456
transform 1 0 35144 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_382
timestamp 18001
transform 1 0 36248 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_388
timestamp 18001
transform 1 0 36800 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_393
timestamp 18001
transform 1 0 37260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_401
timestamp 18001
transform 1 0 37996 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_23
timestamp 18001
transform 1 0 3220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 18001
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_64
timestamp 18001
transform 1 0 6992 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_72
timestamp 18001
transform 1 0 7728 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_94
timestamp 1636986456
transform 1 0 9752 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_106
timestamp 18001
transform 1 0 10856 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_112
timestamp 1636986456
transform 1 0 11408 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_124
timestamp 1636986456
transform 1 0 12512 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_136
timestamp 18001
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_149
timestamp 18001
transform 1 0 14812 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_163
timestamp 18001
transform 1 0 16100 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_169
timestamp 1636986456
transform 1 0 16652 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_187
timestamp 18001
transform 1 0 18308 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_194
timestamp 18001
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_197
timestamp 18001
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_212
timestamp 1636986456
transform 1 0 20608 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_224
timestamp 1636986456
transform 1 0 21712 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_236
timestamp 18001
transform 1 0 22816 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 18001
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_253
timestamp 18001
transform 1 0 24380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_278
timestamp 18001
transform 1 0 26680 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_291
timestamp 18001
transform 1 0 27876 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 18001
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 1636986456
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_321
timestamp 1636986456
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_333
timestamp 1636986456
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_345
timestamp 1636986456
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_357
timestamp 18001
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_363
timestamp 18001
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_365
timestamp 1636986456
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_377
timestamp 1636986456
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_389
timestamp 18001
transform 1 0 36892 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_397
timestamp 18001
transform 1 0 37628 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_408
timestamp 18001
transform 1 0 38640 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_421
timestamp 18001
transform 1 0 39836 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1636986456
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_15
timestamp 18001
transform 1 0 2484 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_33
timestamp 1636986456
transform 1 0 4140 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_45
timestamp 18001
transform 1 0 5244 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_54
timestamp 18001
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_57
timestamp 18001
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_65
timestamp 18001
transform 1 0 7084 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_95
timestamp 18001
transform 1 0 9844 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_101
timestamp 18001
transform 1 0 10396 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_109
timestamp 18001
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_128
timestamp 1636986456
transform 1 0 12880 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_140
timestamp 18001
transform 1 0 13984 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_144
timestamp 18001
transform 1 0 14352 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_152
timestamp 18001
transform 1 0 15088 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_159
timestamp 18001
transform 1 0 15732 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_181
timestamp 1636986456
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_193
timestamp 18001
transform 1 0 18860 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_199
timestamp 18001
transform 1 0 19412 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_210
timestamp 18001
transform 1 0 20424 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 18001
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_233
timestamp 1636986456
transform 1 0 22540 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_245
timestamp 18001
transform 1 0 23644 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_251
timestamp 18001
transform 1 0 24196 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_297
timestamp 18001
transform 1 0 28428 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_302
timestamp 1636986456
transform 1 0 28888 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_314
timestamp 18001
transform 1 0 29992 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_322
timestamp 18001
transform 1 0 30728 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 18001
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1636986456
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 1636986456
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_361
timestamp 18001
transform 1 0 34316 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_369
timestamp 18001
transform 1 0 35052 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_376
timestamp 1636986456
transform 1 0 35696 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_388
timestamp 18001
transform 1 0 36800 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_399
timestamp 18001
transform 1 0 37812 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_415
timestamp 18001
transform 1 0 39284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_421
timestamp 18001
transform 1 0 39836 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_3
timestamp 18001
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_25
timestamp 18001
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_46
timestamp 18001
transform 1 0 5336 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_69
timestamp 18001
transform 1 0 7452 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_73
timestamp 18001
transform 1 0 7820 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 18001
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_93
timestamp 1636986456
transform 1 0 9660 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_105
timestamp 18001
transform 1 0 10764 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_113
timestamp 1636986456
transform 1 0 11500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_125
timestamp 1636986456
transform 1 0 12604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_137
timestamp 18001
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1636986456
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_153
timestamp 18001
transform 1 0 15180 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_159
timestamp 18001
transform 1 0 15732 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_163
timestamp 18001
transform 1 0 16100 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_168
timestamp 1636986456
transform 1 0 16560 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_180
timestamp 18001
transform 1 0 17664 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_186
timestamp 18001
transform 1 0 18216 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_192
timestamp 18001
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_197
timestamp 18001
transform 1 0 19228 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_205
timestamp 18001
transform 1 0 19964 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_211
timestamp 1636986456
transform 1 0 20516 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_223
timestamp 1636986456
transform 1 0 21620 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_235
timestamp 18001
transform 1 0 22724 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_239
timestamp 18001
transform 1 0 23092 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_247
timestamp 18001
transform 1 0 23828 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 18001
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_253
timestamp 18001
transform 1 0 24380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_257
timestamp 18001
transform 1 0 24748 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_280
timestamp 1636986456
transform 1 0 26864 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_292
timestamp 1636986456
transform 1 0 27968 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_304
timestamp 18001
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_309
timestamp 18001
transform 1 0 29532 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_315
timestamp 18001
transform 1 0 30084 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_331
timestamp 18001
transform 1 0 31556 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_338
timestamp 18001
transform 1 0 32200 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_358
timestamp 18001
transform 1 0 34040 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_365
timestamp 18001
transform 1 0 34684 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_371
timestamp 18001
transform 1 0 35236 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_388
timestamp 1636986456
transform 1 0 36800 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_400
timestamp 18001
transform 1 0 37904 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_406
timestamp 1636986456
transform 1 0 38456 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_418
timestamp 18001
transform 1 0 39560 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_421
timestamp 18001
transform 1 0 39836 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_425
timestamp 18001
transform 1 0 40204 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_3
timestamp 18001
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_25
timestamp 18001
transform 1 0 3404 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_73
timestamp 1636986456
transform 1 0 7820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_85
timestamp 1636986456
transform 1 0 8924 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_101
timestamp 18001
transform 1 0 10396 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_109
timestamp 18001
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_118
timestamp 18001
transform 1 0 11960 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_126
timestamp 18001
transform 1 0 12696 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_132
timestamp 18001
transform 1 0 13248 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_149
timestamp 18001
transform 1 0 14812 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_155
timestamp 18001
transform 1 0 15364 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_162
timestamp 18001
transform 1 0 16008 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1636986456
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_181
timestamp 18001
transform 1 0 17756 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_189
timestamp 18001
transform 1 0 18492 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_198
timestamp 1636986456
transform 1 0 19320 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_210
timestamp 1636986456
transform 1 0 20424 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_222
timestamp 18001
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1636986456
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1636986456
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 1636986456
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_261
timestamp 18001
transform 1 0 25116 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_269
timestamp 18001
transform 1 0 25852 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 18001
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 18001
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1636986456
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_293
timestamp 18001
transform 1 0 28060 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_298
timestamp 18001
transform 1 0 28520 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_302
timestamp 18001
transform 1 0 28888 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_325
timestamp 18001
transform 1 0 31004 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_334
timestamp 18001
transform 1 0 31832 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_337
timestamp 18001
transform 1 0 32108 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_342
timestamp 1636986456
transform 1 0 32568 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_354
timestamp 18001
transform 1 0 33672 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_372
timestamp 18001
transform 1 0 35328 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_379
timestamp 1636986456
transform 1 0 35972 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_391
timestamp 18001
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_393
timestamp 18001
transform 1 0 37260 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_407
timestamp 1636986456
transform 1 0 38548 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_419
timestamp 18001
transform 1 0 39652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_425
timestamp 18001
transform 1 0 40204 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1636986456
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_15
timestamp 18001
transform 1 0 2484 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_26
timestamp 18001
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_37
timestamp 18001
transform 1 0 4508 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_45
timestamp 18001
transform 1 0 5244 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_66
timestamp 18001
transform 1 0 7176 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_74
timestamp 18001
transform 1 0 7912 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 18001
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_90
timestamp 18001
transform 1 0 9384 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_94
timestamp 18001
transform 1 0 9752 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_99
timestamp 18001
transform 1 0 10212 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_108
timestamp 18001
transform 1 0 11040 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_113
timestamp 18001
transform 1 0 11500 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_126
timestamp 1636986456
transform 1 0 12696 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_138
timestamp 18001
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_149
timestamp 18001
transform 1 0 14812 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_177
timestamp 18001
transform 1 0 17388 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_186
timestamp 18001
transform 1 0 18216 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_197
timestamp 18001
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_205
timestamp 18001
transform 1 0 19964 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_220
timestamp 18001
transform 1 0 21344 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_228
timestamp 18001
transform 1 0 22080 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_246
timestamp 18001
transform 1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_270
timestamp 18001
transform 1 0 25944 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_282
timestamp 18001
transform 1 0 27048 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_305
timestamp 18001
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_309
timestamp 18001
transform 1 0 29532 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_314
timestamp 1636986456
transform 1 0 29992 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_335
timestamp 18001
transform 1 0 31924 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_345
timestamp 1636986456
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_357
timestamp 18001
transform 1 0 33948 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_378
timestamp 1636986456
transform 1 0 35880 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_390
timestamp 18001
transform 1 0 36984 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_396
timestamp 18001
transform 1 0 37536 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_406
timestamp 1636986456
transform 1 0 38456 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_418
timestamp 18001
transform 1 0 39560 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_421
timestamp 18001
transform 1 0 39836 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1636986456
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1636986456
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_27
timestamp 18001
transform 1 0 3588 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_40
timestamp 18001
transform 1 0 4784 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_48
timestamp 18001
transform 1 0 5520 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_57
timestamp 18001
transform 1 0 6348 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_63
timestamp 1636986456
transform 1 0 6900 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_75
timestamp 18001
transform 1 0 8004 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_88
timestamp 18001
transform 1 0 9200 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_92
timestamp 18001
transform 1 0 9568 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_96
timestamp 18001
transform 1 0 9936 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 18001
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_120
timestamp 1636986456
transform 1 0 12144 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_132
timestamp 18001
transform 1 0 13248 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_137
timestamp 18001
transform 1 0 13708 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_145
timestamp 18001
transform 1 0 14444 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_157
timestamp 18001
transform 1 0 15548 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_165
timestamp 18001
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_177
timestamp 18001
transform 1 0 17388 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_183
timestamp 18001
transform 1 0 17940 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_193
timestamp 18001
transform 1 0 18860 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_202
timestamp 18001
transform 1 0 19688 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_221
timestamp 18001
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_230
timestamp 18001
transform 1 0 22264 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_247
timestamp 18001
transform 1 0 23828 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_259
timestamp 18001
transform 1 0 24932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_263
timestamp 18001
transform 1 0 25300 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_270
timestamp 18001
transform 1 0 25944 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_278
timestamp 18001
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1636986456
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 1636986456
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_305
timestamp 18001
transform 1 0 29164 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_311
timestamp 18001
transform 1 0 29716 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_321
timestamp 18001
transform 1 0 30636 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_330
timestamp 18001
transform 1 0 31464 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_343
timestamp 1636986456
transform 1 0 32660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_355
timestamp 18001
transform 1 0 33764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_361
timestamp 18001
transform 1 0 34316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_365
timestamp 1636986456
transform 1 0 34684 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_377
timestamp 18001
transform 1 0 35788 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_420
timestamp 18001
transform 1 0 39744 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1636986456
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1636986456
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 18001
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_49
timestamp 1636986456
transform 1 0 5612 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_61
timestamp 18001
transform 1 0 6716 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_85
timestamp 18001
transform 1 0 8924 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_95
timestamp 1636986456
transform 1 0 9844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_113
timestamp 18001
transform 1 0 11500 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_121
timestamp 18001
transform 1 0 12236 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_125
timestamp 18001
transform 1 0 12604 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_136
timestamp 18001
transform 1 0 13616 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_141
timestamp 18001
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_150
timestamp 18001
transform 1 0 14904 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_161
timestamp 1636986456
transform 1 0 15916 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_173
timestamp 18001
transform 1 0 17020 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 18001
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_205
timestamp 18001
transform 1 0 19964 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_213
timestamp 1636986456
transform 1 0 20700 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_225
timestamp 1636986456
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_237
timestamp 1636986456
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_249
timestamp 18001
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_253
timestamp 18001
transform 1 0 24380 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_261
timestamp 18001
transform 1 0 25116 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_268
timestamp 1636986456
transform 1 0 25760 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_280
timestamp 1636986456
transform 1 0 26864 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_292
timestamp 1636986456
transform 1 0 27968 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_304
timestamp 18001
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_329
timestamp 18001
transform 1 0 31372 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_345
timestamp 18001
transform 1 0 32844 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_353
timestamp 18001
transform 1 0 33580 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_361
timestamp 18001
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 1636986456
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_377
timestamp 18001
transform 1 0 35788 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_385
timestamp 18001
transform 1 0 36524 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_395
timestamp 1636986456
transform 1 0 37444 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_407
timestamp 18001
transform 1 0 38548 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_413
timestamp 18001
transform 1 0 39100 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_421
timestamp 18001
transform 1 0 39836 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_425
timestamp 18001
transform 1 0 40204 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1636986456
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_44
timestamp 1636986456
transform 1 0 5152 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_66
timestamp 1636986456
transform 1 0 7176 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_78
timestamp 1636986456
transform 1 0 8280 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_90
timestamp 1636986456
transform 1 0 9384 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_102
timestamp 18001
transform 1 0 10488 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_110
timestamp 18001
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_120
timestamp 18001
transform 1 0 12144 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_126
timestamp 18001
transform 1 0 12696 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_151
timestamp 18001
transform 1 0 14996 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_163
timestamp 18001
transform 1 0 16100 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 18001
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_177
timestamp 18001
transform 1 0 17388 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_185
timestamp 18001
transform 1 0 18124 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_196
timestamp 18001
transform 1 0 19136 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_208
timestamp 18001
transform 1 0 20240 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_235
timestamp 18001
transform 1 0 22724 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_239
timestamp 1636986456
transform 1 0 23092 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_251
timestamp 18001
transform 1 0 24196 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_259
timestamp 18001
transform 1 0 24932 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_269
timestamp 18001
transform 1 0 25852 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_277
timestamp 18001
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1636986456
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_293
timestamp 18001
transform 1 0 28060 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_331
timestamp 18001
transform 1 0 31556 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 18001
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_337
timestamp 18001
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_346
timestamp 1636986456
transform 1 0 32936 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_358
timestamp 1636986456
transform 1 0 34040 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_370
timestamp 1636986456
transform 1 0 35144 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_382
timestamp 18001
transform 1 0 36248 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_390
timestamp 18001
transform 1 0 36984 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_393
timestamp 1636986456
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_405
timestamp 1636986456
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_417
timestamp 18001
transform 1 0 39468 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_425
timestamp 18001
transform 1 0 40204 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1636986456
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1636986456
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 18001
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1636986456
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_41
timestamp 18001
transform 1 0 4876 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_47
timestamp 18001
transform 1 0 5428 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_68
timestamp 18001
transform 1 0 7360 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_79
timestamp 18001
transform 1 0 8372 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 18001
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_85
timestamp 18001
transform 1 0 8924 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_89
timestamp 18001
transform 1 0 9292 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_110
timestamp 18001
transform 1 0 11224 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 1636986456
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 18001
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 18001
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_148
timestamp 1636986456
transform 1 0 14720 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_160
timestamp 1636986456
transform 1 0 15824 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_172
timestamp 18001
transform 1 0 16928 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_183
timestamp 1636986456
transform 1 0 17940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 18001
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 1636986456
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_209
timestamp 18001
transform 1 0 20332 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_219
timestamp 18001
transform 1 0 21252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_225
timestamp 18001
transform 1 0 21804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_233
timestamp 18001
transform 1 0 22540 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_246
timestamp 18001
transform 1 0 23736 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_253
timestamp 18001
transform 1 0 24380 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_275
timestamp 18001
transform 1 0 26404 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_282
timestamp 18001
transform 1 0 27048 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_300
timestamp 18001
transform 1 0 28704 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_317
timestamp 18001
transform 1 0 30268 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_322
timestamp 1636986456
transform 1 0 30728 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_334
timestamp 18001
transform 1 0 31832 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_346
timestamp 18001
transform 1 0 32936 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_357
timestamp 18001
transform 1 0 33948 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_362
timestamp 18001
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_365
timestamp 18001
transform 1 0 34684 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_373
timestamp 18001
transform 1 0 35420 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_380
timestamp 1636986456
transform 1 0 36064 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_392
timestamp 18001
transform 1 0 37168 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_400
timestamp 18001
transform 1 0 37904 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_411
timestamp 18001
transform 1 0 38916 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_419
timestamp 18001
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_421
timestamp 18001
transform 1 0 39836 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_425
timestamp 18001
transform 1 0 40204 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1636986456
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1636986456
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_27
timestamp 18001
transform 1 0 3588 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_35
timestamp 18001
transform 1 0 4324 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_57
timestamp 18001
transform 1 0 6348 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_61
timestamp 18001
transform 1 0 6716 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_102
timestamp 18001
transform 1 0 10488 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_118
timestamp 18001
transform 1 0 11960 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_128
timestamp 1636986456
transform 1 0 12880 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_140
timestamp 18001
transform 1 0 13984 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_148
timestamp 18001
transform 1 0 14720 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_163
timestamp 18001
transform 1 0 16100 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 18001
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_185
timestamp 18001
transform 1 0 18124 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_189
timestamp 18001
transform 1 0 18492 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_199
timestamp 18001
transform 1 0 19412 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_203
timestamp 18001
transform 1 0 19780 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_211
timestamp 18001
transform 1 0 20516 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_233
timestamp 18001
transform 1 0 22540 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_270
timestamp 18001
transform 1 0 25944 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_274
timestamp 18001
transform 1 0 26312 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_281
timestamp 18001
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 1636986456
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 1636986456
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_329
timestamp 18001
transform 1 0 31372 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_337
timestamp 18001
transform 1 0 32108 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_346
timestamp 18001
transform 1 0 32936 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_361
timestamp 18001
transform 1 0 34316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_369
timestamp 18001
transform 1 0 35052 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_390
timestamp 18001
transform 1 0 36984 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_399
timestamp 18001
transform 1 0 37812 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1636986456
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1636986456
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 18001
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_58
timestamp 1636986456
transform 1 0 6440 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_70
timestamp 1636986456
transform 1 0 7544 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_82
timestamp 18001
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_85
timestamp 18001
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_93
timestamp 18001
transform 1 0 9660 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_125
timestamp 18001
transform 1 0 12604 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_129
timestamp 18001
transform 1 0 12972 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_138
timestamp 18001
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_147
timestamp 18001
transform 1 0 14628 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_151
timestamp 18001
transform 1 0 14996 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_183
timestamp 18001
transform 1 0 17940 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_202
timestamp 1636986456
transform 1 0 19688 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_214
timestamp 1636986456
transform 1 0 20792 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_226
timestamp 18001
transform 1 0 21896 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_249
timestamp 18001
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_264
timestamp 18001
transform 1 0 25392 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_305
timestamp 18001
transform 1 0 29164 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_309
timestamp 18001
transform 1 0 29532 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_317
timestamp 18001
transform 1 0 30268 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_350
timestamp 18001
transform 1 0 33304 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_363
timestamp 18001
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_371
timestamp 18001
transform 1 0 35236 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_387
timestamp 18001
transform 1 0 36708 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_395
timestamp 18001
transform 1 0 37444 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_421
timestamp 18001
transform 1 0 39836 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_425
timestamp 18001
transform 1 0 40204 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_9
timestamp 18001
transform 1 0 1932 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_23
timestamp 18001
transform 1 0 3220 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_31
timestamp 18001
transform 1 0 3956 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_42
timestamp 1636986456
transform 1 0 4968 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_54
timestamp 18001
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_57
timestamp 18001
transform 1 0 6348 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_65
timestamp 18001
transform 1 0 7084 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_71
timestamp 1636986456
transform 1 0 7636 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_83
timestamp 1636986456
transform 1 0 8740 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_95
timestamp 18001
transform 1 0 9844 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_101
timestamp 18001
transform 1 0 10396 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_108
timestamp 18001
transform 1 0 11040 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_113
timestamp 18001
transform 1 0 11500 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_148
timestamp 18001
transform 1 0 14720 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_175
timestamp 18001
transform 1 0 17204 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_183
timestamp 18001
transform 1 0 17940 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_192
timestamp 1636986456
transform 1 0 18768 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_204
timestamp 1636986456
transform 1 0 19872 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_216
timestamp 18001
transform 1 0 20976 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1636986456
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_245
timestamp 1636986456
transform 1 0 23644 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_257
timestamp 18001
transform 1 0 24748 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_272
timestamp 18001
transform 1 0 26128 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_277
timestamp 18001
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1636986456
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_293
timestamp 18001
transform 1 0 28060 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 18001
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_344
timestamp 18001
transform 1 0 32752 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_350
timestamp 18001
transform 1 0 33304 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_358
timestamp 18001
transform 1 0 34040 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_365
timestamp 1636986456
transform 1 0 34684 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_377
timestamp 18001
transform 1 0 35788 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_381
timestamp 18001
transform 1 0 36156 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_387
timestamp 18001
transform 1 0 36708 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_391
timestamp 18001
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_3
timestamp 18001
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_29
timestamp 18001
transform 1 0 3772 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_42
timestamp 1636986456
transform 1 0 4968 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_57
timestamp 18001
transform 1 0 6348 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_65
timestamp 18001
transform 1 0 7084 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_78
timestamp 18001
transform 1 0 8280 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_82
timestamp 18001
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_85
timestamp 18001
transform 1 0 8924 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_91
timestamp 18001
transform 1 0 9476 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_113
timestamp 1636986456
transform 1 0 11500 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_125
timestamp 18001
transform 1 0 12604 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_129
timestamp 18001
transform 1 0 12972 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 18001
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 18001
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1636986456
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_160
timestamp 1636986456
transform 1 0 15824 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_172
timestamp 18001
transform 1 0 16928 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_180
timestamp 18001
transform 1 0 17664 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_194
timestamp 18001
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_218
timestamp 18001
transform 1 0 21160 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_227
timestamp 18001
transform 1 0 21988 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_235
timestamp 18001
transform 1 0 22724 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_250
timestamp 18001
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_259
timestamp 1636986456
transform 1 0 24932 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_271
timestamp 18001
transform 1 0 26036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_281
timestamp 18001
transform 1 0 26956 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_292
timestamp 18001
transform 1 0 27968 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_304
timestamp 18001
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_334
timestamp 1636986456
transform 1 0 31832 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_346
timestamp 18001
transform 1 0 32936 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_352
timestamp 18001
transform 1 0 33488 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_361
timestamp 18001
transform 1 0 34316 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_365
timestamp 18001
transform 1 0 34684 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_379
timestamp 18001
transform 1 0 35972 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_392
timestamp 18001
transform 1 0 37168 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_402
timestamp 18001
transform 1 0 38088 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_412
timestamp 18001
transform 1 0 39008 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_421
timestamp 18001
transform 1 0 39836 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_425
timestamp 18001
transform 1 0 40204 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1636986456
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_15
timestamp 18001
transform 1 0 2484 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 18001
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 18001
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_83
timestamp 18001
transform 1 0 8740 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_121
timestamp 18001
transform 1 0 12236 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_125
timestamp 18001
transform 1 0 12604 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_136
timestamp 18001
transform 1 0 13616 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_145
timestamp 18001
transform 1 0 14444 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_151
timestamp 18001
transform 1 0 14996 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_164
timestamp 18001
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_181
timestamp 18001
transform 1 0 17756 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_191
timestamp 18001
transform 1 0 18676 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_200
timestamp 18001
transform 1 0 19504 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_234
timestamp 18001
transform 1 0 22632 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_238
timestamp 18001
transform 1 0 23000 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_265
timestamp 18001
transform 1 0 25484 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_271
timestamp 18001
transform 1 0 26036 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_302
timestamp 18001
transform 1 0 28888 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_308
timestamp 18001
transform 1 0 29440 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_312
timestamp 1636986456
transform 1 0 29808 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_324
timestamp 1636986456
transform 1 0 30912 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 1636986456
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_355
timestamp 18001
transform 1 0 33764 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_359
timestamp 18001
transform 1 0 34132 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_370
timestamp 18001
transform 1 0 35144 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_378
timestamp 18001
transform 1 0 35880 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_400
timestamp 18001
transform 1 0 37904 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1636986456
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1636986456
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 18001
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_29
timestamp 18001
transform 1 0 3772 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_35
timestamp 18001
transform 1 0 4324 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_42
timestamp 18001
transform 1 0 4968 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_88
timestamp 18001
transform 1 0 9200 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_96
timestamp 18001
transform 1 0 9936 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_117
timestamp 18001
transform 1 0 11868 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_149
timestamp 18001
transform 1 0 14812 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_173
timestamp 18001
transform 1 0 17020 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 18001
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_197
timestamp 18001
transform 1 0 19228 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_226
timestamp 18001
transform 1 0 21896 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_245
timestamp 18001
transform 1 0 23644 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 18001
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_253
timestamp 18001
transform 1 0 24380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_278
timestamp 18001
transform 1 0 26680 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_304
timestamp 18001
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_314
timestamp 18001
transform 1 0 29992 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_318
timestamp 18001
transform 1 0 30360 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_323
timestamp 18001
transform 1 0 30820 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_351
timestamp 1636986456
transform 1 0 33396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 18001
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_365
timestamp 18001
transform 1 0 34684 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_381
timestamp 18001
transform 1 0 36156 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_403
timestamp 18001
transform 1 0 38180 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_411
timestamp 18001
transform 1 0 38916 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_419
timestamp 18001
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_421
timestamp 18001
transform 1 0 39836 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_425
timestamp 18001
transform 1 0 40204 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_3
timestamp 18001
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_7
timestamp 18001
transform 1 0 1748 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_31
timestamp 1636986456
transform 1 0 3956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_43
timestamp 18001
transform 1 0 5060 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 18001
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_62
timestamp 18001
transform 1 0 6808 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_88
timestamp 1636986456
transform 1 0 9200 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_100
timestamp 1636986456
transform 1 0 10304 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_133
timestamp 18001
transform 1 0 13340 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_156
timestamp 1636986456
transform 1 0 15456 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1636986456
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 1636986456
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_193
timestamp 1636986456
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_205
timestamp 18001
transform 1 0 19964 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_213
timestamp 18001
transform 1 0 20700 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_221
timestamp 18001
transform 1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_246
timestamp 18001
transform 1 0 23736 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_262
timestamp 18001
transform 1 0 25208 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_281
timestamp 18001
transform 1 0 26956 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_289
timestamp 18001
transform 1 0 27692 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_304
timestamp 18001
transform 1 0 29072 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 18001
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_356
timestamp 18001
transform 1 0 33856 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_384
timestamp 18001
transform 1 0 36432 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_400
timestamp 1636986456
transform 1 0 37904 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_412
timestamp 1636986456
transform 1 0 39008 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_424
timestamp 18001
transform 1 0 40112 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_3
timestamp 18001
transform 1 0 1380 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 18001
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_29
timestamp 18001
transform 1 0 3772 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_51
timestamp 18001
transform 1 0 5796 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1636986456
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1636986456
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_109
timestamp 18001
transform 1 0 11132 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_118
timestamp 1636986456
transform 1 0 11960 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_130
timestamp 18001
transform 1 0 13064 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_138
timestamp 18001
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1636986456
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_153
timestamp 18001
transform 1 0 15180 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_160
timestamp 18001
transform 1 0 15824 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_168
timestamp 18001
transform 1 0 16560 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_176
timestamp 18001
transform 1 0 17296 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_188
timestamp 18001
transform 1 0 18400 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1636986456
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 1636986456
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 1636986456
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 1636986456
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_249
timestamp 18001
transform 1 0 24012 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_253
timestamp 18001
transform 1 0 24380 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_261
timestamp 18001
transform 1 0 25116 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_268
timestamp 18001
transform 1 0 25760 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_275
timestamp 1636986456
transform 1 0 26404 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_287
timestamp 18001
transform 1 0 27508 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_295
timestamp 18001
transform 1 0 28244 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_306
timestamp 18001
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_312
timestamp 18001
transform 1 0 29808 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_388
timestamp 1636986456
transform 1 0 36800 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_400
timestamp 1636986456
transform 1 0 37904 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_412
timestamp 18001
transform 1 0 39008 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_421
timestamp 18001
transform 1 0 39836 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_425
timestamp 18001
transform 1 0 40204 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_3
timestamp 18001
transform 1 0 1380 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_11
timestamp 18001
transform 1 0 2116 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1636986456
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_39
timestamp 18001
transform 1 0 4692 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_43
timestamp 18001
transform 1 0 5060 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_69
timestamp 18001
transform 1 0 7452 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_77
timestamp 18001
transform 1 0 8188 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_82
timestamp 18001
transform 1 0 8648 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_96
timestamp 18001
transform 1 0 9936 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_103
timestamp 18001
transform 1 0 10580 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 18001
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1636986456
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1636986456
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_137
timestamp 18001
transform 1 0 13708 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_141
timestamp 18001
transform 1 0 14076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_151
timestamp 18001
transform 1 0 14996 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_159
timestamp 18001
transform 1 0 15732 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 18001
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_169
timestamp 18001
transform 1 0 16652 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_177
timestamp 18001
transform 1 0 17388 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_208
timestamp 1636986456
transform 1 0 20240 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_220
timestamp 18001
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 1636986456
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 1636986456
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_249
timestamp 1636986456
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_261
timestamp 1636986456
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_273
timestamp 18001
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 18001
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_320
timestamp 18001
transform 1 0 30544 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_337
timestamp 18001
transform 1 0 32108 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_349
timestamp 18001
transform 1 0 33212 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_365
timestamp 1636986456
transform 1 0 34684 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_377
timestamp 1636986456
transform 1 0 35788 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_389
timestamp 18001
transform 1 0 36892 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_393
timestamp 1636986456
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_405
timestamp 1636986456
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_417
timestamp 18001
transform 1 0 39468 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_425
timestamp 18001
transform 1 0 40204 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1636986456
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_15
timestamp 18001
transform 1 0 2484 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 18001
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1636986456
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1636986456
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1636986456
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1636986456
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_77
timestamp 18001
transform 1 0 8188 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_99
timestamp 18001
transform 1 0 10212 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_112
timestamp 18001
transform 1 0 11408 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_131
timestamp 18001
transform 1 0 13156 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 18001
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_141
timestamp 18001
transform 1 0 14076 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_166
timestamp 18001
transform 1 0 16376 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_172
timestamp 18001
transform 1 0 16928 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_183
timestamp 18001
transform 1 0 17940 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_194
timestamp 18001
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_197
timestamp 18001
transform 1 0 19228 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_205
timestamp 18001
transform 1 0 19964 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_213
timestamp 18001
transform 1 0 20700 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_221
timestamp 18001
transform 1 0 21436 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_230
timestamp 1636986456
transform 1 0 22264 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_242
timestamp 18001
transform 1 0 23368 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_250
timestamp 18001
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_262
timestamp 1636986456
transform 1 0 25208 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_274
timestamp 1636986456
transform 1 0 26312 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_306
timestamp 18001
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_309
timestamp 18001
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_332
timestamp 18001
transform 1 0 31648 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_336
timestamp 18001
transform 1 0 32016 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_357
timestamp 18001
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 18001
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 1636986456
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_377
timestamp 1636986456
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_389
timestamp 1636986456
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_401
timestamp 1636986456
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_413
timestamp 18001
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_419
timestamp 18001
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_421
timestamp 18001
transform 1 0 39836 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_425
timestamp 18001
transform 1 0 40204 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_3
timestamp 18001
transform 1 0 1380 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_11
timestamp 18001
transform 1 0 2116 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_36
timestamp 1636986456
transform 1 0 4416 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_48
timestamp 18001
transform 1 0 5520 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_65
timestamp 1636986456
transform 1 0 7084 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_77
timestamp 18001
transform 1 0 8188 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_81
timestamp 18001
transform 1 0 8556 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_85
timestamp 18001
transform 1 0 8924 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_91
timestamp 18001
transform 1 0 9476 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_95
timestamp 18001
transform 1 0 9844 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_99
timestamp 18001
transform 1 0 10212 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_113
timestamp 18001
transform 1 0 11500 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_139
timestamp 18001
transform 1 0 13892 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 1636986456
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 18001
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 18001
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_169
timestamp 18001
transform 1 0 16652 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_175
timestamp 18001
transform 1 0 17204 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_180
timestamp 18001
transform 1 0 17664 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_239
timestamp 18001
transform 1 0 23092 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_243
timestamp 18001
transform 1 0 23460 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_267
timestamp 1636986456
transform 1 0 25668 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 18001
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1636986456
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_293
timestamp 18001
transform 1 0 28060 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_304
timestamp 1636986456
transform 1 0 29072 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_323
timestamp 1636986456
transform 1 0 30820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 18001
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1636986456
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1636986456
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_361
timestamp 1636986456
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_373
timestamp 1636986456
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_385
timestamp 18001
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 18001
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_393
timestamp 1636986456
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_405
timestamp 1636986456
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_417
timestamp 18001
transform 1 0 39468 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_425
timestamp 18001
transform 1 0 40204 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_26
timestamp 18001
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_29
timestamp 18001
transform 1 0 3772 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_73
timestamp 18001
transform 1 0 7820 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_92
timestamp 1636986456
transform 1 0 9568 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_104
timestamp 1636986456
transform 1 0 10672 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_116
timestamp 18001
transform 1 0 11776 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_129
timestamp 18001
transform 1 0 12972 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_137
timestamp 18001
transform 1 0 13708 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1636986456
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_153
timestamp 18001
transform 1 0 15180 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_161
timestamp 18001
transform 1 0 15916 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_190
timestamp 18001
transform 1 0 18584 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_205
timestamp 18001
transform 1 0 19964 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_239
timestamp 1636986456
transform 1 0 23092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 18001
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 1636986456
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 1636986456
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_277
timestamp 1636986456
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_289
timestamp 1636986456
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_301
timestamp 18001
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 18001
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1636986456
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1636986456
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 1636986456
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 1636986456
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 18001
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 18001
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 1636986456
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 1636986456
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 1636986456
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_401
timestamp 1636986456
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_413
timestamp 18001
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_419
timestamp 18001
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_421
timestamp 18001
transform 1 0 39836 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_425
timestamp 18001
transform 1 0 40204 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_3
timestamp 18001
transform 1 0 1380 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_38
timestamp 1636986456
transform 1 0 4600 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_50
timestamp 18001
transform 1 0 5704 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_68
timestamp 18001
transform 1 0 7360 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_72
timestamp 18001
transform 1 0 7728 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_92
timestamp 18001
transform 1 0 9568 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_100
timestamp 18001
transform 1 0 10304 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_110
timestamp 18001
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_116
timestamp 18001
transform 1 0 11776 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_120
timestamp 1636986456
transform 1 0 12144 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_132
timestamp 18001
transform 1 0 13248 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_164
timestamp 18001
transform 1 0 16192 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_169
timestamp 18001
transform 1 0 16652 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_173
timestamp 18001
transform 1 0 17020 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_190
timestamp 18001
transform 1 0 18584 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_194
timestamp 18001
transform 1 0 18952 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_204
timestamp 1636986456
transform 1 0 19872 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_236
timestamp 18001
transform 1 0 22816 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_261
timestamp 18001
transform 1 0 25116 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_272
timestamp 18001
transform 1 0 26128 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1636986456
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1636986456
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 1636986456
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 1636986456
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 18001
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 18001
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1636986456
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1636986456
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_361
timestamp 1636986456
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_373
timestamp 1636986456
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_385
timestamp 18001
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 18001
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 1636986456
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_405
timestamp 1636986456
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_417
timestamp 18001
transform 1 0 39468 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_425
timestamp 18001
transform 1 0 40204 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1636986456
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1636986456
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 18001
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_35
timestamp 1636986456
transform 1 0 4324 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_47
timestamp 18001
transform 1 0 5428 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_51
timestamp 18001
transform 1 0 5796 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_61
timestamp 18001
transform 1 0 6716 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_80
timestamp 18001
transform 1 0 8464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_91
timestamp 18001
transform 1 0 9476 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_130
timestamp 18001
transform 1 0 13064 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_138
timestamp 18001
transform 1 0 13800 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_155
timestamp 18001
transform 1 0 15364 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_161
timestamp 1636986456
transform 1 0 15916 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_173
timestamp 1636986456
transform 1 0 17020 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_188
timestamp 18001
transform 1 0 18400 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_197
timestamp 18001
transform 1 0 19228 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_229
timestamp 18001
transform 1 0 22172 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_233
timestamp 18001
transform 1 0 22540 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_253
timestamp 18001
transform 1 0 24380 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_284
timestamp 1636986456
transform 1 0 27232 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_296
timestamp 1636986456
transform 1 0 28336 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1636986456
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1636986456
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_333
timestamp 1636986456
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_345
timestamp 1636986456
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_357
timestamp 18001
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 18001
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 1636986456
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 1636986456
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 1636986456
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_401
timestamp 1636986456
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_413
timestamp 18001
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_419
timestamp 18001
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_421
timestamp 18001
transform 1 0 39836 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_425
timestamp 18001
transform 1 0 40204 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1636986456
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1636986456
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1636986456
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_39
timestamp 18001
transform 1 0 4692 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_47
timestamp 18001
transform 1 0 5428 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_54
timestamp 18001
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_60
timestamp 1636986456
transform 1 0 6624 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_72
timestamp 18001
transform 1 0 7728 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_84
timestamp 1636986456
transform 1 0 8832 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_96
timestamp 18001
transform 1 0 9936 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_109
timestamp 18001
transform 1 0 11132 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_113
timestamp 18001
transform 1 0 11500 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_125
timestamp 18001
transform 1 0 12604 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_150
timestamp 18001
transform 1 0 14904 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_166
timestamp 18001
transform 1 0 16376 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_169
timestamp 18001
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_175
timestamp 18001
transform 1 0 17204 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_181
timestamp 18001
transform 1 0 17756 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_187
timestamp 18001
transform 1 0 18308 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_195
timestamp 1636986456
transform 1 0 19044 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_207
timestamp 1636986456
transform 1 0 20148 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_219
timestamp 18001
transform 1 0 21252 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 18001
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_225
timestamp 18001
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_233
timestamp 18001
transform 1 0 22540 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_247
timestamp 18001
transform 1 0 23828 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_255
timestamp 18001
transform 1 0 24564 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_281
timestamp 1636986456
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_293
timestamp 1636986456
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_305
timestamp 1636986456
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_317
timestamp 1636986456
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 18001
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 18001
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 1636986456
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_349
timestamp 1636986456
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_361
timestamp 1636986456
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_373
timestamp 1636986456
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_385
timestamp 18001
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 18001
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_393
timestamp 1636986456
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_405
timestamp 1636986456
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_417
timestamp 18001
transform 1 0 39468 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_425
timestamp 18001
transform 1 0 40204 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1636986456
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1636986456
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 18001
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1636986456
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_41
timestamp 18001
transform 1 0 4876 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_59
timestamp 1636986456
transform 1 0 6532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_71
timestamp 18001
transform 1 0 7636 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_75
timestamp 18001
transform 1 0 8004 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_82
timestamp 18001
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_91
timestamp 1636986456
transform 1 0 9476 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_103
timestamp 1636986456
transform 1 0 10580 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_115
timestamp 18001
transform 1 0 11684 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_128
timestamp 1636986456
transform 1 0 12880 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_141
timestamp 18001
transform 1 0 14076 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_174
timestamp 18001
transform 1 0 17112 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_185
timestamp 18001
transform 1 0 18124 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_193
timestamp 18001
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_203
timestamp 18001
transform 1 0 19780 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_209
timestamp 18001
transform 1 0 20332 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_217
timestamp 18001
transform 1 0 21068 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_225
timestamp 1636986456
transform 1 0 21804 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_237
timestamp 18001
transform 1 0 22908 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_247
timestamp 18001
transform 1 0 23828 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_251
timestamp 18001
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_253
timestamp 18001
transform 1 0 24380 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_261
timestamp 18001
transform 1 0 25116 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_273
timestamp 1636986456
transform 1 0 26220 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_285
timestamp 1636986456
transform 1 0 27324 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_297
timestamp 18001
transform 1 0 28428 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_305
timestamp 18001
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 1636986456
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 1636986456
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_333
timestamp 1636986456
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_345
timestamp 1636986456
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_357
timestamp 18001
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_363
timestamp 18001
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 1636986456
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 1636986456
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_389
timestamp 1636986456
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_401
timestamp 1636986456
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_413
timestamp 18001
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_419
timestamp 18001
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_421
timestamp 18001
transform 1 0 39836 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_425
timestamp 18001
transform 1 0 40204 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1636986456
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 1636986456
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_27
timestamp 18001
transform 1 0 3588 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_78
timestamp 18001
transform 1 0 8280 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_93
timestamp 1636986456
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_105
timestamp 18001
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_111
timestamp 18001
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_113
timestamp 1636986456
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_125
timestamp 18001
transform 1 0 12604 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_165
timestamp 18001
transform 1 0 16284 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_169
timestamp 18001
transform 1 0 16652 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_177
timestamp 18001
transform 1 0 17388 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_185
timestamp 18001
transform 1 0 18124 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_191
timestamp 18001
transform 1 0 18676 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_229
timestamp 18001
transform 1 0 22172 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_254
timestamp 18001
transform 1 0 24472 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_258
timestamp 18001
transform 1 0 24840 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_268
timestamp 1636986456
transform 1 0 25760 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_281
timestamp 1636986456
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_293
timestamp 1636986456
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_305
timestamp 1636986456
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_317
timestamp 1636986456
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_329
timestamp 18001
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_335
timestamp 18001
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_337
timestamp 1636986456
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_349
timestamp 1636986456
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_361
timestamp 1636986456
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_373
timestamp 1636986456
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_385
timestamp 18001
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_391
timestamp 18001
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_393
timestamp 1636986456
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_405
timestamp 1636986456
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_417
timestamp 18001
transform 1 0 39468 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_425
timestamp 18001
transform 1 0 40204 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 1636986456
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 1636986456
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 18001
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1636986456
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_41
timestamp 18001
transform 1 0 4876 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_51
timestamp 1636986456
transform 1 0 5796 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_63
timestamp 18001
transform 1 0 6900 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_71
timestamp 18001
transform 1 0 7636 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_91
timestamp 18001
transform 1 0 9476 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_97
timestamp 18001
transform 1 0 10028 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_103
timestamp 18001
transform 1 0 10580 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_114
timestamp 18001
transform 1 0 11592 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_122
timestamp 18001
transform 1 0 12328 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_134
timestamp 18001
transform 1 0 13432 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 1636986456
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_153
timestamp 1636986456
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_165
timestamp 1636986456
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_177
timestamp 18001
transform 1 0 17388 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_190
timestamp 18001
transform 1 0 18584 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_197
timestamp 1636986456
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_209
timestamp 18001
transform 1 0 20332 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_218
timestamp 18001
transform 1 0 21160 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_225
timestamp 1636986456
transform 1 0 21804 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_249
timestamp 18001
transform 1 0 24012 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_253
timestamp 18001
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_301
timestamp 18001
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_307
timestamp 18001
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_309
timestamp 1636986456
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_321
timestamp 1636986456
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_333
timestamp 1636986456
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_345
timestamp 1636986456
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_357
timestamp 18001
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_363
timestamp 18001
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_365
timestamp 1636986456
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_377
timestamp 1636986456
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_389
timestamp 1636986456
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_401
timestamp 1636986456
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_413
timestamp 18001
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_419
timestamp 18001
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_421
timestamp 18001
transform 1 0 39836 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_425
timestamp 18001
transform 1 0 40204 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_3
timestamp 1636986456
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_15
timestamp 1636986456
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_27
timestamp 1636986456
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_39
timestamp 1636986456
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_51
timestamp 18001
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 18001
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1636986456
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_69
timestamp 18001
transform 1 0 7452 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_77
timestamp 18001
transform 1 0 8188 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_102
timestamp 18001
transform 1 0 10488 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_110
timestamp 18001
transform 1 0 11224 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_124
timestamp 1636986456
transform 1 0 12512 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_136
timestamp 1636986456
transform 1 0 13616 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_148
timestamp 1636986456
transform 1 0 14720 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_160
timestamp 18001
transform 1 0 15824 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_173
timestamp 18001
transform 1 0 17020 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_181
timestamp 18001
transform 1 0 17756 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_207
timestamp 1636986456
transform 1 0 20148 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_219
timestamp 18001
transform 1 0 21252 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_223
timestamp 18001
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_225
timestamp 18001
transform 1 0 21804 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_233
timestamp 18001
transform 1 0 22540 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_257
timestamp 18001
transform 1 0 24748 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_263
timestamp 18001
transform 1 0 25300 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_273
timestamp 18001
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_279
timestamp 18001
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_281
timestamp 1636986456
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_293
timestamp 1636986456
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_305
timestamp 1636986456
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_317
timestamp 1636986456
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_329
timestamp 18001
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_335
timestamp 18001
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_337
timestamp 1636986456
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_349
timestamp 1636986456
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_361
timestamp 1636986456
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_373
timestamp 1636986456
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_385
timestamp 18001
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_391
timestamp 18001
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_393
timestamp 1636986456
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_405
timestamp 1636986456
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_417
timestamp 18001
transform 1 0 39468 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_425
timestamp 18001
transform 1 0 40204 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_3
timestamp 1636986456
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_15
timestamp 1636986456
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 18001
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_29
timestamp 1636986456
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_41
timestamp 1636986456
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_53
timestamp 1636986456
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_65
timestamp 1636986456
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_77
timestamp 18001
transform 1 0 8188 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_85
timestamp 1636986456
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_97
timestamp 1636986456
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_109
timestamp 18001
transform 1 0 11132 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_116
timestamp 18001
transform 1 0 11776 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_130
timestamp 18001
transform 1 0 13064 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_138
timestamp 18001
transform 1 0 13800 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_141
timestamp 18001
transform 1 0 14076 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_148
timestamp 18001
transform 1 0 14720 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_156
timestamp 18001
transform 1 0 15456 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_169
timestamp 18001
transform 1 0 16652 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_186
timestamp 18001
transform 1 0 18216 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_194
timestamp 18001
transform 1 0 18952 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_197
timestamp 1636986456
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_209
timestamp 1636986456
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_221
timestamp 1636986456
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_233
timestamp 1636986456
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_245
timestamp 18001
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_251
timestamp 18001
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_253
timestamp 1636986456
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_265
timestamp 1636986456
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_277
timestamp 1636986456
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_289
timestamp 1636986456
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_301
timestamp 18001
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_307
timestamp 18001
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_309
timestamp 1636986456
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_321
timestamp 1636986456
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_333
timestamp 1636986456
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_345
timestamp 1636986456
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_357
timestamp 18001
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_363
timestamp 18001
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_365
timestamp 1636986456
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_377
timestamp 1636986456
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_389
timestamp 1636986456
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_401
timestamp 1636986456
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_413
timestamp 18001
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_419
timestamp 18001
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_421
timestamp 18001
transform 1 0 39836 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_425
timestamp 18001
transform 1 0 40204 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_3
timestamp 1636986456
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_15
timestamp 1636986456
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_27
timestamp 1636986456
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_39
timestamp 1636986456
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_51
timestamp 18001
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_55
timestamp 18001
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_57
timestamp 1636986456
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_69
timestamp 1636986456
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_81
timestamp 1636986456
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_93
timestamp 1636986456
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_105
timestamp 18001
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_111
timestamp 18001
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_113
timestamp 18001
transform 1 0 11500 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_123
timestamp 18001
transform 1 0 12420 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_131
timestamp 18001
transform 1 0 13156 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_174
timestamp 1636986456
transform 1 0 17112 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_186
timestamp 1636986456
transform 1 0 18216 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_198
timestamp 1636986456
transform 1 0 19320 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_210
timestamp 1636986456
transform 1 0 20424 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_222
timestamp 18001
transform 1 0 21528 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_225
timestamp 1636986456
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_237
timestamp 1636986456
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_249
timestamp 1636986456
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_261
timestamp 1636986456
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_273
timestamp 18001
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_279
timestamp 18001
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_281
timestamp 1636986456
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_293
timestamp 1636986456
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_305
timestamp 1636986456
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_317
timestamp 1636986456
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_329
timestamp 18001
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_335
timestamp 18001
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_337
timestamp 1636986456
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_349
timestamp 1636986456
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_361
timestamp 1636986456
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_373
timestamp 1636986456
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_385
timestamp 18001
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_391
timestamp 18001
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_393
timestamp 1636986456
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_405
timestamp 1636986456
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_417
timestamp 18001
transform 1 0 39468 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_425
timestamp 18001
transform 1 0 40204 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_3
timestamp 1636986456
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_15
timestamp 1636986456
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_27
timestamp 18001
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_29
timestamp 1636986456
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_41
timestamp 1636986456
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_53
timestamp 1636986456
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_65
timestamp 1636986456
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_77
timestamp 18001
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 18001
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_85
timestamp 1636986456
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_97
timestamp 1636986456
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_109
timestamp 1636986456
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_121
timestamp 1636986456
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_133
timestamp 18001
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_139
timestamp 18001
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_141
timestamp 1636986456
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_153
timestamp 18001
transform 1 0 15180 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_169
timestamp 1636986456
transform 1 0 16652 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_181
timestamp 1636986456
transform 1 0 17756 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_193
timestamp 18001
transform 1 0 18860 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_197
timestamp 1636986456
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_209
timestamp 1636986456
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_221
timestamp 1636986456
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_233
timestamp 1636986456
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_245
timestamp 18001
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_251
timestamp 18001
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_253
timestamp 1636986456
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_265
timestamp 1636986456
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_277
timestamp 1636986456
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_289
timestamp 1636986456
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_301
timestamp 18001
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_307
timestamp 18001
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_309
timestamp 1636986456
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_321
timestamp 1636986456
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_333
timestamp 1636986456
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_345
timestamp 1636986456
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_357
timestamp 18001
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_363
timestamp 18001
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_365
timestamp 1636986456
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_377
timestamp 1636986456
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_389
timestamp 1636986456
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_401
timestamp 1636986456
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_413
timestamp 18001
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_419
timestamp 18001
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_421
timestamp 18001
transform 1 0 39836 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_425
timestamp 18001
transform 1 0 40204 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_3
timestamp 1636986456
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_15
timestamp 1636986456
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_27
timestamp 18001
transform 1 0 3588 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_29
timestamp 1636986456
transform 1 0 3772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_41
timestamp 1636986456
transform 1 0 4876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_53
timestamp 18001
transform 1 0 5980 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 1636986456
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_69
timestamp 1636986456
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_81
timestamp 18001
transform 1 0 8556 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_85
timestamp 1636986456
transform 1 0 8924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_97
timestamp 1636986456
transform 1 0 10028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_109
timestamp 18001
transform 1 0 11132 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_113
timestamp 1636986456
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_125
timestamp 1636986456
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_137
timestamp 18001
transform 1 0 13708 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_141
timestamp 1636986456
transform 1 0 14076 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_153
timestamp 1636986456
transform 1 0 15180 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_165
timestamp 18001
transform 1 0 16284 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_169
timestamp 1636986456
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_181
timestamp 1636986456
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_193
timestamp 18001
transform 1 0 18860 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_197
timestamp 1636986456
transform 1 0 19228 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_209
timestamp 1636986456
transform 1 0 20332 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_221
timestamp 18001
transform 1 0 21436 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_225
timestamp 1636986456
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_237
timestamp 1636986456
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_249
timestamp 18001
transform 1 0 24012 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_253
timestamp 1636986456
transform 1 0 24380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_265
timestamp 1636986456
transform 1 0 25484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_277
timestamp 18001
transform 1 0 26588 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_281
timestamp 1636986456
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_293
timestamp 1636986456
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_305
timestamp 18001
transform 1 0 29164 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_309
timestamp 1636986456
transform 1 0 29532 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_321
timestamp 18001
transform 1 0 30636 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_331
timestamp 18001
transform 1 0 31556 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_335
timestamp 18001
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_337
timestamp 1636986456
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_349
timestamp 1636986456
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_361
timestamp 18001
transform 1 0 34316 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_365
timestamp 1636986456
transform 1 0 34684 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_377
timestamp 1636986456
transform 1 0 35788 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_389
timestamp 18001
transform 1 0 36892 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_393
timestamp 1636986456
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_405
timestamp 1636986456
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_417
timestamp 18001
transform 1 0 39468 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_421
timestamp 18001
transform 1 0 39836 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_425
timestamp 18001
transform 1 0 40204 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 18001
transform 1 0 19964 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 18001
transform -1 0 18124 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 18001
transform -1 0 34224 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 18001
transform -1 0 21896 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 18001
transform -1 0 18676 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 18001
transform -1 0 22356 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 18001
transform -1 0 22540 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 18001
transform 1 0 21988 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 18001
transform 1 0 24564 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 18001
transform -1 0 26956 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 18001
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 18001
transform 1 0 19320 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 18001
transform -1 0 12328 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 18001
transform -1 0 14076 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 18001
transform -1 0 9384 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 18001
transform -1 0 11316 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 18001
transform -1 0 4508 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 18001
transform -1 0 8832 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 18001
transform -1 0 5888 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 18001
transform -1 0 11132 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 18001
transform -1 0 5980 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 18001
transform -1 0 13524 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 18001
transform -1 0 7912 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 18001
transform -1 0 15916 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 18001
transform -1 0 5612 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 18001
transform -1 0 19780 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 18001
transform -1 0 14812 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 18001
transform -1 0 16192 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 18001
transform -1 0 17848 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 18001
transform -1 0 3680 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 18001
transform 1 0 28796 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 18001
transform -1 0 13892 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 18001
transform -1 0 5244 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 18001
transform -1 0 5336 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 18001
transform -1 0 13064 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 18001
transform -1 0 6072 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 18001
transform -1 0 5060 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 18001
transform -1 0 32844 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 18001
transform -1 0 13432 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 18001
transform -1 0 6256 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 18001
transform -1 0 9660 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 18001
transform 1 0 28336 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 18001
transform -1 0 14720 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 18001
transform -1 0 19504 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 18001
transform -1 0 4140 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 18001
transform -1 0 4508 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 18001
transform -1 0 6348 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 18001
transform 1 0 9384 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 18001
transform 1 0 34776 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 18001
transform -1 0 4508 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 18001
transform -1 0 31464 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 18001
transform -1 0 9384 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 18001
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 18001
transform 1 0 29532 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 18001
transform -1 0 39744 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input2
timestamp 18001
transform 1 0 31004 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 18001
transform -1 0 40296 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 18001
transform 1 0 1380 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 18001
transform -1 0 40296 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 18001
transform 1 0 39376 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input7
timestamp 18001
transform -1 0 39744 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 18001
transform -1 0 40296 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 18001
transform -1 0 40296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 18001
transform -1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 18001
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 18001
transform 1 0 14260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 18001
transform -1 0 11408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 18001
transform 1 0 15272 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 18001
transform -1 0 13708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 18001
transform 1 0 11592 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 18001
transform -1 0 15272 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 18001
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_72
timestamp 18001
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 18001
transform -1 0 40572 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_73
timestamp 18001
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 18001
transform -1 0 40572 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_74
timestamp 18001
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 18001
transform -1 0 40572 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_75
timestamp 18001
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 18001
transform -1 0 40572 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_76
timestamp 18001
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 18001
transform -1 0 40572 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_77
timestamp 18001
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 18001
transform -1 0 40572 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_78
timestamp 18001
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 18001
transform -1 0 40572 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_79
timestamp 18001
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 18001
transform -1 0 40572 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_80
timestamp 18001
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 18001
transform -1 0 40572 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_81
timestamp 18001
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 18001
transform -1 0 40572 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_82
timestamp 18001
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 18001
transform -1 0 40572 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_83
timestamp 18001
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 18001
transform -1 0 40572 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_84
timestamp 18001
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 18001
transform -1 0 40572 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_85
timestamp 18001
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 18001
transform -1 0 40572 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_86
timestamp 18001
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 18001
transform -1 0 40572 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_87
timestamp 18001
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 18001
transform -1 0 40572 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_88
timestamp 18001
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 18001
transform -1 0 40572 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_89
timestamp 18001
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 18001
transform -1 0 40572 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_90
timestamp 18001
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 18001
transform -1 0 40572 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_91
timestamp 18001
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 18001
transform -1 0 40572 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_92
timestamp 18001
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 18001
transform -1 0 40572 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_93
timestamp 18001
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 18001
transform -1 0 40572 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_94
timestamp 18001
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 18001
transform -1 0 40572 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_95
timestamp 18001
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 18001
transform -1 0 40572 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_96
timestamp 18001
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 18001
transform -1 0 40572 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_97
timestamp 18001
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 18001
transform -1 0 40572 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_98
timestamp 18001
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 18001
transform -1 0 40572 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_99
timestamp 18001
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 18001
transform -1 0 40572 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_100
timestamp 18001
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 18001
transform -1 0 40572 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_101
timestamp 18001
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 18001
transform -1 0 40572 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_102
timestamp 18001
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 18001
transform -1 0 40572 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_103
timestamp 18001
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 18001
transform -1 0 40572 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_104
timestamp 18001
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 18001
transform -1 0 40572 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_105
timestamp 18001
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 18001
transform -1 0 40572 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_106
timestamp 18001
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 18001
transform -1 0 40572 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_107
timestamp 18001
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 18001
transform -1 0 40572 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_108
timestamp 18001
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 18001
transform -1 0 40572 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_109
timestamp 18001
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 18001
transform -1 0 40572 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_110
timestamp 18001
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 18001
transform -1 0 40572 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_111
timestamp 18001
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 18001
transform -1 0 40572 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_112
timestamp 18001
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 18001
transform -1 0 40572 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_113
timestamp 18001
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 18001
transform -1 0 40572 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_114
timestamp 18001
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 18001
transform -1 0 40572 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_115
timestamp 18001
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 18001
transform -1 0 40572 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_116
timestamp 18001
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 18001
transform -1 0 40572 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_117
timestamp 18001
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 18001
transform -1 0 40572 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_118
timestamp 18001
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 18001
transform -1 0 40572 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_119
timestamp 18001
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 18001
transform -1 0 40572 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_120
timestamp 18001
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 18001
transform -1 0 40572 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_121
timestamp 18001
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 18001
transform -1 0 40572 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_122
timestamp 18001
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 18001
transform -1 0 40572 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_123
timestamp 18001
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 18001
transform -1 0 40572 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_124
timestamp 18001
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 18001
transform -1 0 40572 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_125
timestamp 18001
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 18001
transform -1 0 40572 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_126
timestamp 18001
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 18001
transform -1 0 40572 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_127
timestamp 18001
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 18001
transform -1 0 40572 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_128
timestamp 18001
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 18001
transform -1 0 40572 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_129
timestamp 18001
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 18001
transform -1 0 40572 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_130
timestamp 18001
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 18001
transform -1 0 40572 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_131
timestamp 18001
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 18001
transform -1 0 40572 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_132
timestamp 18001
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 18001
transform -1 0 40572 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_133
timestamp 18001
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 18001
transform -1 0 40572 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_134
timestamp 18001
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 18001
transform -1 0 40572 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_135
timestamp 18001
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 18001
transform -1 0 40572 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_136
timestamp 18001
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 18001
transform -1 0 40572 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_137
timestamp 18001
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp 18001
transform -1 0 40572 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Left_138
timestamp 18001
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Right_66
timestamp 18001
transform -1 0 40572 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_139
timestamp 18001
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_67
timestamp 18001
transform -1 0 40572 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_140
timestamp 18001
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_68
timestamp 18001
transform -1 0 40572 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_141
timestamp 18001
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_69
timestamp 18001
transform -1 0 40572 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_142
timestamp 18001
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_70
timestamp 18001
transform -1 0 40572 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_143
timestamp 18001
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_71
timestamp 18001
transform -1 0 40572 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_144
timestamp 18001
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_145
timestamp 18001
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_146
timestamp 18001
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_147
timestamp 18001
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_148
timestamp 18001
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_149
timestamp 18001
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_150
timestamp 18001
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_151
timestamp 18001
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_152
timestamp 18001
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_153
timestamp 18001
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_154
timestamp 18001
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_155
timestamp 18001
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_156
timestamp 18001
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_157
timestamp 18001
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_158
timestamp 18001
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_159
timestamp 18001
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_160
timestamp 18001
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_161
timestamp 18001
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_162
timestamp 18001
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_163
timestamp 18001
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_164
timestamp 18001
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_165
timestamp 18001
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_166
timestamp 18001
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_167
timestamp 18001
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_168
timestamp 18001
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_169
timestamp 18001
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_170
timestamp 18001
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_171
timestamp 18001
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_172
timestamp 18001
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_173
timestamp 18001
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_174
timestamp 18001
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_175
timestamp 18001
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_176
timestamp 18001
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_177
timestamp 18001
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_178
timestamp 18001
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_179
timestamp 18001
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_180
timestamp 18001
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_181
timestamp 18001
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_182
timestamp 18001
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_183
timestamp 18001
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_184
timestamp 18001
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_185
timestamp 18001
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_186
timestamp 18001
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_187
timestamp 18001
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_188
timestamp 18001
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_189
timestamp 18001
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_190
timestamp 18001
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_191
timestamp 18001
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_192
timestamp 18001
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_193
timestamp 18001
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_194
timestamp 18001
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_195
timestamp 18001
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_196
timestamp 18001
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_197
timestamp 18001
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_198
timestamp 18001
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_199
timestamp 18001
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_200
timestamp 18001
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_201
timestamp 18001
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_202
timestamp 18001
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_203
timestamp 18001
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_204
timestamp 18001
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_205
timestamp 18001
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_206
timestamp 18001
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_207
timestamp 18001
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_208
timestamp 18001
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_209
timestamp 18001
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_210
timestamp 18001
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_211
timestamp 18001
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_212
timestamp 18001
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_213
timestamp 18001
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_214
timestamp 18001
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_215
timestamp 18001
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_216
timestamp 18001
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_217
timestamp 18001
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_218
timestamp 18001
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_219
timestamp 18001
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_220
timestamp 18001
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_221
timestamp 18001
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_222
timestamp 18001
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_223
timestamp 18001
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_224
timestamp 18001
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_225
timestamp 18001
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_226
timestamp 18001
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_227
timestamp 18001
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_228
timestamp 18001
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_229
timestamp 18001
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_230
timestamp 18001
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_231
timestamp 18001
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_232
timestamp 18001
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_233
timestamp 18001
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_234
timestamp 18001
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_235
timestamp 18001
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_236
timestamp 18001
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_237
timestamp 18001
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_238
timestamp 18001
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_239
timestamp 18001
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_240
timestamp 18001
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_241
timestamp 18001
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_242
timestamp 18001
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_243
timestamp 18001
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_244
timestamp 18001
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_245
timestamp 18001
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_246
timestamp 18001
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_247
timestamp 18001
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_248
timestamp 18001
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_249
timestamp 18001
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_250
timestamp 18001
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_251
timestamp 18001
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_252
timestamp 18001
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_253
timestamp 18001
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_254
timestamp 18001
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_255
timestamp 18001
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_256
timestamp 18001
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_257
timestamp 18001
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_258
timestamp 18001
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_259
timestamp 18001
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_260
timestamp 18001
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_261
timestamp 18001
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_262
timestamp 18001
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_263
timestamp 18001
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_264
timestamp 18001
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_265
timestamp 18001
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_266
timestamp 18001
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_267
timestamp 18001
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_268
timestamp 18001
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_269
timestamp 18001
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_270
timestamp 18001
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_271
timestamp 18001
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_272
timestamp 18001
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_273
timestamp 18001
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_274
timestamp 18001
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_275
timestamp 18001
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_276
timestamp 18001
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_277
timestamp 18001
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_278
timestamp 18001
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_279
timestamp 18001
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_280
timestamp 18001
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_281
timestamp 18001
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_282
timestamp 18001
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_283
timestamp 18001
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_284
timestamp 18001
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_285
timestamp 18001
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_286
timestamp 18001
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_287
timestamp 18001
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_288
timestamp 18001
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_289
timestamp 18001
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_290
timestamp 18001
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_291
timestamp 18001
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_292
timestamp 18001
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_293
timestamp 18001
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_294
timestamp 18001
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_295
timestamp 18001
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_296
timestamp 18001
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_297
timestamp 18001
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_298
timestamp 18001
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_299
timestamp 18001
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_300
timestamp 18001
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_301
timestamp 18001
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_302
timestamp 18001
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_303
timestamp 18001
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_304
timestamp 18001
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_305
timestamp 18001
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_306
timestamp 18001
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_307
timestamp 18001
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_308
timestamp 18001
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_309
timestamp 18001
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_310
timestamp 18001
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_311
timestamp 18001
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_312
timestamp 18001
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_313
timestamp 18001
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_314
timestamp 18001
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_315
timestamp 18001
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_316
timestamp 18001
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_317
timestamp 18001
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_318
timestamp 18001
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_319
timestamp 18001
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_320
timestamp 18001
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_321
timestamp 18001
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_322
timestamp 18001
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_323
timestamp 18001
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_324
timestamp 18001
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_325
timestamp 18001
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_326
timestamp 18001
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_327
timestamp 18001
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_328
timestamp 18001
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_329
timestamp 18001
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_330
timestamp 18001
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_331
timestamp 18001
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_332
timestamp 18001
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_333
timestamp 18001
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_334
timestamp 18001
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_335
timestamp 18001
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_336
timestamp 18001
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_337
timestamp 18001
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_338
timestamp 18001
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_339
timestamp 18001
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_340
timestamp 18001
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_341
timestamp 18001
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_342
timestamp 18001
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_343
timestamp 18001
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_344
timestamp 18001
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_345
timestamp 18001
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_346
timestamp 18001
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_347
timestamp 18001
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_348
timestamp 18001
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_349
timestamp 18001
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_350
timestamp 18001
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_351
timestamp 18001
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_352
timestamp 18001
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_353
timestamp 18001
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_354
timestamp 18001
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_355
timestamp 18001
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_356
timestamp 18001
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_357
timestamp 18001
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_358
timestamp 18001
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_359
timestamp 18001
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_360
timestamp 18001
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_361
timestamp 18001
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_362
timestamp 18001
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_363
timestamp 18001
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_364
timestamp 18001
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_365
timestamp 18001
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_366
timestamp 18001
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_367
timestamp 18001
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_368
timestamp 18001
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_369
timestamp 18001
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_370
timestamp 18001
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_371
timestamp 18001
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_372
timestamp 18001
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_373
timestamp 18001
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_374
timestamp 18001
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_375
timestamp 18001
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_376
timestamp 18001
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_377
timestamp 18001
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_378
timestamp 18001
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_379
timestamp 18001
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_380
timestamp 18001
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_381
timestamp 18001
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_382
timestamp 18001
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_383
timestamp 18001
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_384
timestamp 18001
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_385
timestamp 18001
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_386
timestamp 18001
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_387
timestamp 18001
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_388
timestamp 18001
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_389
timestamp 18001
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_390
timestamp 18001
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_391
timestamp 18001
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_392
timestamp 18001
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_393
timestamp 18001
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_394
timestamp 18001
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_395
timestamp 18001
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_396
timestamp 18001
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_397
timestamp 18001
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_398
timestamp 18001
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_399
timestamp 18001
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_400
timestamp 18001
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_401
timestamp 18001
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_402
timestamp 18001
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_403
timestamp 18001
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_404
timestamp 18001
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_405
timestamp 18001
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_406
timestamp 18001
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_407
timestamp 18001
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_408
timestamp 18001
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_409
timestamp 18001
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_410
timestamp 18001
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_411
timestamp 18001
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_412
timestamp 18001
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_413
timestamp 18001
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_414
timestamp 18001
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_415
timestamp 18001
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_416
timestamp 18001
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_417
timestamp 18001
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_418
timestamp 18001
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_419
timestamp 18001
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_420
timestamp 18001
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_421
timestamp 18001
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_422
timestamp 18001
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_423
timestamp 18001
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_424
timestamp 18001
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_425
timestamp 18001
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_426
timestamp 18001
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_427
timestamp 18001
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_428
timestamp 18001
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_429
timestamp 18001
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_430
timestamp 18001
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_431
timestamp 18001
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_432
timestamp 18001
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_433
timestamp 18001
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_434
timestamp 18001
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_435
timestamp 18001
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_436
timestamp 18001
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_437
timestamp 18001
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_438
timestamp 18001
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_439
timestamp 18001
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_440
timestamp 18001
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_441
timestamp 18001
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_442
timestamp 18001
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_443
timestamp 18001
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_444
timestamp 18001
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_445
timestamp 18001
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_446
timestamp 18001
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_447
timestamp 18001
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_448
timestamp 18001
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_449
timestamp 18001
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_450
timestamp 18001
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_451
timestamp 18001
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_452
timestamp 18001
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_453
timestamp 18001
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_454
timestamp 18001
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_455
timestamp 18001
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_456
timestamp 18001
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_457
timestamp 18001
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_458
timestamp 18001
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_459
timestamp 18001
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_460
timestamp 18001
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_461
timestamp 18001
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_462
timestamp 18001
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_463
timestamp 18001
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_464
timestamp 18001
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_465
timestamp 18001
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_466
timestamp 18001
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_467
timestamp 18001
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_468
timestamp 18001
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_469
timestamp 18001
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_470
timestamp 18001
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_471
timestamp 18001
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_472
timestamp 18001
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_473
timestamp 18001
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_474
timestamp 18001
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_475
timestamp 18001
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_476
timestamp 18001
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_477
timestamp 18001
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_478
timestamp 18001
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_479
timestamp 18001
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_480
timestamp 18001
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_481
timestamp 18001
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_482
timestamp 18001
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_483
timestamp 18001
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_484
timestamp 18001
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_485
timestamp 18001
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_486
timestamp 18001
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_487
timestamp 18001
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_488
timestamp 18001
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_489
timestamp 18001
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_490
timestamp 18001
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_491
timestamp 18001
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_492
timestamp 18001
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_493
timestamp 18001
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_494
timestamp 18001
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_495
timestamp 18001
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_496
timestamp 18001
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_497
timestamp 18001
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_498
timestamp 18001
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_499
timestamp 18001
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_500
timestamp 18001
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_501
timestamp 18001
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_502
timestamp 18001
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_503
timestamp 18001
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_504
timestamp 18001
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_505
timestamp 18001
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_506
timestamp 18001
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_507
timestamp 18001
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_508
timestamp 18001
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_509
timestamp 18001
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_510
timestamp 18001
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_511
timestamp 18001
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_512
timestamp 18001
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_513
timestamp 18001
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_514
timestamp 18001
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_515
timestamp 18001
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_516
timestamp 18001
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_517
timestamp 18001
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_518
timestamp 18001
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_519
timestamp 18001
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_520
timestamp 18001
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_521
timestamp 18001
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_522
timestamp 18001
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_523
timestamp 18001
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_524
timestamp 18001
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_525
timestamp 18001
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_526
timestamp 18001
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_527
timestamp 18001
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_528
timestamp 18001
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_529
timestamp 18001
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_530
timestamp 18001
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_531
timestamp 18001
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_532
timestamp 18001
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_533
timestamp 18001
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_534
timestamp 18001
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_535
timestamp 18001
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_536
timestamp 18001
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_537
timestamp 18001
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_538
timestamp 18001
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_539
timestamp 18001
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_540
timestamp 18001
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_541
timestamp 18001
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_542
timestamp 18001
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_543
timestamp 18001
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_544
timestamp 18001
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_545
timestamp 18001
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_546
timestamp 18001
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_547
timestamp 18001
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_548
timestamp 18001
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_549
timestamp 18001
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_550
timestamp 18001
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_551
timestamp 18001
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_552
timestamp 18001
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_553
timestamp 18001
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_554
timestamp 18001
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_555
timestamp 18001
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_556
timestamp 18001
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_557
timestamp 18001
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_558
timestamp 18001
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_559
timestamp 18001
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_560
timestamp 18001
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_561
timestamp 18001
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_562
timestamp 18001
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_563
timestamp 18001
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_564
timestamp 18001
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_565
timestamp 18001
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_566
timestamp 18001
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_567
timestamp 18001
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_568
timestamp 18001
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_569
timestamp 18001
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_570
timestamp 18001
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_571
timestamp 18001
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_572
timestamp 18001
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_573
timestamp 18001
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_574
timestamp 18001
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_575
timestamp 18001
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_576
timestamp 18001
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_577
timestamp 18001
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_578
timestamp 18001
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_579
timestamp 18001
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_580
timestamp 18001
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_581
timestamp 18001
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_582
timestamp 18001
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_583
timestamp 18001
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_584
timestamp 18001
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_585
timestamp 18001
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_586
timestamp 18001
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_587
timestamp 18001
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_588
timestamp 18001
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_589
timestamp 18001
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_590
timestamp 18001
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_591
timestamp 18001
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_592
timestamp 18001
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_593
timestamp 18001
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_594
timestamp 18001
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_595
timestamp 18001
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_596
timestamp 18001
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_597
timestamp 18001
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_598
timestamp 18001
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_599
timestamp 18001
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_600
timestamp 18001
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_601
timestamp 18001
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_602
timestamp 18001
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_603
timestamp 18001
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_604
timestamp 18001
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_605
timestamp 18001
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_606
timestamp 18001
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_607
timestamp 18001
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_608
timestamp 18001
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_609
timestamp 18001
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_610
timestamp 18001
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_611
timestamp 18001
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_612
timestamp 18001
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_613
timestamp 18001
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_614
timestamp 18001
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_615
timestamp 18001
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_616
timestamp 18001
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_617
timestamp 18001
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_618
timestamp 18001
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_619
timestamp 18001
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_620
timestamp 18001
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_621
timestamp 18001
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_622
timestamp 18001
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_623
timestamp 18001
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_624
timestamp 18001
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_625
timestamp 18001
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_626
timestamp 18001
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_627
timestamp 18001
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_628
timestamp 18001
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_629
timestamp 18001
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_630
timestamp 18001
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_631
timestamp 18001
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_632
timestamp 18001
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_633
timestamp 18001
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_634
timestamp 18001
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_635
timestamp 18001
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_636
timestamp 18001
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_637
timestamp 18001
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_638
timestamp 18001
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_639
timestamp 18001
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_640
timestamp 18001
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_641
timestamp 18001
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_642
timestamp 18001
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_643
timestamp 18001
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_644
timestamp 18001
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_645
timestamp 18001
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_646
timestamp 18001
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_647
timestamp 18001
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_648
timestamp 18001
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_649
timestamp 18001
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_650
timestamp 18001
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_651
timestamp 18001
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_652
timestamp 18001
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_653
timestamp 18001
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_654
timestamp 18001
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_655
timestamp 18001
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_656
timestamp 18001
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_657
timestamp 18001
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_658
timestamp 18001
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_659
timestamp 18001
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_660
timestamp 18001
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_661
timestamp 18001
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_662
timestamp 18001
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_663
timestamp 18001
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_664
timestamp 18001
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_665
timestamp 18001
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_666
timestamp 18001
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_667
timestamp 18001
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_668
timestamp 18001
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_669
timestamp 18001
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_670
timestamp 18001
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_671
timestamp 18001
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_672
timestamp 18001
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_673
timestamp 18001
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_674
timestamp 18001
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_675
timestamp 18001
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_676
timestamp 18001
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_677
timestamp 18001
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_678
timestamp 18001
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_679
timestamp 18001
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_680
timestamp 18001
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_681
timestamp 18001
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_682
timestamp 18001
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_683
timestamp 18001
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_684
timestamp 18001
transform 1 0 3680 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_685
timestamp 18001
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_686
timestamp 18001
transform 1 0 8832 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_687
timestamp 18001
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_688
timestamp 18001
transform 1 0 13984 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_689
timestamp 18001
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_690
timestamp 18001
transform 1 0 19136 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_691
timestamp 18001
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_692
timestamp 18001
transform 1 0 24288 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_693
timestamp 18001
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_694
timestamp 18001
transform 1 0 29440 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_695
timestamp 18001
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_696
timestamp 18001
transform 1 0 34592 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_697
timestamp 18001
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_698
timestamp 18001
transform 1 0 39744 0 -1 41344
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 41392 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 41392 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 41392 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 34928 2128 35248 41392 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 38768 800 38888 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 cs
port 3 nsew signal input
flabel metal3 s 40957 23808 41757 23928 0 FreeSans 480 0 0 0 dataBusIn[0]
port 4 nsew signal input
flabel metal2 s 30930 43101 30986 43901 0 FreeSans 224 90 0 0 dataBusIn[1]
port 5 nsew signal input
flabel metal3 s 40957 24488 41757 24608 0 FreeSans 480 0 0 0 dataBusIn[2]
port 6 nsew signal input
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 dataBusIn[3]
port 7 nsew signal input
flabel metal3 s 40957 26528 41757 26648 0 FreeSans 480 0 0 0 dataBusIn[4]
port 8 nsew signal input
flabel metal3 s 40957 17688 41757 17808 0 FreeSans 480 0 0 0 dataBusIn[5]
port 9 nsew signal input
flabel metal3 s 40957 27208 41757 27328 0 FreeSans 480 0 0 0 dataBusIn[6]
port 10 nsew signal input
flabel metal3 s 40957 25848 41757 25968 0 FreeSans 480 0 0 0 dataBusIn[7]
port 11 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 dataBusOut[0]
port 12 nsew signal output
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 dataBusOut[1]
port 13 nsew signal output
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 dataBusOut[2]
port 14 nsew signal output
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 dataBusOut[3]
port 15 nsew signal output
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 dataBusOut[4]
port 16 nsew signal output
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 dataBusOut[5]
port 17 nsew signal output
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 dataBusOut[6]
port 18 nsew signal output
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 dataBusOut[7]
port 19 nsew signal output
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 dataBusSelect
port 20 nsew signal output
flabel metal3 s 0 33328 800 33448 0 FreeSans 480 0 0 0 gpio[0]
port 21 nsew signal bidirectional
flabel metal2 s 23846 43101 23902 43901 0 FreeSans 224 90 0 0 gpio[10]
port 22 nsew signal bidirectional
flabel metal2 s 26422 43101 26478 43901 0 FreeSans 224 90 0 0 gpio[11]
port 23 nsew signal bidirectional
flabel metal2 s 24490 43101 24546 43901 0 FreeSans 224 90 0 0 gpio[12]
port 24 nsew signal bidirectional
flabel metal2 s 25134 43101 25190 43901 0 FreeSans 224 90 0 0 gpio[13]
port 25 nsew signal bidirectional
flabel metal2 s 28354 43101 28410 43901 0 FreeSans 224 90 0 0 gpio[14]
port 26 nsew signal bidirectional
flabel metal2 s 25778 43101 25834 43901 0 FreeSans 224 90 0 0 gpio[15]
port 27 nsew signal bidirectional
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 gpio[16]
port 28 nsew signal bidirectional
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 gpio[17]
port 29 nsew signal bidirectional
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 gpio[18]
port 30 nsew signal bidirectional
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 gpio[19]
port 31 nsew signal bidirectional
flabel metal3 s 0 31288 800 31408 0 FreeSans 480 0 0 0 gpio[1]
port 32 nsew signal bidirectional
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 gpio[20]
port 33 nsew signal bidirectional
flabel metal3 s 40957 16328 41757 16448 0 FreeSans 480 0 0 0 gpio[21]
port 34 nsew signal bidirectional
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 gpio[22]
port 35 nsew signal bidirectional
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 gpio[23]
port 36 nsew signal bidirectional
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 gpio[24]
port 37 nsew signal bidirectional
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 gpio[25]
port 38 nsew signal bidirectional
flabel metal3 s 0 30608 800 30728 0 FreeSans 480 0 0 0 gpio[2]
port 39 nsew signal bidirectional
flabel metal3 s 0 32648 800 32768 0 FreeSans 480 0 0 0 gpio[3]
port 40 nsew signal bidirectional
flabel metal3 s 0 34008 800 34128 0 FreeSans 480 0 0 0 gpio[4]
port 41 nsew signal bidirectional
flabel metal2 s 7102 43101 7158 43901 0 FreeSans 224 90 0 0 gpio[5]
port 42 nsew signal bidirectional
flabel metal3 s 0 34688 800 34808 0 FreeSans 480 0 0 0 gpio[6]
port 43 nsew signal bidirectional
flabel metal3 s 0 36048 800 36168 0 FreeSans 480 0 0 0 gpio[7]
port 44 nsew signal bidirectional
flabel metal2 s 27710 43101 27766 43901 0 FreeSans 224 90 0 0 gpio[8]
port 45 nsew signal bidirectional
flabel metal2 s 27066 43101 27122 43901 0 FreeSans 224 90 0 0 gpio[9]
port 46 nsew signal bidirectional
flabel metal3 s 40957 3408 41757 3528 0 FreeSans 480 0 0 0 nrst
port 47 nsew signal input
rlabel metal1 20838 41344 20838 41344 0 VGND
rlabel metal1 20838 40800 20838 40800 0 VPWR
rlabel metal2 32246 32436 32246 32436 0 _0000_
rlabel metal2 36110 32164 36110 32164 0 _0001_
rlabel metal1 29946 33626 29946 33626 0 _0002_
rlabel metal1 35512 32538 35512 32538 0 _0003_
rlabel metal2 38870 31518 38870 31518 0 _0004_
rlabel metal1 32430 29546 32430 29546 0 _0005_
rlabel metal1 28520 33082 28520 33082 0 _0006_
rlabel metal1 37959 31994 37959 31994 0 _0007_
rlabel metal1 30038 30158 30038 30158 0 _0008_
rlabel metal2 38502 29461 38502 29461 0 _0009_
rlabel via1 38502 30141 38502 30141 0 _0010_
rlabel metal2 32706 33762 32706 33762 0 _0011_
rlabel metal1 30728 31994 30728 31994 0 _0012_
rlabel metal2 29210 28186 29210 28186 0 _0013_
rlabel metal1 25024 5270 25024 5270 0 _0014_
rlabel metal2 27278 5916 27278 5916 0 _0015_
rlabel metal1 29394 5780 29394 5780 0 _0016_
rlabel metal1 30958 6392 30958 6392 0 _0017_
rlabel metal1 25116 4522 25116 4522 0 _0018_
rlabel metal1 28290 5134 28290 5134 0 _0019_
rlabel metal1 38640 7446 38640 7446 0 _0020_
rlabel metal2 39422 10200 39422 10200 0 _0021_
rlabel metal1 37634 6970 37634 6970 0 _0022_
rlabel metal1 38686 8534 38686 8534 0 _0023_
rlabel metal1 38364 23290 38364 23290 0 _0024_
rlabel metal1 37076 14042 37076 14042 0 _0025_
rlabel metal2 20838 30940 20838 30940 0 _0026_
rlabel metal1 19688 31450 19688 31450 0 _0027_
rlabel metal1 28612 4114 28612 4114 0 _0028_
rlabel metal2 18354 4250 18354 4250 0 _0029_
rlabel metal1 17020 5270 17020 5270 0 _0030_
rlabel metal2 20470 6052 20470 6052 0 _0031_
rlabel metal1 19228 5814 19228 5814 0 _0032_
rlabel metal1 22034 4012 22034 4012 0 _0033_
rlabel metal1 16652 2890 16652 2890 0 _0034_
rlabel metal2 14122 3230 14122 3230 0 _0035_
rlabel metal1 12236 4794 12236 4794 0 _0036_
rlabel metal2 10718 5848 10718 5848 0 _0037_
rlabel metal2 12558 3230 12558 3230 0 _0038_
rlabel metal1 11868 2346 11868 2346 0 _0039_
rlabel metal1 11040 3434 11040 3434 0 _0040_
rlabel metal2 14306 4964 14306 4964 0 _0041_
rlabel metal2 13294 38046 13294 38046 0 _0042_
rlabel metal2 13754 35802 13754 35802 0 _0043_
rlabel metal2 15318 37468 15318 37468 0 _0044_
rlabel metal1 19182 38522 19182 38522 0 _0045_
rlabel metal1 19918 37774 19918 37774 0 _0046_
rlabel metal1 19872 35802 19872 35802 0 _0047_
rlabel metal1 19734 34646 19734 34646 0 _0048_
rlabel metal1 18170 33082 18170 33082 0 _0049_
rlabel metal1 12558 23290 12558 23290 0 _0050_
rlabel metal2 7590 24990 7590 24990 0 _0051_
rlabel metal1 4370 23562 4370 23562 0 _0052_
rlabel metal1 2254 24922 2254 24922 0 _0053_
rlabel metal1 4278 25466 4278 25466 0 _0054_
rlabel metal2 1886 26078 1886 26078 0 _0055_
rlabel metal1 2116 23834 2116 23834 0 _0056_
rlabel metal1 10304 21658 10304 21658 0 _0057_
rlabel metal1 11684 20570 11684 20570 0 _0058_
rlabel metal2 7682 21284 7682 21284 0 _0059_
rlabel metal1 3680 21658 3680 21658 0 _0060_
rlabel metal1 3818 21420 3818 21420 0 _0061_
rlabel metal1 4140 20366 4140 20366 0 _0062_
rlabel metal1 2438 20298 2438 20298 0 _0063_
rlabel metal1 2017 22202 2017 22202 0 _0064_
rlabel metal2 9338 20196 9338 20196 0 _0065_
rlabel metal1 22540 5338 22540 5338 0 _0066_
rlabel metal2 25070 36958 25070 36958 0 _0067_
rlabel metal1 27968 38386 27968 38386 0 _0068_
rlabel metal1 22862 37434 22862 37434 0 _0069_
rlabel metal2 24978 38114 24978 38114 0 _0070_
rlabel metal2 23230 38760 23230 38760 0 _0071_
rlabel metal1 23322 35768 23322 35768 0 _0072_
rlabel metal1 25392 35802 25392 35802 0 _0073_
rlabel metal1 24150 34170 24150 34170 0 _0074_
rlabel metal2 14766 34204 14766 34204 0 _0075_
rlabel metal1 12190 34510 12190 34510 0 _0076_
rlabel metal1 7452 32946 7452 32946 0 _0077_
rlabel metal1 4692 32946 4692 32946 0 _0078_
rlabel metal1 6210 34986 6210 34986 0 _0079_
rlabel metal1 6578 37434 6578 37434 0 _0080_
rlabel metal1 8694 38522 8694 38522 0 _0081_
rlabel metal2 10626 36312 10626 36312 0 _0082_
rlabel metal2 12834 18020 12834 18020 0 _0083_
rlabel metal1 7360 28730 7360 28730 0 _0084_
rlabel metal1 6118 28186 6118 28186 0 _0085_
rlabel metal1 3588 27982 3588 27982 0 _0086_
rlabel metal1 5237 28934 5237 28934 0 _0087_
rlabel metal1 4048 27098 4048 27098 0 _0088_
rlabel metal2 4094 29852 4094 29852 0 _0089_
rlabel metal2 8418 27370 8418 27370 0 _0090_
rlabel metal2 3634 32878 3634 32878 0 _0091_
rlabel metal1 4600 30906 4600 30906 0 _0092_
rlabel metal2 3358 30464 3358 30464 0 _0093_
rlabel metal2 2898 33150 2898 33150 0 _0094_
rlabel metal1 3588 34170 3588 34170 0 _0095_
rlabel metal2 4462 38046 4462 38046 0 _0096_
rlabel metal2 3174 35292 3174 35292 0 _0097_
rlabel metal2 4278 35870 4278 35870 0 _0098_
rlabel metal2 15226 11934 15226 11934 0 _0099_
rlabel metal1 3312 12750 3312 12750 0 _0100_
rlabel metal1 6164 15674 6164 15674 0 _0101_
rlabel metal2 3818 11934 3818 11934 0 _0102_
rlabel metal1 4048 16014 4048 16014 0 _0103_
rlabel metal1 5474 8058 5474 8058 0 _0104_
rlabel metal1 5329 10234 5329 10234 0 _0105_
rlabel metal2 9522 7582 9522 7582 0 _0106_
rlabel metal1 11454 18394 11454 18394 0 _0107_
rlabel metal2 7682 19108 7682 19108 0 _0108_
rlabel metal2 4094 18462 4094 18462 0 _0109_
rlabel metal1 3542 19244 3542 19244 0 _0110_
rlabel metal1 5934 18394 5934 18394 0 _0111_
rlabel metal2 2806 17374 2806 17374 0 _0112_
rlabel metal1 2300 18394 2300 18394 0 _0113_
rlabel metal2 9522 19108 9522 19108 0 _0114_
rlabel metal1 17802 31858 17802 31858 0 _0115_
rlabel metal2 30222 33796 30222 33796 0 _0116_
rlabel metal1 15870 6222 15870 6222 0 _0117_
rlabel metal1 8234 11118 8234 11118 0 _0118_
rlabel metal1 7774 11118 7774 11118 0 _0119_
rlabel metal1 8464 11050 8464 11050 0 _0120_
rlabel metal1 6670 19958 6670 19958 0 _0121_
rlabel metal1 6440 22134 6440 22134 0 _0122_
rlabel metal1 6486 21114 6486 21114 0 _0123_
rlabel metal2 6670 21590 6670 21590 0 _0124_
rlabel metal1 12190 31348 12190 31348 0 _0125_
rlabel metal1 10350 30736 10350 30736 0 _0126_
rlabel metal1 13386 26520 13386 26520 0 _0127_
rlabel metal2 19458 8211 19458 8211 0 _0128_
rlabel metal1 18446 23290 18446 23290 0 _0129_
rlabel metal1 12098 26316 12098 26316 0 _0130_
rlabel metal2 12098 24854 12098 24854 0 _0131_
rlabel metal1 9890 30770 9890 30770 0 _0132_
rlabel metal1 7590 17204 7590 17204 0 _0133_
rlabel metal1 7452 16490 7452 16490 0 _0134_
rlabel metal1 11086 15980 11086 15980 0 _0135_
rlabel metal2 12926 5168 12926 5168 0 _0136_
rlabel metal1 7682 16014 7682 16014 0 _0137_
rlabel metal1 7084 25874 7084 25874 0 _0138_
rlabel metal1 7452 26010 7452 26010 0 _0139_
rlabel metal1 7360 17646 7360 17646 0 _0140_
rlabel metal2 7314 17136 7314 17136 0 _0141_
rlabel via1 7306 16422 7306 16422 0 _0142_
rlabel metal2 6854 16048 6854 16048 0 _0143_
rlabel metal2 7038 16082 7038 16082 0 _0144_
rlabel metal2 6026 14144 6026 14144 0 _0145_
rlabel metal1 6762 14994 6762 14994 0 _0146_
rlabel metal2 6762 20468 6762 20468 0 _0147_
rlabel metal1 5980 20570 5980 20570 0 _0148_
rlabel metal1 6808 21046 6808 21046 0 _0149_
rlabel metal1 10626 22406 10626 22406 0 _0150_
rlabel metal2 12374 29818 12374 29818 0 _0151_
rlabel metal1 9752 28526 9752 28526 0 _0152_
rlabel metal2 14766 26622 14766 26622 0 _0153_
rlabel metal1 10166 26384 10166 26384 0 _0154_
rlabel metal1 10212 26486 10212 26486 0 _0155_
rlabel metal1 10120 28390 10120 28390 0 _0156_
rlabel metal1 8740 14926 8740 14926 0 _0157_
rlabel metal1 14398 7820 14398 7820 0 _0158_
rlabel metal1 12006 6698 12006 6698 0 _0159_
rlabel metal1 9614 16490 9614 16490 0 _0160_
rlabel metal2 6026 26554 6026 26554 0 _0161_
rlabel metal1 6762 26554 6762 26554 0 _0162_
rlabel metal1 2645 33490 2645 33490 0 _0163_
rlabel metal1 9430 16660 9430 16660 0 _0164_
rlabel metal1 8832 15130 8832 15130 0 _0165_
rlabel metal1 7406 13362 7406 13362 0 _0166_
rlabel metal2 16146 27098 16146 27098 0 _0167_
rlabel metal2 16790 26112 16790 26112 0 _0168_
rlabel metal2 10350 24480 10350 24480 0 _0169_
rlabel metal2 10810 27506 10810 27506 0 _0170_
rlabel metal1 6164 19278 6164 19278 0 _0171_
rlabel metal2 6394 23290 6394 23290 0 _0172_
rlabel metal1 6486 22746 6486 22746 0 _0173_
rlabel metal1 10304 29614 10304 29614 0 _0174_
rlabel metal2 13846 29240 13846 29240 0 _0175_
rlabel metal2 10442 28730 10442 28730 0 _0176_
rlabel metal1 4646 19244 4646 19244 0 _0177_
rlabel metal2 10074 16490 10074 16490 0 _0178_
rlabel metal1 12788 16082 12788 16082 0 _0179_
rlabel metal1 11960 15402 11960 15402 0 _0180_
rlabel metal2 11822 15674 11822 15674 0 _0181_
rlabel metal1 10948 15538 10948 15538 0 _0182_
rlabel metal1 11362 25160 11362 25160 0 _0183_
rlabel metal2 7866 24004 7866 24004 0 _0184_
rlabel metal1 9016 18734 9016 18734 0 _0185_
rlabel metal1 10074 15674 10074 15674 0 _0186_
rlabel metal1 10488 14382 10488 14382 0 _0187_
rlabel metal1 14306 25874 14306 25874 0 _0188_
rlabel metal1 14398 25772 14398 25772 0 _0189_
rlabel metal1 13570 25840 13570 25840 0 _0190_
rlabel metal1 14030 25670 14030 25670 0 _0191_
rlabel metal1 14030 31382 14030 31382 0 _0192_
rlabel metal1 8418 22678 8418 22678 0 _0193_
rlabel metal1 8648 22610 8648 22610 0 _0194_
rlabel metal1 8648 22202 8648 22202 0 _0195_
rlabel metal2 14306 22848 14306 22848 0 _0196_
rlabel metal1 14996 31858 14996 31858 0 _0197_
rlabel metal1 13524 31790 13524 31790 0 _0198_
rlabel metal2 12650 18445 12650 18445 0 _0199_
rlabel metal2 12466 14416 12466 14416 0 _0200_
rlabel metal1 13800 16626 13800 16626 0 _0201_
rlabel metal1 13708 6834 13708 6834 0 _0202_
rlabel metal1 13202 16456 13202 16456 0 _0203_
rlabel metal1 9154 23290 9154 23290 0 _0204_
rlabel metal2 9798 24956 9798 24956 0 _0205_
rlabel metal1 8872 24174 8872 24174 0 _0206_
rlabel metal2 7406 27404 7406 27404 0 _0207_
rlabel metal2 12512 16422 12512 16422 0 _0208_
rlabel metal1 12190 13906 12190 13906 0 _0209_
rlabel metal1 11776 12818 11776 12818 0 _0210_
rlabel metal1 12926 21930 12926 21930 0 _0211_
rlabel metal2 13386 20944 13386 20944 0 _0212_
rlabel metal1 12972 21386 12972 21386 0 _0213_
rlabel metal1 12742 30124 12742 30124 0 _0214_
rlabel metal1 13156 29546 13156 29546 0 _0215_
rlabel metal2 17066 29580 17066 29580 0 _0216_
rlabel metal1 17158 29172 17158 29172 0 _0217_
rlabel metal2 14398 29444 14398 29444 0 _0218_
rlabel metal1 13984 29750 13984 29750 0 _0219_
rlabel metal1 15042 26860 15042 26860 0 _0220_
rlabel metal2 14950 27132 14950 27132 0 _0221_
rlabel metal2 14858 26724 14858 26724 0 _0222_
rlabel metal1 14260 29614 14260 29614 0 _0223_
rlabel metal1 13662 29648 13662 29648 0 _0224_
rlabel metal1 13064 17578 13064 17578 0 _0225_
rlabel metal1 14030 16422 14030 16422 0 _0226_
rlabel metal1 14306 16558 14306 16558 0 _0227_
rlabel metal1 14858 6630 14858 6630 0 _0228_
rlabel metal2 17066 3536 17066 3536 0 _0229_
rlabel metal1 13478 15912 13478 15912 0 _0230_
rlabel metal1 13984 16014 13984 16014 0 _0231_
rlabel metal1 14628 24378 14628 24378 0 _0232_
rlabel metal2 15226 24208 15226 24208 0 _0233_
rlabel metal2 16606 23426 16606 23426 0 _0234_
rlabel metal1 14352 17238 14352 17238 0 _0235_
rlabel metal1 13547 33422 13547 33422 0 _0236_
rlabel metal2 13662 16524 13662 16524 0 _0237_
rlabel metal1 13432 14994 13432 14994 0 _0238_
rlabel metal1 13570 13838 13570 13838 0 _0239_
rlabel metal2 12880 13906 12880 13906 0 _0240_
rlabel metal1 13064 12410 13064 12410 0 _0241_
rlabel metal1 21252 21862 21252 21862 0 _0242_
rlabel metal1 20608 21658 20608 21658 0 _0243_
rlabel metal1 20884 21998 20884 21998 0 _0244_
rlabel metal1 21482 12818 21482 12818 0 _0245_
rlabel metal1 21528 12614 21528 12614 0 _0246_
rlabel metal2 21022 17442 21022 17442 0 _0247_
rlabel via2 27002 31195 27002 31195 0 _0248_
rlabel metal1 21528 22066 21528 22066 0 _0249_
rlabel metal1 20654 21930 20654 21930 0 _0250_
rlabel metal1 19872 13906 19872 13906 0 _0251_
rlabel metal1 12972 13906 12972 13906 0 _0252_
rlabel metal2 12466 13430 12466 13430 0 _0253_
rlabel metal2 11546 13056 11546 13056 0 _0254_
rlabel metal1 9982 13260 9982 13260 0 _0255_
rlabel metal2 10074 14858 10074 14858 0 _0256_
rlabel metal1 10074 13906 10074 13906 0 _0257_
rlabel metal1 7130 13328 7130 13328 0 _0258_
rlabel via1 8234 13243 8234 13243 0 _0259_
rlabel metal2 7774 13056 7774 13056 0 _0260_
rlabel metal2 5934 13940 5934 13940 0 _0261_
rlabel metal2 6578 14892 6578 14892 0 _0262_
rlabel metal1 6762 14246 6762 14246 0 _0263_
rlabel metal1 7682 10438 7682 10438 0 _0264_
rlabel metal2 10258 10234 10258 10234 0 _0265_
rlabel metal2 11086 9724 11086 9724 0 _0266_
rlabel metal1 12006 9520 12006 9520 0 _0267_
rlabel metal1 14812 9690 14812 9690 0 _0268_
rlabel metal2 14490 10166 14490 10166 0 _0269_
rlabel metal1 14490 10200 14490 10200 0 _0270_
rlabel metal1 7222 12614 7222 12614 0 _0271_
rlabel metal1 14214 11560 14214 11560 0 _0272_
rlabel metal1 12926 14246 12926 14246 0 _0273_
rlabel metal1 11684 14790 11684 14790 0 _0274_
rlabel metal2 10902 8908 10902 8908 0 _0275_
rlabel metal1 9246 13396 9246 13396 0 _0276_
rlabel metal1 8142 12682 8142 12682 0 _0277_
rlabel metal1 5980 13158 5980 13158 0 _0278_
rlabel metal1 6302 12750 6302 12750 0 _0279_
rlabel metal2 4784 13294 4784 13294 0 _0280_
rlabel metal2 7498 11356 7498 11356 0 _0281_
rlabel metal2 4646 14722 4646 14722 0 _0282_
rlabel metal2 7038 9996 7038 9996 0 _0283_
rlabel metal1 11316 7990 11316 7990 0 _0284_
rlabel metal2 9062 8908 9062 8908 0 _0285_
rlabel metal1 8142 8874 8142 8874 0 _0286_
rlabel metal1 7452 9554 7452 9554 0 _0287_
rlabel metal1 7038 8942 7038 8942 0 _0288_
rlabel metal1 8280 7922 8280 7922 0 _0289_
rlabel metal1 11592 8058 11592 8058 0 _0290_
rlabel metal1 9798 7956 9798 7956 0 _0291_
rlabel metal1 10626 8432 10626 8432 0 _0292_
rlabel metal1 10396 8466 10396 8466 0 _0293_
rlabel metal1 10580 8330 10580 8330 0 _0294_
rlabel metal3 16813 20740 16813 20740 0 _0295_
rlabel metal2 17986 7956 17986 7956 0 _0296_
rlabel metal2 17710 7820 17710 7820 0 _0297_
rlabel metal2 18814 8262 18814 8262 0 _0298_
rlabel metal1 17572 7514 17572 7514 0 _0299_
rlabel metal2 15870 8058 15870 8058 0 _0300_
rlabel metal1 16376 7514 16376 7514 0 _0301_
rlabel metal1 23414 14926 23414 14926 0 _0302_
rlabel metal2 20746 13124 20746 13124 0 _0303_
rlabel metal2 15318 7548 15318 7548 0 _0304_
rlabel metal1 14766 7412 14766 7412 0 _0305_
rlabel metal1 14168 6766 14168 6766 0 _0306_
rlabel metal1 14214 6664 14214 6664 0 _0307_
rlabel metal1 13478 6868 13478 6868 0 _0308_
rlabel metal1 15732 6902 15732 6902 0 _0309_
rlabel metal2 18446 7718 18446 7718 0 _0310_
rlabel metal1 20332 5678 20332 5678 0 _0311_
rlabel metal1 14904 8058 14904 8058 0 _0312_
rlabel via2 15686 8483 15686 8483 0 _0313_
rlabel metal2 15318 8262 15318 8262 0 _0314_
rlabel metal1 12466 9452 12466 9452 0 _0315_
rlabel metal1 13386 9350 13386 9350 0 _0316_
rlabel metal1 15042 9554 15042 9554 0 _0317_
rlabel metal1 16928 9350 16928 9350 0 _0318_
rlabel metal1 16560 9554 16560 9554 0 _0319_
rlabel metal1 18538 5066 18538 5066 0 _0320_
rlabel metal1 15226 9588 15226 9588 0 _0321_
rlabel metal1 19964 30906 19964 30906 0 _0322_
rlabel metal1 20516 32198 20516 32198 0 _0323_
rlabel metal1 21712 5678 21712 5678 0 _0324_
rlabel metal2 18722 4930 18722 4930 0 _0325_
rlabel metal1 20470 5712 20470 5712 0 _0326_
rlabel metal1 19642 3978 19642 3978 0 _0327_
rlabel metal2 22402 4522 22402 4522 0 _0328_
rlabel metal1 18308 19210 18308 19210 0 _0329_
rlabel metal1 19228 20570 19228 20570 0 _0330_
rlabel metal1 19044 20842 19044 20842 0 _0331_
rlabel metal1 25668 28186 25668 28186 0 _0332_
rlabel metal1 24886 28560 24886 28560 0 _0333_
rlabel metal1 25254 26554 25254 26554 0 _0334_
rlabel metal2 19918 34170 19918 34170 0 _0335_
rlabel metal1 25438 24922 25438 24922 0 _0336_
rlabel metal2 25898 24820 25898 24820 0 _0337_
rlabel metal2 24518 24990 24518 24990 0 _0338_
rlabel metal1 27186 21896 27186 21896 0 _0339_
rlabel metal1 26312 22066 26312 22066 0 _0340_
rlabel metal1 26772 22678 26772 22678 0 _0341_
rlabel metal1 25668 20502 25668 20502 0 _0342_
rlabel metal1 25530 21896 25530 21896 0 _0343_
rlabel metal2 26266 23341 26266 23341 0 _0344_
rlabel metal1 26496 20434 26496 20434 0 _0345_
rlabel metal2 25714 23664 25714 23664 0 _0346_
rlabel metal2 24426 25092 24426 25092 0 _0347_
rlabel via2 24886 25483 24886 25483 0 _0348_
rlabel metal2 23138 28985 23138 28985 0 _0349_
rlabel metal1 23184 30906 23184 30906 0 _0350_
rlabel metal2 22862 31280 22862 31280 0 _0351_
rlabel metal1 16422 33048 16422 33048 0 _0352_
rlabel metal1 22494 26418 22494 26418 0 _0353_
rlabel metal2 16514 32929 16514 32929 0 _0354_
rlabel metal2 15318 34068 15318 34068 0 _0355_
rlabel metal2 15686 34306 15686 34306 0 _0356_
rlabel metal1 22770 31450 22770 31450 0 _0357_
rlabel metal1 11592 35734 11592 35734 0 _0358_
rlabel metal2 12190 39610 12190 39610 0 _0359_
rlabel metal1 11914 39508 11914 39508 0 _0360_
rlabel metal2 11546 38964 11546 38964 0 _0361_
rlabel metal1 11822 38964 11822 38964 0 _0362_
rlabel metal1 11224 38862 11224 38862 0 _0363_
rlabel metal1 10120 38522 10120 38522 0 _0364_
rlabel metal1 9430 38318 9430 38318 0 _0365_
rlabel metal1 8832 38318 8832 38318 0 _0366_
rlabel metal1 9430 37808 9430 37808 0 _0367_
rlabel metal2 9154 37434 9154 37434 0 _0368_
rlabel metal1 9016 36754 9016 36754 0 _0369_
rlabel metal1 8786 35258 8786 35258 0 _0370_
rlabel metal2 9154 35258 9154 35258 0 _0371_
rlabel metal1 9016 35122 9016 35122 0 _0372_
rlabel metal2 9154 34170 9154 34170 0 _0373_
rlabel metal1 9430 34000 9430 34000 0 _0374_
rlabel metal1 10074 33626 10074 33626 0 _0375_
rlabel metal1 10534 33456 10534 33456 0 _0376_
rlabel metal1 10488 33966 10488 33966 0 _0377_
rlabel metal2 10994 34306 10994 34306 0 _0378_
rlabel metal1 12558 34170 12558 34170 0 _0379_
rlabel metal1 10718 34170 10718 34170 0 _0380_
rlabel metal1 10166 34034 10166 34034 0 _0381_
rlabel metal1 9338 35156 9338 35156 0 _0382_
rlabel metal2 8510 36958 8510 36958 0 _0383_
rlabel via2 9062 38301 9062 38301 0 _0384_
rlabel metal2 9430 38964 9430 38964 0 _0385_
rlabel metal1 11730 39610 11730 39610 0 _0386_
rlabel metal2 13662 39746 13662 39746 0 _0387_
rlabel metal1 12834 39338 12834 39338 0 _0388_
rlabel metal2 13018 38828 13018 38828 0 _0389_
rlabel metal1 7360 33490 7360 33490 0 _0390_
rlabel metal2 7406 34204 7406 34204 0 _0391_
rlabel metal1 8188 36210 8188 36210 0 _0392_
rlabel metal2 14030 36924 14030 36924 0 _0393_
rlabel metal2 14674 30107 14674 30107 0 _0394_
rlabel metal2 12558 32436 12558 32436 0 _0395_
rlabel metal1 12131 30226 12131 30226 0 _0396_
rlabel metal2 13294 30430 13294 30430 0 _0397_
rlabel metal1 13616 30226 13616 30226 0 _0398_
rlabel metal1 15778 35734 15778 35734 0 _0399_
rlabel metal1 5566 32402 5566 32402 0 _0400_
rlabel metal1 6302 33490 6302 33490 0 _0401_
rlabel metal1 12834 36176 12834 36176 0 _0402_
rlabel metal1 15686 35734 15686 35734 0 _0403_
rlabel metal2 12282 36890 12282 36890 0 _0404_
rlabel metal1 16330 36788 16330 36788 0 _0405_
rlabel metal1 12604 36890 12604 36890 0 _0406_
rlabel metal2 12650 37876 12650 37876 0 _0407_
rlabel metal2 19458 35734 19458 35734 0 _0408_
rlabel via1 10833 34578 10833 34578 0 _0409_
rlabel metal1 13938 40052 13938 40052 0 _0410_
rlabel metal1 14214 39950 14214 39950 0 _0411_
rlabel metal1 14398 36822 14398 36822 0 _0412_
rlabel metal1 14168 32334 14168 32334 0 _0413_
rlabel metal1 14168 31450 14168 31450 0 _0414_
rlabel metal1 17066 36788 17066 36788 0 _0415_
rlabel metal1 14076 36074 14076 36074 0 _0416_
rlabel metal1 13202 36686 13202 36686 0 _0417_
rlabel metal1 13800 36550 13800 36550 0 _0418_
rlabel metal2 14582 36380 14582 36380 0 _0419_
rlabel metal1 16238 40494 16238 40494 0 _0420_
rlabel metal1 15594 39882 15594 39882 0 _0421_
rlabel metal2 14674 39168 14674 39168 0 _0422_
rlabel metal1 16100 40358 16100 40358 0 _0423_
rlabel metal1 15410 39406 15410 39406 0 _0424_
rlabel metal2 15870 38556 15870 38556 0 _0425_
rlabel metal1 15778 37876 15778 37876 0 _0426_
rlabel metal1 15594 36754 15594 36754 0 _0427_
rlabel metal2 15686 36992 15686 36992 0 _0428_
rlabel metal2 11362 29444 11362 29444 0 _0429_
rlabel metal1 19550 37128 19550 37128 0 _0430_
rlabel metal1 15272 36346 15272 36346 0 _0431_
rlabel metal1 15180 37434 15180 37434 0 _0432_
rlabel metal2 17158 39712 17158 39712 0 _0433_
rlabel metal1 16698 40630 16698 40630 0 _0434_
rlabel metal2 17986 38794 17986 38794 0 _0435_
rlabel metal1 17894 36652 17894 36652 0 _0436_
rlabel metal2 16146 35428 16146 35428 0 _0437_
rlabel metal1 17664 37434 17664 37434 0 _0438_
rlabel metal1 11500 28730 11500 28730 0 _0439_
rlabel metal1 14904 35122 14904 35122 0 _0440_
rlabel metal1 19826 37638 19826 37638 0 _0441_
rlabel metal2 17342 37604 17342 37604 0 _0442_
rlabel metal1 17940 37978 17940 37978 0 _0443_
rlabel metal1 21574 38284 21574 38284 0 _0444_
rlabel metal1 21620 37434 21620 37434 0 _0445_
rlabel metal2 22126 38080 22126 38080 0 _0446_
rlabel metal1 20838 37264 20838 37264 0 _0447_
rlabel metal2 16974 39372 16974 39372 0 _0448_
rlabel metal2 16698 39134 16698 39134 0 _0449_
rlabel metal1 19918 37298 19918 37298 0 _0450_
rlabel metal1 19872 37434 19872 37434 0 _0451_
rlabel metal2 18262 37060 18262 37060 0 _0452_
rlabel metal1 19090 37094 19090 37094 0 _0453_
rlabel metal2 10994 32164 10994 32164 0 _0454_
rlabel metal1 16054 34986 16054 34986 0 _0455_
rlabel metal1 23322 38250 23322 38250 0 _0456_
rlabel metal1 19228 36686 19228 36686 0 _0457_
rlabel metal2 18998 37366 18998 37366 0 _0458_
rlabel metal2 21942 36890 21942 36890 0 _0459_
rlabel metal2 22310 35700 22310 35700 0 _0460_
rlabel viali 21573 35666 21573 35666 0 _0461_
rlabel metal1 22218 36210 22218 36210 0 _0462_
rlabel metal1 21574 36244 21574 36244 0 _0463_
rlabel metal1 12649 31790 12649 31790 0 _0464_
rlabel metal2 17066 33796 17066 33796 0 _0465_
rlabel metal2 17986 35802 17986 35802 0 _0466_
rlabel metal1 17158 35632 17158 35632 0 _0467_
rlabel metal1 17986 35666 17986 35666 0 _0468_
rlabel metal1 18308 35598 18308 35598 0 _0469_
rlabel metal1 19090 35598 19090 35598 0 _0470_
rlabel via1 21850 34493 21850 34493 0 _0471_
rlabel via2 21482 35020 21482 35020 0 _0472_
rlabel metal1 21436 34034 21436 34034 0 _0473_
rlabel metal1 21620 34102 21620 34102 0 _0474_
rlabel metal1 17802 35190 17802 35190 0 _0475_
rlabel metal1 18446 34714 18446 34714 0 _0476_
rlabel metal2 11086 32368 11086 32368 0 _0477_
rlabel metal1 16698 34578 16698 34578 0 _0478_
rlabel metal1 18722 34170 18722 34170 0 _0479_
rlabel metal1 18768 34578 18768 34578 0 _0480_
rlabel metal1 21160 33966 21160 33966 0 _0481_
rlabel metal2 20194 33830 20194 33830 0 _0482_
rlabel metal1 17802 32912 17802 32912 0 _0483_
rlabel metal1 17710 34646 17710 34646 0 _0484_
rlabel metal2 17434 34170 17434 34170 0 _0485_
rlabel metal2 12466 29750 12466 29750 0 _0486_
rlabel metal1 18124 34034 18124 34034 0 _0487_
rlabel metal1 17434 34034 17434 34034 0 _0488_
rlabel metal2 17618 33354 17618 33354 0 _0489_
rlabel metal2 22402 17850 22402 17850 0 _0490_
rlabel metal1 20792 17714 20792 17714 0 _0491_
rlabel metal1 29440 20366 29440 20366 0 _0492_
rlabel via2 16330 20451 16330 20451 0 _0493_
rlabel metal1 13202 20434 13202 20434 0 _0494_
rlabel metal2 22402 5406 22402 5406 0 _0495_
rlabel metal1 25885 22610 25885 22610 0 _0496_
rlabel metal1 25254 24718 25254 24718 0 _0497_
rlabel metal1 29072 23834 29072 23834 0 _0498_
rlabel metal2 28014 24412 28014 24412 0 _0499_
rlabel metal1 28842 24072 28842 24072 0 _0500_
rlabel metal1 28704 24310 28704 24310 0 _0501_
rlabel metal1 26312 24650 26312 24650 0 _0502_
rlabel metal2 26542 31110 26542 31110 0 _0503_
rlabel metal1 26128 31450 26128 31450 0 _0504_
rlabel metal1 25392 32334 25392 32334 0 _0505_
rlabel metal1 25116 34034 25116 34034 0 _0506_
rlabel metal1 14260 33626 14260 33626 0 _0507_
rlabel metal1 7866 30634 7866 30634 0 _0508_
rlabel metal1 8602 30634 8602 30634 0 _0509_
rlabel metal2 8602 31076 8602 31076 0 _0510_
rlabel metal2 11040 31892 11040 31892 0 _0511_
rlabel metal1 12144 34170 12144 34170 0 _0512_
rlabel metal2 11362 34748 11362 34748 0 _0513_
rlabel metal1 8004 30906 8004 30906 0 _0514_
rlabel metal2 7406 32266 7406 32266 0 _0515_
rlabel metal2 10258 33932 10258 33932 0 _0516_
rlabel metal1 8050 33524 8050 33524 0 _0517_
rlabel metal1 7728 32538 7728 32538 0 _0518_
rlabel metal2 5842 32538 5842 32538 0 _0519_
rlabel metal1 9476 33354 9476 33354 0 _0520_
rlabel metal1 7866 33626 7866 33626 0 _0521_
rlabel metal1 6486 32538 6486 32538 0 _0522_
rlabel metal1 6026 33626 6026 33626 0 _0523_
rlabel metal1 9108 34714 9108 34714 0 _0524_
rlabel metal1 8004 35190 8004 35190 0 _0525_
rlabel via1 6026 35802 6026 35802 0 _0526_
rlabel metal2 6578 34748 6578 34748 0 _0527_
rlabel metal1 5612 32198 5612 32198 0 _0528_
rlabel metal1 6394 33558 6394 33558 0 _0529_
rlabel metal1 7084 34714 7084 34714 0 _0530_
rlabel metal2 7222 35258 7222 35258 0 _0531_
rlabel metal2 5842 36924 5842 36924 0 _0532_
rlabel metal1 5934 37264 5934 37264 0 _0533_
rlabel metal2 6026 37060 6026 37060 0 _0534_
rlabel metal2 8418 37060 8418 37060 0 _0535_
rlabel metal1 5750 37196 5750 37196 0 _0536_
rlabel metal1 8234 38522 8234 38522 0 _0537_
rlabel metal2 8326 38794 8326 38794 0 _0538_
rlabel metal1 6854 36142 6854 36142 0 _0539_
rlabel metal2 7590 35938 7590 35938 0 _0540_
rlabel metal1 9798 36176 9798 36176 0 _0541_
rlabel metal1 7360 36074 7360 36074 0 _0542_
rlabel metal2 7866 36788 7866 36788 0 _0543_
rlabel metal1 8004 37434 8004 37434 0 _0544_
rlabel metal2 11086 39100 11086 39100 0 _0545_
rlabel metal1 10994 36788 10994 36788 0 _0546_
rlabel metal1 10534 35598 10534 35598 0 _0547_
rlabel metal1 10856 35802 10856 35802 0 _0548_
rlabel metal2 11178 36142 11178 36142 0 _0549_
rlabel metal1 24656 15130 24656 15130 0 _0550_
rlabel metal1 25530 15504 25530 15504 0 _0551_
rlabel metal1 16422 17714 16422 17714 0 _0552_
rlabel metal1 27462 24208 27462 24208 0 _0553_
rlabel metal1 27830 23834 27830 23834 0 _0554_
rlabel metal1 28106 22542 28106 22542 0 _0555_
rlabel metal2 27554 23392 27554 23392 0 _0556_
rlabel metal1 27140 24378 27140 24378 0 _0557_
rlabel metal1 24932 24786 24932 24786 0 _0558_
rlabel metal1 25208 31246 25208 31246 0 _0559_
rlabel metal2 2254 34578 2254 34578 0 _0560_
rlabel metal1 13800 11118 13800 11118 0 _0561_
rlabel metal1 14674 11322 14674 11322 0 _0562_
rlabel metal1 14444 13158 14444 13158 0 _0563_
rlabel metal1 10258 14450 10258 14450 0 _0564_
rlabel metal1 12926 11152 12926 11152 0 _0565_
rlabel metal1 13018 13328 13018 13328 0 _0566_
rlabel metal1 14214 13906 14214 13906 0 _0567_
rlabel metal2 14122 13158 14122 13158 0 _0568_
rlabel metal2 12834 13498 12834 13498 0 _0569_
rlabel metal2 13754 12988 13754 12988 0 _0570_
rlabel metal1 14766 12682 14766 12682 0 _0571_
rlabel metal1 19366 12954 19366 12954 0 _0572_
rlabel metal1 16330 13328 16330 13328 0 _0573_
rlabel metal1 16008 13498 16008 13498 0 _0574_
rlabel metal2 15870 14790 15870 14790 0 _0575_
rlabel metal1 15134 14858 15134 14858 0 _0576_
rlabel metal1 4876 13158 4876 13158 0 _0577_
rlabel metal1 7774 12410 7774 12410 0 _0578_
rlabel metal2 12558 13464 12558 13464 0 _0579_
rlabel metal1 10534 12818 10534 12818 0 _0580_
rlabel metal1 10948 12818 10948 12818 0 _0581_
rlabel metal1 7774 12852 7774 12852 0 _0582_
rlabel metal1 4830 12818 4830 12818 0 _0583_
rlabel metal2 4600 12716 4600 12716 0 _0584_
rlabel metal2 4692 12852 4692 12852 0 _0585_
rlabel metal1 14352 12614 14352 12614 0 _0586_
rlabel metal1 4508 13498 4508 13498 0 _0587_
rlabel metal1 3818 13498 3818 13498 0 _0588_
rlabel metal1 4232 14042 4232 14042 0 _0589_
rlabel metal1 10304 14586 10304 14586 0 _0590_
rlabel metal1 9338 14892 9338 14892 0 _0591_
rlabel metal1 9384 14586 9384 14586 0 _0592_
rlabel metal1 5382 14960 5382 14960 0 _0593_
rlabel metal1 5428 15130 5428 15130 0 _0594_
rlabel metal1 5198 14586 5198 14586 0 _0595_
rlabel metal1 6118 12614 6118 12614 0 _0596_
rlabel metal1 5842 12104 5842 12104 0 _0597_
rlabel metal1 6072 11866 6072 11866 0 _0598_
rlabel metal1 7866 13328 7866 13328 0 _0599_
rlabel metal2 8326 12988 8326 12988 0 _0600_
rlabel metal1 7130 12138 7130 12138 0 _0601_
rlabel metal2 6486 14620 6486 14620 0 _0602_
rlabel metal2 7222 14586 7222 14586 0 _0603_
rlabel metal1 6762 14484 6762 14484 0 _0604_
rlabel metal2 6302 14960 6302 14960 0 _0605_
rlabel metal2 4646 15232 4646 15232 0 _0606_
rlabel metal2 5474 15878 5474 15878 0 _0607_
rlabel metal1 8924 11186 8924 11186 0 _0608_
rlabel metal2 8694 11424 8694 11424 0 _0609_
rlabel metal2 7130 10642 7130 10642 0 _0610_
rlabel metal1 7498 10064 7498 10064 0 _0611_
rlabel metal2 7314 9418 7314 9418 0 _0612_
rlabel metal1 7038 8466 7038 8466 0 _0613_
rlabel metal1 6900 8398 6900 8398 0 _0614_
rlabel metal2 6670 8636 6670 8636 0 _0615_
rlabel metal1 6026 7854 6026 7854 0 _0616_
rlabel metal1 9476 10234 9476 10234 0 _0617_
rlabel metal2 9338 9758 9338 9758 0 _0618_
rlabel metal1 10120 10778 10120 10778 0 _0619_
rlabel metal1 10212 11118 10212 11118 0 _0620_
rlabel metal2 9430 10302 9430 10302 0 _0621_
rlabel metal1 8832 9690 8832 9690 0 _0622_
rlabel metal2 7774 8772 7774 8772 0 _0623_
rlabel metal1 7958 7990 7958 7990 0 _0624_
rlabel metal1 7130 7922 7130 7922 0 _0625_
rlabel metal1 7176 7990 7176 7990 0 _0626_
rlabel metal1 7084 8602 7084 8602 0 _0627_
rlabel metal1 13064 9554 13064 9554 0 _0628_
rlabel metal1 13018 9146 13018 9146 0 _0629_
rlabel metal2 12650 10438 12650 10438 0 _0630_
rlabel metal2 12466 10948 12466 10948 0 _0631_
rlabel metal2 13478 9996 13478 9996 0 _0632_
rlabel metal1 12742 9384 12742 9384 0 _0633_
rlabel metal1 10166 7922 10166 7922 0 _0634_
rlabel metal1 9108 7854 9108 7854 0 _0635_
rlabel metal1 25576 14586 25576 14586 0 _0636_
rlabel metal2 12282 17204 12282 17204 0 _0637_
rlabel metal1 18308 30362 18308 30362 0 _0638_
rlabel metal2 30130 32844 30130 32844 0 _0639_
rlabel metal1 18170 6834 18170 6834 0 _0640_
rlabel via2 24702 13957 24702 13957 0 _0641_
rlabel metal2 28658 8160 28658 8160 0 _0642_
rlabel metal1 28336 26010 28336 26010 0 _0643_
rlabel metal1 25300 31858 25300 31858 0 _0644_
rlabel metal1 15870 7378 15870 7378 0 _0645_
rlabel metal1 17802 10030 17802 10030 0 _0646_
rlabel metal3 19412 15164 19412 15164 0 _0647_
rlabel metal2 32154 27200 32154 27200 0 _0648_
rlabel via1 19918 5678 19918 5678 0 _0649_
rlabel metal1 32108 31858 32108 31858 0 _0650_
rlabel metal1 28750 32368 28750 32368 0 _0651_
rlabel metal1 31924 32538 31924 32538 0 _0652_
rlabel metal1 21850 4148 21850 4148 0 _0653_
rlabel metal2 33810 9282 33810 9282 0 _0654_
rlabel metal1 13248 13906 13248 13906 0 _0655_
rlabel metal1 23920 14042 23920 14042 0 _0656_
rlabel metal1 32844 7922 32844 7922 0 _0657_
rlabel metal1 30314 8262 30314 8262 0 _0658_
rlabel metal2 20700 21998 20700 21998 0 _0659_
rlabel metal2 37674 9350 37674 9350 0 _0660_
rlabel metal1 22854 7514 22854 7514 0 _0661_
rlabel metal1 26726 8262 26726 8262 0 _0662_
rlabel metal2 22954 19125 22954 19125 0 _0663_
rlabel metal1 23046 14416 23046 14416 0 _0664_
rlabel metal1 15502 14348 15502 14348 0 _0665_
rlabel metal2 34270 8755 34270 8755 0 _0666_
rlabel metal1 28566 23664 28566 23664 0 _0667_
rlabel via2 37766 8483 37766 8483 0 _0668_
rlabel metal1 25024 7174 25024 7174 0 _0669_
rlabel metal2 31878 17765 31878 17765 0 _0670_
rlabel metal2 28382 16490 28382 16490 0 _0671_
rlabel metal1 33718 6834 33718 6834 0 _0672_
rlabel metal1 19136 10098 19136 10098 0 _0673_
rlabel metal1 32062 10234 32062 10234 0 _0674_
rlabel metal1 30774 20842 30774 20842 0 _0675_
rlabel metal1 26864 18938 26864 18938 0 _0676_
rlabel metal1 25714 31926 25714 31926 0 _0677_
rlabel metal1 18032 19414 18032 19414 0 _0678_
rlabel metal1 24886 27302 24886 27302 0 _0679_
rlabel metal1 23000 23698 23000 23698 0 _0680_
rlabel metal1 24610 22406 24610 22406 0 _0681_
rlabel metal2 32614 16915 32614 16915 0 _0682_
rlabel metal1 26726 8942 26726 8942 0 _0683_
rlabel metal2 20516 19924 20516 19924 0 _0684_
rlabel metal1 30268 11322 30268 11322 0 _0685_
rlabel metal1 25346 12852 25346 12852 0 _0686_
rlabel metal1 25868 8874 25868 8874 0 _0687_
rlabel metal1 19090 10200 19090 10200 0 _0688_
rlabel metal2 32982 14178 32982 14178 0 _0689_
rlabel metal2 33902 11730 33902 11730 0 _0690_
rlabel metal1 25760 12614 25760 12614 0 _0691_
rlabel metal2 26542 13566 26542 13566 0 _0692_
rlabel metal2 29854 10336 29854 10336 0 _0693_
rlabel metal1 37030 14450 37030 14450 0 _0694_
rlabel via3 34707 13124 34707 13124 0 _0695_
rlabel metal1 12972 12818 12972 12818 0 _0696_
rlabel metal2 25622 13022 25622 13022 0 _0697_
rlabel metal2 18538 18326 18538 18326 0 _0698_
rlabel metal2 23874 15436 23874 15436 0 _0699_
rlabel metal1 33994 20366 33994 20366 0 _0700_
rlabel metal1 31142 21318 31142 21318 0 _0701_
rlabel metal3 37237 21012 37237 21012 0 _0702_
rlabel metal2 18722 8976 18722 8976 0 _0703_
rlabel metal3 26841 28492 26841 28492 0 _0704_
rlabel via1 28298 7718 28298 7718 0 _0705_
rlabel metal1 27554 12750 27554 12750 0 _0706_
rlabel metal2 36478 21318 36478 21318 0 _0707_
rlabel metal1 26266 13804 26266 13804 0 _0708_
rlabel metal1 24196 12682 24196 12682 0 _0709_
rlabel metal1 24150 12886 24150 12886 0 _0710_
rlabel metal1 21896 2346 21896 2346 0 _0711_
rlabel metal4 17756 12036 17756 12036 0 _0712_
rlabel metal1 23368 27098 23368 27098 0 _0713_
rlabel metal1 24702 5338 24702 5338 0 _0714_
rlabel metal1 21942 4080 21942 4080 0 _0715_
rlabel metal2 16652 17204 16652 17204 0 _0716_
rlabel metal2 34362 7871 34362 7871 0 _0717_
rlabel metal1 35236 8466 35236 8466 0 _0718_
rlabel metal2 28750 8772 28750 8772 0 _0719_
rlabel via2 33626 11747 33626 11747 0 _0720_
rlabel metal3 38157 18020 38157 18020 0 _0721_
rlabel metal2 28658 8738 28658 8738 0 _0722_
rlabel metal1 33189 9622 33189 9622 0 _0723_
rlabel metal1 19274 24718 19274 24718 0 _0724_
rlabel metal2 25714 8636 25714 8636 0 _0725_
rlabel metal1 25622 7990 25622 7990 0 _0726_
rlabel metal2 25254 8636 25254 8636 0 _0727_
rlabel metal2 25070 7616 25070 7616 0 _0728_
rlabel metal1 25070 7786 25070 7786 0 _0729_
rlabel metal1 24886 8432 24886 8432 0 _0730_
rlabel metal1 24886 7514 24886 7514 0 _0731_
rlabel metal1 25208 24174 25208 24174 0 _0732_
rlabel via2 24702 8075 24702 8075 0 _0733_
rlabel metal1 26588 24718 26588 24718 0 _0734_
rlabel metal1 16514 20774 16514 20774 0 _0735_
rlabel metal1 27278 26350 27278 26350 0 _0736_
rlabel metal1 26726 17646 26726 17646 0 _0737_
rlabel metal1 29256 21862 29256 21862 0 _0738_
rlabel metal1 34592 19414 34592 19414 0 _0739_
rlabel metal1 26726 18054 26726 18054 0 _0740_
rlabel metal2 24242 17340 24242 17340 0 _0741_
rlabel metal2 18446 15674 18446 15674 0 _0742_
rlabel metal2 26864 15334 26864 15334 0 _0743_
rlabel metal2 29670 22899 29670 22899 0 _0744_
rlabel metal2 20102 8160 20102 8160 0 _0745_
rlabel metal1 20654 9384 20654 9384 0 _0746_
rlabel metal1 22862 14348 22862 14348 0 _0747_
rlabel metal2 22494 15334 22494 15334 0 _0748_
rlabel metal1 22632 16558 22632 16558 0 _0749_
rlabel metal1 20378 18870 20378 18870 0 _0750_
rlabel metal1 35098 16490 35098 16490 0 _0751_
rlabel metal1 25806 16587 25806 16587 0 _0752_
rlabel metal1 23046 9520 23046 9520 0 _0753_
rlabel metal1 23690 17102 23690 17102 0 _0754_
rlabel metal1 31142 13906 31142 13906 0 _0755_
rlabel metal1 32062 13192 32062 13192 0 _0756_
rlabel metal2 20470 7599 20470 7599 0 _0757_
rlabel metal1 27462 21964 27462 21964 0 _0758_
rlabel metal2 25714 16388 25714 16388 0 _0759_
rlabel metal1 25898 20230 25898 20230 0 _0760_
rlabel via1 25438 20298 25438 20298 0 _0761_
rlabel metal1 25254 20366 25254 20366 0 _0762_
rlabel metal2 25990 20570 25990 20570 0 _0763_
rlabel metal1 26450 19822 26450 19822 0 _0764_
rlabel metal3 34316 16456 34316 16456 0 _0765_
rlabel metal2 29854 20332 29854 20332 0 _0766_
rlabel metal2 31970 20910 31970 20910 0 _0767_
rlabel metal1 29118 17646 29118 17646 0 _0768_
rlabel metal2 28842 18224 28842 18224 0 _0769_
rlabel metal1 28336 7990 28336 7990 0 _0770_
rlabel metal2 25070 20162 25070 20162 0 _0771_
rlabel metal2 28842 17476 28842 17476 0 _0772_
rlabel metal1 27416 17714 27416 17714 0 _0773_
rlabel metal1 20470 11594 20470 11594 0 _0774_
rlabel metal1 18860 12206 18860 12206 0 _0775_
rlabel metal2 33626 15470 33626 15470 0 _0776_
rlabel metal1 28888 14450 28888 14450 0 _0777_
rlabel metal1 27646 14348 27646 14348 0 _0778_
rlabel metal2 26450 14824 26450 14824 0 _0779_
rlabel metal2 32430 22236 32430 22236 0 _0780_
rlabel metal1 29854 15538 29854 15538 0 _0781_
rlabel metal1 30498 12954 30498 12954 0 _0782_
rlabel metal2 27554 20247 27554 20247 0 _0783_
rlabel metal2 28934 14926 28934 14926 0 _0784_
rlabel via2 28566 14603 28566 14603 0 _0785_
rlabel metal1 23506 17578 23506 17578 0 _0786_
rlabel via2 21850 10659 21850 10659 0 _0787_
rlabel metal1 24242 17238 24242 17238 0 _0788_
rlabel metal1 25898 14042 25898 14042 0 _0789_
rlabel metal2 30038 16354 30038 16354 0 _0790_
rlabel metal1 33166 13328 33166 13328 0 _0791_
rlabel metal2 30314 14586 30314 14586 0 _0792_
rlabel metal2 24518 11815 24518 11815 0 _0793_
rlabel metal2 18538 11169 18538 11169 0 _0794_
rlabel via1 28290 11322 28290 11322 0 _0795_
rlabel via2 37214 19771 37214 19771 0 _0796_
rlabel metal2 28474 14960 28474 14960 0 _0797_
rlabel metal2 24426 17442 24426 17442 0 _0798_
rlabel metal1 28198 14348 28198 14348 0 _0799_
rlabel metal1 28152 14042 28152 14042 0 _0800_
rlabel metal1 27876 14586 27876 14586 0 _0801_
rlabel metal2 27186 17340 27186 17340 0 _0802_
rlabel metal1 33948 26350 33948 26350 0 _0803_
rlabel metal1 33442 31246 33442 31246 0 _0804_
rlabel metal1 27186 31348 27186 31348 0 _0805_
rlabel metal1 26910 26316 26910 26316 0 _0806_
rlabel metal2 25162 29410 25162 29410 0 _0807_
rlabel metal1 26266 24072 26266 24072 0 _0808_
rlabel metal1 22609 30226 22609 30226 0 _0809_
rlabel via1 28579 29206 28579 29206 0 _0810_
rlabel metal1 28842 29648 28842 29648 0 _0811_
rlabel metal2 21942 27302 21942 27302 0 _0812_
rlabel metal1 27784 29070 27784 29070 0 _0813_
rlabel via2 25346 29597 25346 29597 0 _0814_
rlabel metal2 26266 29818 26266 29818 0 _0815_
rlabel metal1 26450 31688 26450 31688 0 _0816_
rlabel metal3 27117 17748 27117 17748 0 _0817_
rlabel metal1 27232 29002 27232 29002 0 _0818_
rlabel metal1 29624 32334 29624 32334 0 _0819_
rlabel metal1 29624 6698 29624 6698 0 _0820_
rlabel metal1 29854 25330 29854 25330 0 _0821_
rlabel metal2 39146 27166 39146 27166 0 _0822_
rlabel metal1 29946 27098 29946 27098 0 _0823_
rlabel via2 21390 5355 21390 5355 0 _0824_
rlabel metal1 21390 5644 21390 5644 0 _0825_
rlabel metal1 38865 19482 38865 19482 0 _0826_
rlabel metal2 38870 29070 38870 29070 0 _0827_
rlabel metal1 35374 29002 35374 29002 0 _0828_
rlabel metal1 31234 30192 31234 30192 0 _0829_
rlabel metal1 38272 30634 38272 30634 0 _0830_
rlabel metal2 34270 28730 34270 28730 0 _0831_
rlabel metal1 35834 30770 35834 30770 0 _0832_
rlabel metal1 37996 29614 37996 29614 0 _0833_
rlabel metal1 38318 28730 38318 28730 0 _0834_
rlabel metal1 38318 29070 38318 29070 0 _0835_
rlabel metal3 32361 13668 32361 13668 0 _0836_
rlabel metal1 38640 20910 38640 20910 0 _0837_
rlabel via1 36746 29206 36746 29206 0 _0838_
rlabel viali 33625 29138 33625 29138 0 _0839_
rlabel metal1 36064 30906 36064 30906 0 _0840_
rlabel metal1 37214 30906 37214 30906 0 _0841_
rlabel metal1 38226 31110 38226 31110 0 _0842_
rlabel metal1 35988 29546 35988 29546 0 _0843_
rlabel metal1 34040 29614 34040 29614 0 _0844_
rlabel metal1 36248 29818 36248 29818 0 _0845_
rlabel metal1 36708 31314 36708 31314 0 _0846_
rlabel metal1 37444 31450 37444 31450 0 _0847_
rlabel metal1 35374 25194 35374 25194 0 _0848_
rlabel metal1 38180 30906 38180 30906 0 _0849_
rlabel metal1 39238 15470 39238 15470 0 _0850_
rlabel metal1 36984 30022 36984 30022 0 _0851_
rlabel metal1 31418 30634 31418 30634 0 _0852_
rlabel metal2 32338 17068 32338 17068 0 _0853_
rlabel metal1 30866 30294 30866 30294 0 _0854_
rlabel metal1 30958 30226 30958 30226 0 _0855_
rlabel metal3 34960 26180 34960 26180 0 _0856_
rlabel metal1 29716 33490 29716 33490 0 _0857_
rlabel metal1 29624 33082 29624 33082 0 _0858_
rlabel metal1 33580 28934 33580 28934 0 _0859_
rlabel via1 32724 29138 32724 29138 0 _0860_
rlabel metal1 32430 28526 32430 28526 0 _0861_
rlabel metal2 32154 27676 32154 27676 0 _0862_
rlabel metal1 32660 20434 32660 20434 0 _0863_
rlabel metal1 32798 31790 32798 31790 0 _0864_
rlabel metal1 32430 31756 32430 31756 0 _0865_
rlabel metal1 31326 19856 31326 19856 0 _0866_
rlabel metal1 32982 29138 32982 29138 0 _0867_
rlabel metal1 32522 29274 32522 29274 0 _0868_
rlabel metal1 35236 31858 35236 31858 0 _0869_
rlabel metal1 31464 30090 31464 30090 0 _0870_
rlabel metal1 34730 21624 34730 21624 0 _0871_
rlabel metal2 33626 31008 33626 31008 0 _0872_
rlabel metal1 31556 31790 31556 31790 0 _0873_
rlabel metal1 36340 21590 36340 21590 0 _0874_
rlabel metal1 36892 14382 36892 14382 0 _0875_
rlabel metal1 35420 26962 35420 26962 0 _0876_
rlabel metal2 31878 25738 31878 25738 0 _0877_
rlabel metal1 32292 20434 32292 20434 0 _0878_
rlabel metal1 32246 25330 32246 25330 0 _0879_
rlabel metal1 33994 23732 33994 23732 0 _0880_
rlabel metal2 35006 16218 35006 16218 0 _0881_
rlabel metal1 33258 23698 33258 23698 0 _0882_
rlabel via1 36202 17646 36202 17646 0 _0883_
rlabel metal1 36754 19754 36754 19754 0 _0884_
rlabel metal1 34730 23800 34730 23800 0 _0885_
rlabel metal1 38594 20842 38594 20842 0 _0886_
rlabel metal1 39146 18802 39146 18802 0 _0887_
rlabel metal2 33074 23324 33074 23324 0 _0888_
rlabel metal1 33534 28390 33534 28390 0 _0889_
rlabel metal2 32890 22780 32890 22780 0 _0890_
rlabel metal1 38042 22440 38042 22440 0 _0891_
rlabel metal1 31648 26554 31648 26554 0 _0892_
rlabel metal1 31188 19822 31188 19822 0 _0893_
rlabel metal1 33488 23630 33488 23630 0 _0894_
rlabel metal2 37582 28016 37582 28016 0 _0895_
rlabel metal2 37490 27132 37490 27132 0 _0896_
rlabel metal1 33718 16082 33718 16082 0 _0897_
rlabel metal1 36892 23018 36892 23018 0 _0898_
rlabel metal2 38042 22780 38042 22780 0 _0899_
rlabel metal1 39100 22406 39100 22406 0 _0900_
rlabel metal1 32062 22474 32062 22474 0 _0901_
rlabel metal1 32982 17816 32982 17816 0 _0902_
rlabel metal1 32614 17646 32614 17646 0 _0903_
rlabel metal1 31326 16014 31326 16014 0 _0904_
rlabel metal1 32798 17680 32798 17680 0 _0905_
rlabel metal1 37766 15470 37766 15470 0 _0906_
rlabel metal1 35558 19346 35558 19346 0 _0907_
rlabel via1 36644 16558 36644 16558 0 _0908_
rlabel metal1 35512 18734 35512 18734 0 _0909_
rlabel metal1 35512 19482 35512 19482 0 _0910_
rlabel metal1 35420 24786 35420 24786 0 _0911_
rlabel metal1 36570 24786 36570 24786 0 _0912_
rlabel metal1 35282 26384 35282 26384 0 _0913_
rlabel metal1 34638 26350 34638 26350 0 _0914_
rlabel metal1 34592 25874 34592 25874 0 _0915_
rlabel metal1 36938 25466 36938 25466 0 _0916_
rlabel metal1 34592 21522 34592 21522 0 _0917_
rlabel metal1 36754 26928 36754 26928 0 _0918_
rlabel metal1 38088 26010 38088 26010 0 _0919_
rlabel metal2 38042 25466 38042 25466 0 _0920_
rlabel metal2 37628 18020 37628 18020 0 _0921_
rlabel metal1 33672 17306 33672 17306 0 _0922_
rlabel metal1 34914 13294 34914 13294 0 _0923_
rlabel metal1 36938 12954 36938 12954 0 _0924_
rlabel metal1 39054 14042 39054 14042 0 _0925_
rlabel metal2 31234 18938 31234 18938 0 _0926_
rlabel metal2 31878 18496 31878 18496 0 _0927_
rlabel metal1 32292 18258 32292 18258 0 _0928_
rlabel metal2 34086 17986 34086 17986 0 _0929_
rlabel metal2 31786 19482 31786 19482 0 _0930_
rlabel metal1 32706 10166 32706 10166 0 _0931_
rlabel metal2 32798 10608 32798 10608 0 _0932_
rlabel metal1 32890 13940 32890 13940 0 _0933_
rlabel metal1 36432 10030 36432 10030 0 _0934_
rlabel metal1 34454 13498 34454 13498 0 _0935_
rlabel metal1 35144 9690 35144 9690 0 _0936_
rlabel metal1 35650 22610 35650 22610 0 _0937_
rlabel metal1 35006 9554 35006 9554 0 _0938_
rlabel metal1 37628 10574 37628 10574 0 _0939_
rlabel metal1 37306 10744 37306 10744 0 _0940_
rlabel metal1 38502 10472 38502 10472 0 _0941_
rlabel metal1 34822 15538 34822 15538 0 _0942_
rlabel metal2 36570 16507 36570 16507 0 _0943_
rlabel metal1 31510 15436 31510 15436 0 _0944_
rlabel metal1 32384 13702 32384 13702 0 _0945_
rlabel metal1 32844 10642 32844 10642 0 _0946_
rlabel metal1 35742 10234 35742 10234 0 _0947_
rlabel metal2 37306 13974 37306 13974 0 _0948_
rlabel metal1 38226 17136 38226 17136 0 _0949_
rlabel metal1 36984 11050 36984 11050 0 _0950_
rlabel metal2 38318 10812 38318 10812 0 _0951_
rlabel metal1 36616 11526 36616 11526 0 _0952_
rlabel metal1 37076 10098 37076 10098 0 _0953_
rlabel metal1 37490 20910 37490 20910 0 _0954_
rlabel metal1 39192 20230 39192 20230 0 _0955_
rlabel metal1 33902 14960 33902 14960 0 _0956_
rlabel metal2 35006 15402 35006 15402 0 _0957_
rlabel metal2 34822 16592 34822 16592 0 _0958_
rlabel metal1 35604 15062 35604 15062 0 _0959_
rlabel metal1 37398 14790 37398 14790 0 _0960_
rlabel metal1 36570 21080 36570 21080 0 _0961_
rlabel metal1 37582 17646 37582 17646 0 _0962_
rlabel metal2 38318 15810 38318 15810 0 _0963_
rlabel metal1 36892 20978 36892 20978 0 _0964_
rlabel metal1 38962 12648 38962 12648 0 _0965_
rlabel metal1 36432 20842 36432 20842 0 _0966_
rlabel metal1 37628 11866 37628 11866 0 _0967_
rlabel metal2 32798 13600 32798 13600 0 _0968_
rlabel metal1 35351 13430 35351 13430 0 _0969_
rlabel metal1 38640 12410 38640 12410 0 _0970_
rlabel metal1 39008 10710 39008 10710 0 _0971_
rlabel metal1 32614 13872 32614 13872 0 _0972_
rlabel metal2 36202 18394 36202 18394 0 _0973_
rlabel metal2 38594 18428 38594 18428 0 _0974_
rlabel metal3 34385 19244 34385 19244 0 _0975_
rlabel metal2 38686 27268 38686 27268 0 _0976_
rlabel metal1 39514 26826 39514 26826 0 _0977_
rlabel metal1 34960 19822 34960 19822 0 _0978_
rlabel via1 36938 19822 36938 19822 0 _0979_
rlabel metal1 38088 18122 38088 18122 0 _0980_
rlabel metal1 38870 18054 38870 18054 0 _0981_
rlabel metal1 39192 13226 39192 13226 0 _0982_
rlabel metal1 38364 13158 38364 13158 0 _0983_
rlabel metal1 36432 16558 36432 16558 0 _0984_
rlabel metal1 37260 16694 37260 16694 0 _0985_
rlabel metal2 38042 10676 38042 10676 0 _0986_
rlabel metal1 38686 15538 38686 15538 0 _0987_
rlabel metal2 37490 14654 37490 14654 0 _0988_
rlabel metal2 38686 15164 38686 15164 0 _0989_
rlabel metal2 38962 11849 38962 11849 0 _0990_
rlabel metal1 39054 11832 39054 11832 0 _0991_
rlabel metal1 39330 24582 39330 24582 0 _0992_
rlabel metal1 36662 15674 36662 15674 0 _0993_
rlabel metal2 38134 17340 38134 17340 0 _0994_
rlabel metal2 33074 16694 33074 16694 0 _0995_
rlabel metal1 36202 17238 36202 17238 0 _0996_
rlabel metal2 38410 18411 38410 18411 0 _0997_
rlabel metal1 38686 22134 38686 22134 0 _0998_
rlabel metal2 38686 22610 38686 22610 0 _0999_
rlabel metal1 37260 24650 37260 24650 0 _1000_
rlabel metal2 37950 24548 37950 24548 0 _1001_
rlabel metal2 36386 25466 36386 25466 0 _1002_
rlabel metal2 33534 24106 33534 24106 0 _1003_
rlabel metal2 37766 24956 37766 24956 0 _1004_
rlabel metal2 36938 14603 36938 14603 0 _1005_
rlabel metal1 37260 13974 37260 13974 0 _1006_
rlabel metal1 36938 13736 36938 13736 0 _1007_
rlabel metal2 34730 13634 34730 13634 0 _1008_
rlabel metal1 35972 13498 35972 13498 0 _1009_
rlabel metal2 18538 12988 18538 12988 0 _1010_
rlabel metal2 19366 14144 19366 14144 0 _1011_
rlabel metal1 17434 12784 17434 12784 0 _1012_
rlabel metal1 17756 12614 17756 12614 0 _1013_
rlabel metal1 21712 20774 21712 20774 0 _1014_
rlabel metal2 20102 14144 20102 14144 0 _1015_
rlabel metal1 17066 12648 17066 12648 0 _1016_
rlabel metal1 16836 7242 16836 7242 0 _1017_
rlabel via1 25072 32402 25072 32402 0 _1018_
rlabel metal2 23598 28866 23598 28866 0 _1019_
rlabel metal1 23506 30906 23506 30906 0 _1020_
rlabel metal2 23414 29818 23414 29818 0 _1021_
rlabel metal2 22494 29002 22494 29002 0 _1022_
rlabel metal1 21436 28730 21436 28730 0 _1023_
rlabel metal1 15088 16082 15088 16082 0 _1024_
rlabel metal1 17342 19482 17342 19482 0 _1025_
rlabel metal1 20470 15470 20470 15470 0 _1026_
rlabel metal1 20654 15436 20654 15436 0 _1027_
rlabel metal2 17802 15096 17802 15096 0 _1028_
rlabel metal2 18078 17102 18078 17102 0 _1029_
rlabel metal1 17894 14926 17894 14926 0 _1030_
rlabel metal2 22218 18428 22218 18428 0 _1031_
rlabel metal1 19918 22168 19918 22168 0 _1032_
rlabel metal2 16882 14722 16882 14722 0 _1033_
rlabel metal1 16054 16116 16054 16116 0 _1034_
rlabel metal2 14766 21760 14766 21760 0 _1035_
rlabel metal1 17664 16558 17664 16558 0 _1036_
rlabel metal1 17526 22066 17526 22066 0 _1037_
rlabel metal2 17986 13651 17986 13651 0 _1038_
rlabel metal2 17710 12274 17710 12274 0 _1039_
rlabel metal2 21666 19108 21666 19108 0 _1040_
rlabel metal1 20746 18938 20746 18938 0 _1041_
rlabel metal1 17618 15470 17618 15470 0 _1042_
rlabel metal2 16238 16660 16238 16660 0 _1043_
rlabel metal2 17066 18904 17066 18904 0 _1044_
rlabel metal2 17526 13090 17526 13090 0 _1045_
rlabel metal2 17066 14212 17066 14212 0 _1046_
rlabel metal1 14950 14960 14950 14960 0 _1047_
rlabel metal1 14444 13362 14444 13362 0 _1048_
rlabel metal1 25020 32538 25020 32538 0 _1049_
rlabel metal1 24058 32878 24058 32878 0 _1050_
rlabel metal2 26450 32606 26450 32606 0 _1051_
rlabel metal1 24334 32300 24334 32300 0 _1052_
rlabel metal1 24012 32402 24012 32402 0 _1053_
rlabel metal1 20148 20026 20148 20026 0 _1054_
rlabel metal1 19550 22202 19550 22202 0 _1055_
rlabel metal1 20010 23494 20010 23494 0 _1056_
rlabel metal1 22494 32436 22494 32436 0 _1057_
rlabel metal1 17204 18190 17204 18190 0 _1058_
rlabel metal2 17020 15028 17020 15028 0 _1059_
rlabel metal1 16238 13396 16238 13396 0 _1060_
rlabel metal1 16054 13158 16054 13158 0 _1061_
rlabel metal1 18216 11118 18216 11118 0 _1062_
rlabel metal1 17434 14450 17434 14450 0 _1063_
rlabel metal1 19274 13260 19274 13260 0 _1064_
rlabel metal1 17388 14382 17388 14382 0 _1065_
rlabel metal1 16376 14314 16376 14314 0 _1066_
rlabel metal1 15548 14518 15548 14518 0 _1067_
rlabel metal1 21298 32334 21298 32334 0 _1068_
rlabel metal1 22724 32266 22724 32266 0 _1069_
rlabel via2 15594 18275 15594 18275 0 _1070_
rlabel metal2 13294 17918 13294 17918 0 _1071_
rlabel metal1 7866 14994 7866 14994 0 _1072_
rlabel metal1 20838 14484 20838 14484 0 _1073_
rlabel via3 21827 26316 21827 26316 0 _1074_
rlabel metal2 22034 15759 22034 15759 0 _1075_
rlabel metal1 18078 26962 18078 26962 0 _1076_
rlabel metal1 12972 32334 12972 32334 0 _1077_
rlabel metal1 28014 10778 28014 10778 0 _1078_
rlabel metal1 26128 11186 26128 11186 0 _1079_
rlabel metal1 24610 11288 24610 11288 0 _1080_
rlabel metal1 22540 9690 22540 9690 0 _1081_
rlabel metal1 21942 10506 21942 10506 0 _1082_
rlabel metal1 21160 11118 21160 11118 0 _1083_
rlabel metal1 22816 23086 22816 23086 0 _1084_
rlabel metal1 21390 11050 21390 11050 0 _1085_
rlabel metal2 21942 10778 21942 10778 0 _1086_
rlabel metal1 22540 10778 22540 10778 0 _1087_
rlabel via2 22494 21981 22494 21981 0 _1088_
rlabel metal2 22218 23834 22218 23834 0 _1089_
rlabel metal1 20286 20944 20286 20944 0 _1090_
rlabel metal1 20102 22508 20102 22508 0 _1091_
rlabel metal1 11178 22644 11178 22644 0 _1092_
rlabel metal1 21344 26350 21344 26350 0 _1093_
rlabel metal1 20976 26418 20976 26418 0 _1094_
rlabel metal2 20470 25126 20470 25126 0 _1095_
rlabel metal2 18354 26758 18354 26758 0 _1096_
rlabel metal2 20102 26758 20102 26758 0 _1097_
rlabel via1 19734 27285 19734 27285 0 _1098_
rlabel metal1 20332 24922 20332 24922 0 _1099_
rlabel metal2 20654 26452 20654 26452 0 _1100_
rlabel metal1 21390 28118 21390 28118 0 _1101_
rlabel metal2 20516 22202 20516 22202 0 _1102_
rlabel metal2 21850 19346 21850 19346 0 _1103_
rlabel metal1 20102 27438 20102 27438 0 _1104_
rlabel metal1 20332 26962 20332 26962 0 _1105_
rlabel metal2 20838 27302 20838 27302 0 _1106_
rlabel metal1 22402 28016 22402 28016 0 _1107_
rlabel metal2 19274 9758 19274 9758 0 _1108_
rlabel metal1 19734 10132 19734 10132 0 _1109_
rlabel metal2 19550 14688 19550 14688 0 _1110_
rlabel metal2 19826 12920 19826 12920 0 _1111_
rlabel metal1 20608 15130 20608 15130 0 _1112_
rlabel metal1 19688 14314 19688 14314 0 _1113_
rlabel via2 19826 14603 19826 14603 0 _1114_
rlabel metal2 19274 27438 19274 27438 0 _1115_
rlabel metal1 19274 26962 19274 26962 0 _1116_
rlabel metal2 17894 27744 17894 27744 0 _1117_
rlabel metal1 19780 27982 19780 27982 0 _1118_
rlabel metal2 18722 27710 18722 27710 0 _1119_
rlabel metal1 17457 28050 17457 28050 0 _1120_
rlabel metal2 18814 27166 18814 27166 0 _1121_
rlabel metal2 16698 27812 16698 27812 0 _1122_
rlabel metal1 16882 15640 16882 15640 0 _1123_
rlabel metal1 17066 17136 17066 17136 0 _1124_
rlabel metal2 16606 17986 16606 17986 0 _1125_
rlabel metal1 16008 18394 16008 18394 0 _1126_
rlabel metal2 15134 26350 15134 26350 0 _1127_
rlabel metal2 11914 25942 11914 25942 0 _1128_
rlabel metal1 15870 26962 15870 26962 0 _1129_
rlabel metal1 16974 28152 16974 28152 0 _1130_
rlabel metal2 16054 26826 16054 26826 0 _1131_
rlabel metal2 18170 27166 18170 27166 0 _1132_
rlabel metal1 17940 26350 17940 26350 0 _1133_
rlabel metal1 14030 25942 14030 25942 0 _1134_
rlabel metal1 12420 25670 12420 25670 0 _1135_
rlabel metal1 10994 27438 10994 27438 0 _1136_
rlabel metal2 12650 27302 12650 27302 0 _1137_
rlabel metal2 18906 27812 18906 27812 0 _1138_
rlabel via1 19191 28934 19191 28934 0 _1139_
rlabel metal1 20194 29206 20194 29206 0 _1140_
rlabel metal2 19550 29376 19550 29376 0 _1141_
rlabel metal1 14628 31994 14628 31994 0 _1142_
rlabel via1 11728 31314 11728 31314 0 _1143_
rlabel metal1 12742 29546 12742 29546 0 _1144_
rlabel metal1 20746 20400 20746 20400 0 _1145_
rlabel metal2 15962 18938 15962 18938 0 _1146_
rlabel metal1 15916 19346 15916 19346 0 _1147_
rlabel metal1 15226 19822 15226 19822 0 _1148_
rlabel metal1 24150 10642 24150 10642 0 _1149_
rlabel metal1 23506 14790 23506 14790 0 _1150_
rlabel metal1 21252 16762 21252 16762 0 _1151_
rlabel metal1 21298 16490 21298 16490 0 _1152_
rlabel via2 22954 16779 22954 16779 0 _1153_
rlabel metal1 22862 17748 22862 17748 0 _1154_
rlabel metal2 22310 16320 22310 16320 0 _1155_
rlabel metal1 22862 16660 22862 16660 0 _1156_
rlabel metal1 22908 16422 22908 16422 0 _1157_
rlabel metal2 21850 23953 21850 23953 0 _1158_
rlabel metal1 14306 20026 14306 20026 0 _1159_
rlabel metal1 14214 20502 14214 20502 0 _1160_
rlabel metal1 28704 21522 28704 21522 0 _1161_
rlabel metal1 26082 20978 26082 20978 0 _1162_
rlabel metal1 29532 20842 29532 20842 0 _1163_
rlabel metal2 29118 20094 29118 20094 0 _1164_
rlabel metal1 26358 20910 26358 20910 0 _1165_
rlabel metal2 15502 20774 15502 20774 0 _1166_
rlabel metal2 18262 11832 18262 11832 0 _1167_
rlabel via2 18722 12733 18722 12733 0 _1168_
rlabel metal2 18354 15878 18354 15878 0 _1169_
rlabel via1 14968 19822 14968 19822 0 _1170_
rlabel metal1 14766 20230 14766 20230 0 _1171_
rlabel metal1 14628 20434 14628 20434 0 _1172_
rlabel metal2 28106 31994 28106 31994 0 _1173_
rlabel metal1 27876 31926 27876 31926 0 _1174_
rlabel metal3 21643 20604 21643 20604 0 _1175_
rlabel metal1 29026 19176 29026 19176 0 _1176_
rlabel metal2 21390 20196 21390 20196 0 _1177_
rlabel metal2 15686 20060 15686 20060 0 _1178_
rlabel metal1 15134 19686 15134 19686 0 _1179_
rlabel metal2 13938 20638 13938 20638 0 _1180_
rlabel metal2 14398 20604 14398 20604 0 _1181_
rlabel metal2 12558 19686 12558 19686 0 _1182_
rlabel metal1 6670 19278 6670 19278 0 _1183_
rlabel metal2 13110 21828 13110 21828 0 _1184_
rlabel metal1 14398 22168 14398 22168 0 _1185_
rlabel viali 12831 21522 12831 21522 0 _1186_
rlabel metal1 12742 20808 12742 20808 0 _1187_
rlabel metal2 13018 20876 13018 20876 0 _1188_
rlabel metal2 13570 21012 13570 21012 0 _1189_
rlabel metal1 10212 20026 10212 20026 0 _1190_
rlabel metal2 10902 21556 10902 21556 0 _1191_
rlabel metal1 11408 21998 11408 21998 0 _1192_
rlabel metal1 11868 23086 11868 23086 0 _1193_
rlabel metal1 27876 12614 27876 12614 0 _1194_
rlabel metal1 26128 21998 26128 21998 0 _1195_
rlabel metal1 26726 16218 26726 16218 0 _1196_
rlabel metal1 28796 18666 28796 18666 0 _1197_
rlabel metal1 26634 20026 26634 20026 0 _1198_
rlabel metal1 27646 19788 27646 19788 0 _1199_
rlabel metal1 28060 19958 28060 19958 0 _1200_
rlabel metal2 28934 24208 28934 24208 0 _1201_
rlabel metal2 28014 20774 28014 20774 0 _1202_
rlabel metal1 28152 16762 28152 16762 0 _1203_
rlabel metal2 27370 19958 27370 19958 0 _1204_
rlabel metal2 27462 19686 27462 19686 0 _1205_
rlabel metal1 27830 20026 27830 20026 0 _1206_
rlabel metal1 27968 20434 27968 20434 0 _1207_
rlabel metal1 27462 19890 27462 19890 0 _1208_
rlabel metal1 24150 14586 24150 14586 0 _1209_
rlabel metal1 26358 18938 26358 18938 0 _1210_
rlabel metal1 26128 25262 26128 25262 0 _1211_
rlabel metal1 25944 26010 25944 26010 0 _1212_
rlabel metal2 20930 9401 20930 9401 0 _1213_
rlabel metal2 26818 26758 26818 26758 0 _1214_
rlabel metal2 23046 28492 23046 28492 0 _1215_
rlabel metal2 23322 27404 23322 27404 0 _1216_
rlabel metal1 23460 26826 23460 26826 0 _1217_
rlabel metal2 17894 28866 17894 28866 0 _1218_
rlabel metal3 23529 20740 23529 20740 0 _1219_
rlabel metal2 24426 21760 24426 21760 0 _1220_
rlabel metal1 25024 26282 25024 26282 0 _1221_
rlabel metal1 24242 26554 24242 26554 0 _1222_
rlabel metal1 25668 29138 25668 29138 0 _1223_
rlabel metal1 25070 26962 25070 26962 0 _1224_
rlabel metal1 24234 28390 24234 28390 0 _1225_
rlabel metal1 17802 28594 17802 28594 0 _1226_
rlabel metal1 16882 29104 16882 29104 0 _1227_
rlabel metal1 17158 28594 17158 28594 0 _1228_
rlabel metal1 16192 24174 16192 24174 0 _1229_
rlabel metal1 19136 19822 19136 19822 0 _1230_
rlabel metal1 18952 24174 18952 24174 0 _1231_
rlabel metal1 20194 24378 20194 24378 0 _1232_
rlabel metal1 17894 29648 17894 29648 0 _1233_
rlabel metal1 15272 29614 15272 29614 0 _1234_
rlabel metal1 13800 29138 13800 29138 0 _1235_
rlabel metal2 11730 28220 11730 28220 0 _1236_
rlabel metal2 9982 18122 9982 18122 0 _1237_
rlabel metal1 11270 11118 11270 11118 0 _1238_
rlabel metal1 10534 11152 10534 11152 0 _1239_
rlabel metal1 13616 13906 13616 13906 0 _1240_
rlabel metal1 19826 32334 19826 32334 0 _1241_
rlabel metal1 19642 31314 19642 31314 0 _1242_
rlabel metal1 17250 21046 17250 21046 0 _1243_
rlabel metal1 17480 19278 17480 19278 0 _1244_
rlabel metal1 15364 17170 15364 17170 0 _1245_
rlabel metal2 9522 16422 9522 16422 0 _1246_
rlabel metal1 16376 14042 16376 14042 0 _1247_
rlabel metal2 16974 16218 16974 16218 0 _1248_
rlabel metal2 17434 15844 17434 15844 0 _1249_
rlabel metal1 16836 15470 16836 15470 0 _1250_
rlabel metal2 16422 15878 16422 15878 0 _1251_
rlabel metal1 15548 16082 15548 16082 0 _1252_
rlabel metal2 14582 16354 14582 16354 0 _1253_
rlabel metal2 12926 10472 12926 10472 0 _1254_
rlabel metal2 14214 7038 14214 7038 0 _1255_
rlabel metal1 14352 16150 14352 16150 0 _1256_
rlabel metal1 11822 16218 11822 16218 0 _1257_
rlabel metal1 18538 23834 18538 23834 0 _1258_
rlabel metal2 17342 24990 17342 24990 0 _1259_
rlabel metal1 26266 31994 26266 31994 0 _1260_
rlabel metal1 25070 27030 25070 27030 0 _1261_
rlabel metal1 24334 24174 24334 24174 0 _1262_
rlabel metal2 18446 20638 18446 20638 0 _1263_
rlabel metal2 23782 24106 23782 24106 0 _1264_
rlabel metal1 23782 24208 23782 24208 0 _1265_
rlabel metal2 24150 25670 24150 25670 0 _1266_
rlabel metal1 23966 26350 23966 26350 0 _1267_
rlabel metal2 23138 25704 23138 25704 0 _1268_
rlabel metal1 24012 27030 24012 27030 0 _1269_
rlabel metal1 17480 25262 17480 25262 0 _1270_
rlabel viali 14489 24174 14489 24174 0 _1271_
rlabel metal1 15870 25466 15870 25466 0 _1272_
rlabel metal1 26680 24378 26680 24378 0 _1273_
rlabel metal1 26358 25228 26358 25228 0 _1274_
rlabel metal2 17434 25092 17434 25092 0 _1275_
rlabel metal2 15502 24956 15502 24956 0 _1276_
rlabel metal2 15962 24072 15962 24072 0 _1277_
rlabel metal1 16054 23698 16054 23698 0 _1278_
rlabel metal2 15502 23936 15502 23936 0 _1279_
rlabel metal1 7222 25228 7222 25228 0 _1280_
rlabel metal1 9522 24752 9522 24752 0 _1281_
rlabel metal1 8280 23698 8280 23698 0 _1282_
rlabel metal1 11316 24786 11316 24786 0 _1283_
rlabel metal1 6486 25942 6486 25942 0 _1284_
rlabel metal1 12236 24786 12236 24786 0 _1285_
rlabel metal2 12558 17714 12558 17714 0 _1286_
rlabel metal2 12006 16524 12006 16524 0 _1287_
rlabel metal1 11500 15878 11500 15878 0 _1288_
rlabel metal2 12374 9316 12374 9316 0 _1289_
rlabel metal1 12742 11016 12742 11016 0 _1290_
rlabel viali 12833 11118 12833 11118 0 _1291_
rlabel metal1 12512 9962 12512 9962 0 _1292_
rlabel metal2 17342 27404 17342 27404 0 _1293_
rlabel metal1 16606 27098 16606 27098 0 _1294_
rlabel metal1 10718 26962 10718 26962 0 _1295_
rlabel metal1 11408 31790 11408 31790 0 _1296_
rlabel metal2 6394 21325 6394 21325 0 _1297_
rlabel metal2 5658 23358 5658 23358 0 _1298_
rlabel metal1 5428 23222 5428 23222 0 _1299_
rlabel metal1 11132 32878 11132 32878 0 _1300_
rlabel metal1 13938 31858 13938 31858 0 _1301_
rlabel metal2 10810 31110 10810 31110 0 _1302_
rlabel metal1 3450 18394 3450 18394 0 _1303_
rlabel metal1 8970 17510 8970 17510 0 _1304_
rlabel metal1 7498 24378 7498 24378 0 _1305_
rlabel metal1 9016 26554 9016 26554 0 _1306_
rlabel metal1 2162 35632 2162 35632 0 _1307_
rlabel metal2 15410 9180 15410 9180 0 _1308_
rlabel metal1 10212 17170 10212 17170 0 _1309_
rlabel metal1 9154 17170 9154 17170 0 _1310_
rlabel metal1 9522 16966 9522 16966 0 _1311_
rlabel metal1 9982 10608 9982 10608 0 _1312_
rlabel metal1 9936 11118 9936 11118 0 _1313_
rlabel metal2 8418 10064 8418 10064 0 _1314_
rlabel metal1 6026 21556 6026 21556 0 _1315_
rlabel metal1 5980 24582 5980 24582 0 _1316_
rlabel metal1 5980 20026 5980 20026 0 _1317_
rlabel metal1 7360 21658 7360 21658 0 _1318_
rlabel metal1 13294 31280 13294 31280 0 _1319_
rlabel metal1 13386 27404 13386 27404 0 _1320_
rlabel metal1 13340 26826 13340 26826 0 _1321_
rlabel metal1 13754 27404 13754 27404 0 _1322_
rlabel metal1 13524 27506 13524 27506 0 _1323_
rlabel metal2 13018 29444 13018 29444 0 _1324_
rlabel metal2 12282 27115 12282 27115 0 _1325_
rlabel metal2 9614 29308 9614 29308 0 _1326_
rlabel metal2 2714 21760 2714 21760 0 _1327_
rlabel metal1 7636 16626 7636 16626 0 _1328_
rlabel metal2 12742 5610 12742 5610 0 _1329_
rlabel metal1 8510 16116 8510 16116 0 _1330_
rlabel via1 8234 16490 8234 16490 0 _1331_
rlabel metal2 6394 25670 6394 25670 0 _1332_
rlabel metal2 7038 25466 7038 25466 0 _1333_
rlabel metal1 7038 17170 7038 17170 0 _1334_
rlabel metal1 7774 16762 7774 16762 0 _1335_
rlabel via2 20838 20859 20838 20859 0 clk
rlabel via2 22034 20757 22034 20757 0 clknet_0_clk
rlabel metal1 12466 7480 12466 7480 0 clknet_4_0_0_clk
rlabel metal1 37490 7922 37490 7922 0 clknet_4_10_0_clk
rlabel metal1 38318 7412 38318 7412 0 clknet_4_11_0_clk
rlabel metal1 17480 33422 17480 33422 0 clknet_4_12_0_clk
rlabel metal1 19826 37910 19826 37910 0 clknet_4_13_0_clk
rlabel metal1 38180 31790 38180 31790 0 clknet_4_14_0_clk
rlabel metal1 29072 34034 29072 34034 0 clknet_4_15_0_clk
rlabel metal1 2162 12886 2162 12886 0 clknet_4_1_0_clk
rlabel metal1 16928 2482 16928 2482 0 clknet_4_2_0_clk
rlabel metal1 14858 18122 14858 18122 0 clknet_4_3_0_clk
rlabel metal1 1656 19278 1656 19278 0 clknet_4_4_0_clk
rlabel metal1 2530 27914 2530 27914 0 clknet_4_5_0_clk
rlabel metal1 5842 31790 5842 31790 0 clknet_4_6_0_clk
rlabel metal1 13018 37706 13018 37706 0 clknet_4_7_0_clk
rlabel metal1 23000 2482 23000 2482 0 clknet_4_8_0_clk
rlabel metal1 17250 18734 17250 18734 0 clknet_4_9_0_clk
rlabel metal2 39698 24021 39698 24021 0 dataBusIn[0]
rlabel metal1 31004 41106 31004 41106 0 dataBusIn[1]
rlabel metal2 40250 24667 40250 24667 0 dataBusIn[2]
rlabel metal3 751 29988 751 29988 0 dataBusIn[3]
rlabel metal2 40250 26775 40250 26775 0 dataBusIn[4]
rlabel metal2 39422 17969 39422 17969 0 dataBusIn[5]
rlabel metal2 39606 27319 39606 27319 0 dataBusIn[6]
rlabel metal1 40112 26350 40112 26350 0 dataBusIn[7]
rlabel metal2 16790 1520 16790 1520 0 dataBusOut[0]
rlabel metal2 16146 1520 16146 1520 0 dataBusOut[1]
rlabel metal2 14214 1520 14214 1520 0 dataBusOut[2]
rlabel metal2 11638 1520 11638 1520 0 dataBusOut[3]
rlabel metal2 13570 1656 13570 1656 0 dataBusOut[4]
rlabel metal2 12926 1656 12926 1656 0 dataBusOut[5]
rlabel metal2 12282 1095 12282 1095 0 dataBusOut[6]
rlabel metal2 14858 1520 14858 1520 0 dataBusOut[7]
rlabel metal2 21298 1520 21298 1520 0 dataBusSelect
rlabel via2 1702 33405 1702 33405 0 gpio[0]
rlabel metal1 24150 37774 24150 37774 0 gpio[10]
rlabel metal1 26542 38386 26542 38386 0 gpio[11]
rlabel metal1 24610 38998 24610 38998 0 gpio[12]
rlabel metal1 25116 35734 25116 35734 0 gpio[13]
rlabel metal1 27784 36210 27784 36210 0 gpio[14]
rlabel metal2 25806 42283 25806 42283 0 gpio[15]
rlabel metal1 15594 3026 15594 3026 0 gpio[16]
rlabel metal2 19366 1588 19366 1588 0 gpio[17]
rlabel metal2 20654 1588 20654 1588 0 gpio[18]
rlabel metal2 23230 1761 23230 1761 0 gpio[19]
rlabel metal2 3266 31008 3266 31008 0 gpio[1]
rlabel metal2 18078 1761 18078 1761 0 gpio[20]
rlabel metal1 34224 29478 34224 29478 0 gpio[21]
rlabel metal2 21942 1860 21942 1860 0 gpio[22]
rlabel metal3 1280 10948 1280 10948 0 gpio[23]
rlabel metal2 23874 1520 23874 1520 0 gpio[24]
rlabel via2 1610 30651 1610 30651 0 gpio[2]
rlabel metal2 1518 32759 1518 32759 0 gpio[3]
rlabel metal2 1702 33983 1702 33983 0 gpio[4]
rlabel metal2 7130 42283 7130 42283 0 gpio[5]
rlabel metal1 1380 34986 1380 34986 0 gpio[6]
rlabel metal2 2990 35870 2990 35870 0 gpio[7]
rlabel metal1 27278 36822 27278 36822 0 gpio[8]
rlabel metal1 26910 38386 26910 38386 0 gpio[9]
rlabel metal2 16882 26367 16882 26367 0 net1
rlabel metal1 16974 2414 16974 2414 0 net10
rlabel metal1 37260 8942 37260 8942 0 net100
rlabel metal1 26634 13804 26634 13804 0 net101
rlabel metal2 26910 9520 26910 9520 0 net102
rlabel metal1 37490 8942 37490 8942 0 net103
rlabel metal1 35282 7956 35282 7956 0 net104
rlabel metal2 18032 19244 18032 19244 0 net105
rlabel via2 22770 23715 22770 23715 0 net106
rlabel metal1 19734 17136 19734 17136 0 net107
rlabel metal1 21298 8534 21298 8534 0 net108
rlabel metal2 24518 15504 24518 15504 0 net109
rlabel metal1 15916 2414 15916 2414 0 net11
rlabel metal1 29532 7514 29532 7514 0 net110
rlabel metal1 17710 19448 17710 19448 0 net111
rlabel metal2 28750 19142 28750 19142 0 net112
rlabel metal1 25668 30022 25668 30022 0 net113
rlabel metal2 18538 21495 18538 21495 0 net114
rlabel metal1 25668 27370 25668 27370 0 net115
rlabel metal1 20654 8534 20654 8534 0 net116
rlabel metal1 17894 8976 17894 8976 0 net117
rlabel metal2 18998 12036 18998 12036 0 net118
rlabel metal1 23920 19278 23920 19278 0 net119
rlabel metal1 14076 4590 14076 4590 0 net12
rlabel metal2 19274 18292 19274 18292 0 net120
rlabel metal1 29762 12818 29762 12818 0 net121
rlabel metal1 29716 19822 29716 19822 0 net122
rlabel metal1 21482 29070 21482 29070 0 net123
rlabel metal1 23046 27506 23046 27506 0 net124
rlabel metal1 30636 27098 30636 27098 0 net125
rlabel metal1 27554 30736 27554 30736 0 net126
rlabel metal2 29026 20604 29026 20604 0 net127
rlabel metal1 22816 30294 22816 30294 0 net128
rlabel metal2 3818 13056 3818 13056 0 net129
rlabel metal1 11776 5542 11776 5542 0 net13
rlabel metal2 4186 12971 4186 12971 0 net130
rlabel metal1 14589 8534 14589 8534 0 net131
rlabel metal2 16790 9690 16790 9690 0 net132
rlabel metal1 17112 6086 17112 6086 0 net133
rlabel metal1 3365 21998 3365 21998 0 net134
rlabel metal2 8234 21692 8234 21692 0 net135
rlabel metal2 2714 34850 2714 34850 0 net136
rlabel metal1 10987 36074 10987 36074 0 net137
rlabel metal1 20109 38998 20109 38998 0 net138
rlabel metal1 19235 33558 19235 33558 0 net139
rlabel metal1 14582 2346 14582 2346 0 net14
rlabel metal1 13846 3502 13846 3502 0 net140
rlabel metal2 21574 3230 21574 3230 0 net141
rlabel metal2 37490 7310 37490 7310 0 net142
rlabel metal1 24663 38930 24663 38930 0 net143
rlabel metal2 39606 23494 39606 23494 0 net144
rlabel metal1 36117 32810 36117 32810 0 net145
rlabel metal1 33120 29614 33120 29614 0 net146
rlabel metal1 37996 19754 37996 19754 0 net147
rlabel metal2 17894 26911 17894 26911 0 net148
rlabel metal1 20424 2618 20424 2618 0 net149
rlabel metal1 13846 2414 13846 2414 0 net15
rlabel metal2 17434 2924 17434 2924 0 net150
rlabel metal1 33304 33558 33304 33558 0 net151
rlabel metal1 20654 31450 20654 31450 0 net152
rlabel metal1 17756 5542 17756 5542 0 net153
rlabel metal1 21620 3706 21620 3706 0 net154
rlabel metal2 21298 4590 21298 4590 0 net155
rlabel metal2 22678 4386 22678 4386 0 net156
rlabel metal1 25438 2890 25438 2890 0 net157
rlabel metal1 26082 3434 26082 3434 0 net158
rlabel metal1 20010 3706 20010 3706 0 net159
rlabel metal2 11638 3366 11638 3366 0 net16
rlabel metal2 19550 4828 19550 4828 0 net160
rlabel metal1 11822 4250 11822 4250 0 net161
rlabel metal2 13018 3740 13018 3740 0 net162
rlabel metal1 8372 20910 8372 20910 0 net163
rlabel metal1 10258 18734 10258 18734 0 net164
rlabel metal1 3450 20026 3450 20026 0 net165
rlabel metal1 8096 18734 8096 18734 0 net166
rlabel metal2 4738 18938 4738 18938 0 net167
rlabel metal1 9844 19822 9844 19822 0 net168
rlabel metal1 5060 20842 5060 20842 0 net169
rlabel metal1 15318 2482 15318 2482 0 net17
rlabel metal2 12834 20672 12834 20672 0 net170
rlabel metal1 6992 18258 6992 18258 0 net171
rlabel metal2 14858 3740 14858 3740 0 net172
rlabel metal1 4554 21658 4554 21658 0 net173
rlabel metal1 18952 4046 18952 4046 0 net174
rlabel metal1 13478 4114 13478 4114 0 net175
rlabel metal1 14766 4692 14766 4692 0 net176
rlabel metal2 17158 3536 17158 3536 0 net177
rlabel metal2 2622 22848 2622 22848 0 net178
rlabel metal1 29348 32946 29348 32946 0 net179
rlabel metal1 21298 2414 21298 2414 0 net18
rlabel metal1 13018 4454 13018 4454 0 net180
rlabel metal2 3910 19584 3910 19584 0 net181
rlabel metal1 4416 17578 4416 17578 0 net182
rlabel metal1 12190 6290 12190 6290 0 net183
rlabel metal1 5290 21658 5290 21658 0 net184
rlabel metal1 3404 18258 3404 18258 0 net185
rlabel metal2 31878 32028 31878 32028 0 net186
rlabel metal2 12742 18496 12742 18496 0 net187
rlabel metal1 5244 25262 5244 25262 0 net188
rlabel metal1 8326 25160 8326 25160 0 net189
rlabel metal2 19274 37553 19274 37553 0 net19
rlabel metal1 29440 33558 29440 33558 0 net190
rlabel metal1 13524 23086 13524 23086 0 net191
rlabel metal1 18722 31246 18722 31246 0 net192
rlabel metal1 2944 23834 2944 23834 0 net193
rlabel metal1 3450 26282 3450 26282 0 net194
rlabel metal1 5336 23834 5336 23834 0 net195
rlabel metal1 9936 21658 9936 21658 0 net196
rlabel metal1 35834 31858 35834 31858 0 net197
rlabel metal1 3404 24922 3404 24922 0 net198
rlabel metal1 30636 33490 30636 33490 0 net199
rlabel metal2 16146 32164 16146 32164 0 net2
rlabel metal1 14996 37842 14996 37842 0 net20
rlabel metal1 8372 28526 8372 28526 0 net200
rlabel metal1 14812 12206 14812 12206 0 net201
rlabel metal2 30314 30396 30314 30396 0 net202
rlabel metal1 37490 20502 37490 20502 0 net21
rlabel metal1 6762 34612 6762 34612 0 net22
rlabel metal2 12282 39440 12282 39440 0 net23
rlabel metal1 13386 39916 13386 39916 0 net24
rlabel metal1 16238 39984 16238 39984 0 net25
rlabel metal1 16468 39406 16468 39406 0 net26
rlabel metal1 9246 35632 9246 35632 0 net27
rlabel metal1 13616 15130 13616 15130 0 net28
rlabel metal1 31924 30294 31924 30294 0 net29
rlabel via2 15502 29699 15502 29699 0 net3
rlabel metal1 13754 30702 13754 30702 0 net30
rlabel metal3 11638 31756 11638 31756 0 net31
rlabel metal1 7498 12818 7498 12818 0 net32
rlabel metal1 14260 12818 14260 12818 0 net33
rlabel metal2 35558 9452 35558 9452 0 net34
rlabel metal1 36478 14348 36478 14348 0 net35
rlabel metal1 32890 20400 32890 20400 0 net36
rlabel metal1 35604 20774 35604 20774 0 net37
rlabel metal2 32246 20570 32246 20570 0 net38
rlabel metal1 34459 23630 34459 23630 0 net39
rlabel metal1 15226 30260 15226 30260 0 net4
rlabel metal2 36570 21726 36570 21726 0 net40
rlabel metal2 32614 27693 32614 27693 0 net41
rlabel metal1 39514 29648 39514 29648 0 net42
rlabel metal2 32384 32742 32384 32742 0 net43
rlabel metal1 34776 18802 34776 18802 0 net44
rlabel metal2 10718 28730 10718 28730 0 net45
rlabel metal2 14214 36958 14214 36958 0 net46
rlabel metal1 19642 35190 19642 35190 0 net47
rlabel metal2 15778 19635 15778 19635 0 net48
rlabel metal1 19458 13906 19458 13906 0 net49
rlabel metal1 38134 29546 38134 29546 0 net5
rlabel metal1 19780 20910 19780 20910 0 net50
rlabel metal1 31970 26996 31970 26996 0 net51
rlabel metal3 32775 24956 32775 24956 0 net52
rlabel metal1 14490 19278 14490 19278 0 net53
rlabel metal1 38732 19142 38732 19142 0 net54
rlabel metal1 30406 26860 30406 26860 0 net55
rlabel metal3 21689 19924 21689 19924 0 net56
rlabel metal2 21482 7038 21482 7038 0 net57
rlabel metal2 15318 13804 15318 13804 0 net58
rlabel metal1 16606 18258 16606 18258 0 net59
rlabel metal1 38870 19788 38870 19788 0 net6
rlabel metal1 21482 8262 21482 8262 0 net60
rlabel metal2 32062 27353 32062 27353 0 net61
rlabel metal1 37168 27506 37168 27506 0 net62
rlabel metal2 17802 18292 17802 18292 0 net63
rlabel via1 17615 19346 17615 19346 0 net64
rlabel metal1 18354 20910 18354 20910 0 net65
rlabel metal1 18078 20774 18078 20774 0 net66
rlabel metal1 21574 27948 21574 27948 0 net67
rlabel metal1 17158 21556 17158 21556 0 net68
rlabel metal1 20930 2346 20930 2346 0 net69
rlabel via1 17249 26962 17249 26962 0 net7
rlabel metal1 21436 26894 21436 26894 0 net70
rlabel metal1 26956 31314 26956 31314 0 net71
rlabel metal1 20240 14382 20240 14382 0 net72
rlabel metal1 21758 30634 21758 30634 0 net73
rlabel metal1 20408 8874 20408 8874 0 net74
rlabel metal2 21252 13294 21252 13294 0 net75
rlabel metal2 18722 14654 18722 14654 0 net76
rlabel metal1 34730 19414 34730 19414 0 net77
rlabel metal2 30314 19380 30314 19380 0 net78
rlabel metal1 19136 16966 19136 16966 0 net79
rlabel metal1 36294 26928 36294 26928 0 net8
rlabel metal1 30498 19278 30498 19278 0 net80
rlabel metal1 33534 21556 33534 21556 0 net81
rlabel metal2 32798 20162 32798 20162 0 net82
rlabel metal2 21022 8874 21022 8874 0 net83
rlabel metal1 20976 22746 20976 22746 0 net84
rlabel metal1 30314 23052 30314 23052 0 net85
rlabel metal1 25070 18938 25070 18938 0 net86
rlabel metal2 33902 20264 33902 20264 0 net87
rlabel metal2 20838 8772 20838 8772 0 net88
rlabel metal1 20562 14790 20562 14790 0 net89
rlabel metal1 20470 4998 20470 4998 0 net9
rlabel metal2 35742 21284 35742 21284 0 net90
rlabel metal1 35604 8942 35604 8942 0 net91
rlabel metal1 28980 10234 28980 10234 0 net92
rlabel metal1 31142 9520 31142 9520 0 net93
rlabel metal1 37582 9894 37582 9894 0 net94
rlabel metal1 28888 10030 28888 10030 0 net95
rlabel metal1 30728 9554 30728 9554 0 net96
rlabel metal2 36202 8738 36202 8738 0 net97
rlabel metal2 26450 10370 26450 10370 0 net98
rlabel metal1 31188 9622 31188 9622 0 net99
rlabel via2 40158 3451 40158 3451 0 nrst
rlabel metal2 21390 21913 21390 21913 0 top8227.PSRCurrentValue\[0\]
rlabel metal2 14122 7905 14122 7905 0 top8227.PSRCurrentValue\[1\]
rlabel metal2 16284 19482 16284 19482 0 top8227.PSRCurrentValue\[2\]
rlabel metal2 14904 17204 14904 17204 0 top8227.PSRCurrentValue\[3\]
rlabel via2 16882 10251 16882 10251 0 top8227.PSRCurrentValue\[6\]
rlabel via2 16422 6443 16422 6443 0 top8227.PSRCurrentValue\[7\]
rlabel metal2 19090 25602 19090 25602 0 top8227.branchBackward
rlabel metal1 19918 30770 19918 30770 0 top8227.branchForward
rlabel metal2 31418 33660 31418 33660 0 top8227.demux.isAddressing
rlabel metal1 19228 4182 19228 4182 0 top8227.demux.nmi
rlabel metal2 20654 7378 20654 7378 0 top8227.demux.reset
rlabel metal1 20884 7378 20884 7378 0 top8227.demux.setInterruptFlag
rlabel metal1 33925 33082 33925 33082 0 top8227.demux.state_machine.currentAddress\[0\]
rlabel metal1 34730 32198 34730 32198 0 top8227.demux.state_machine.currentAddress\[10\]
rlabel metal1 29716 31790 29716 31790 0 top8227.demux.state_machine.currentAddress\[11\]
rlabel metal1 34730 32946 34730 32946 0 top8227.demux.state_machine.currentAddress\[12\]
rlabel metal1 39422 31450 39422 31450 0 top8227.demux.state_machine.currentAddress\[1\]
rlabel metal1 32154 29240 32154 29240 0 top8227.demux.state_machine.currentAddress\[2\]
rlabel metal1 28750 33422 28750 33422 0 top8227.demux.state_machine.currentAddress\[3\]
rlabel metal1 35512 31314 35512 31314 0 top8227.demux.state_machine.currentAddress\[4\]
rlabel metal1 29026 30158 29026 30158 0 top8227.demux.state_machine.currentAddress\[5\]
rlabel metal1 38640 29546 38640 29546 0 top8227.demux.state_machine.currentAddress\[6\]
rlabel metal1 38410 28628 38410 28628 0 top8227.demux.state_machine.currentAddress\[7\]
rlabel metal2 34086 33660 34086 33660 0 top8227.demux.state_machine.currentAddress\[8\]
rlabel metal1 31602 32232 31602 32232 0 top8227.demux.state_machine.currentAddress\[9\]
rlabel metal1 40020 7514 40020 7514 0 top8227.demux.state_machine.currentInstruction\[0\]
rlabel metal2 37950 9418 37950 9418 0 top8227.demux.state_machine.currentInstruction\[1\]
rlabel metal1 28842 9520 28842 9520 0 top8227.demux.state_machine.currentInstruction\[2\]
rlabel metal2 33350 8330 33350 8330 0 top8227.demux.state_machine.currentInstruction\[3\]
rlabel metal1 33994 6936 33994 6936 0 top8227.demux.state_machine.currentInstruction\[4\]
rlabel via2 21114 7395 21114 7395 0 top8227.demux.state_machine.currentInstruction\[5\]
rlabel metal1 29992 19890 29992 19890 0 top8227.demux.state_machine.timeState\[0\]
rlabel metal1 23230 17544 23230 17544 0 top8227.demux.state_machine.timeState\[1\]
rlabel metal2 28382 18615 28382 18615 0 top8227.demux.state_machine.timeState\[2\]
rlabel metal4 36156 14416 36156 14416 0 top8227.demux.state_machine.timeState\[3\]
rlabel metal1 29670 18700 29670 18700 0 top8227.demux.state_machine.timeState\[4\]
rlabel metal2 25438 5950 25438 5950 0 top8227.demux.state_machine.timeState\[5\]
rlabel metal1 26910 5338 26910 5338 0 top8227.demux.state_machine.timeState\[6\]
rlabel metal1 21436 31858 21436 31858 0 top8227.freeCarry
rlabel metal1 18860 2958 18860 2958 0 top8227.instructionLoader.interruptInjector.interruptRequest
rlabel metal1 21344 4794 21344 4794 0 top8227.instructionLoader.interruptInjector.irqGenerated
rlabel metal2 21666 3332 21666 3332 0 top8227.instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ
rlabel metal1 19918 2482 19918 2482 0 top8227.instructionLoader.interruptInjector.irqSync.nextQ2
rlabel metal1 19826 4794 19826 4794 0 top8227.instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning
rlabel metal1 19090 2618 19090 2618 0 top8227.instructionLoader.interruptInjector.nmiGeneratedFF.synchronizedNMI
rlabel metal2 15778 3264 15778 3264 0 top8227.instructionLoader.interruptInjector.nmiSync.in
rlabel metal1 17664 3570 17664 3570 0 top8227.instructionLoader.interruptInjector.nmiSync.nextQ2
rlabel via2 29210 5219 29210 5219 0 top8227.instructionLoader.interruptInjector.resetDetected
rlabel metal1 14490 19210 14490 19210 0 top8227.internalDataflow.accRegToDB\[0\]
rlabel metal1 12926 28016 12926 28016 0 top8227.internalDataflow.accRegToDB\[1\]
rlabel metal1 6854 27914 6854 27914 0 top8227.internalDataflow.accRegToDB\[2\]
rlabel metal1 13662 28084 13662 28084 0 top8227.internalDataflow.accRegToDB\[3\]
rlabel metal2 6210 28866 6210 28866 0 top8227.internalDataflow.accRegToDB\[4\]
rlabel metal1 6026 27574 6026 27574 0 top8227.internalDataflow.accRegToDB\[5\]
rlabel metal2 16054 28526 16054 28526 0 top8227.internalDataflow.accRegToDB\[6\]
rlabel metal1 8786 27472 8786 27472 0 top8227.internalDataflow.accRegToDB\[7\]
rlabel metal1 15134 37774 15134 37774 0 top8227.internalDataflow.addressHighBusModule.busInputs\[16\]
rlabel metal1 15502 35564 15502 35564 0 top8227.internalDataflow.addressHighBusModule.busInputs\[17\]
rlabel metal1 15318 37808 15318 37808 0 top8227.internalDataflow.addressHighBusModule.busInputs\[18\]
rlabel via1 15870 39389 15870 39389 0 top8227.internalDataflow.addressHighBusModule.busInputs\[19\]
rlabel metal1 19550 37774 19550 37774 0 top8227.internalDataflow.addressHighBusModule.busInputs\[20\]
rlabel metal1 16008 31314 16008 31314 0 top8227.internalDataflow.addressHighBusModule.busInputs\[21\]
rlabel metal1 19320 34578 19320 34578 0 top8227.internalDataflow.addressHighBusModule.busInputs\[22\]
rlabel metal2 18170 32708 18170 32708 0 top8227.internalDataflow.addressHighBusModule.busInputs\[23\]
rlabel metal1 16284 33830 16284 33830 0 top8227.internalDataflow.addressLowBusModule.busInputs\[16\]
rlabel metal1 13294 34442 13294 34442 0 top8227.internalDataflow.addressLowBusModule.busInputs\[17\]
rlabel metal2 9614 34034 9614 34034 0 top8227.internalDataflow.addressLowBusModule.busInputs\[18\]
rlabel metal2 8510 34238 8510 34238 0 top8227.internalDataflow.addressLowBusModule.busInputs\[19\]
rlabel metal1 4830 35258 4830 35258 0 top8227.internalDataflow.addressLowBusModule.busInputs\[20\]
rlabel metal1 8050 37638 8050 37638 0 top8227.internalDataflow.addressLowBusModule.busInputs\[21\]
rlabel metal2 10258 36890 10258 36890 0 top8227.internalDataflow.addressLowBusModule.busInputs\[22\]
rlabel metal1 12788 25874 12788 25874 0 top8227.internalDataflow.addressLowBusModule.busInputs\[23\]
rlabel metal2 13984 18156 13984 18156 0 top8227.internalDataflow.addressLowBusModule.busInputs\[24\]
rlabel metal1 4692 12614 4692 12614 0 top8227.internalDataflow.addressLowBusModule.busInputs\[25\]
rlabel metal2 6578 17000 6578 17000 0 top8227.internalDataflow.addressLowBusModule.busInputs\[26\]
rlabel metal2 6210 17697 6210 17697 0 top8227.internalDataflow.addressLowBusModule.busInputs\[27\]
rlabel metal1 6210 16218 6210 16218 0 top8227.internalDataflow.addressLowBusModule.busInputs\[28\]
rlabel metal1 5612 19822 5612 19822 0 top8227.internalDataflow.addressLowBusModule.busInputs\[29\]
rlabel metal2 5750 10217 5750 10217 0 top8227.internalDataflow.addressLowBusModule.busInputs\[30\]
rlabel metal2 10718 18972 10718 18972 0 top8227.internalDataflow.addressLowBusModule.busInputs\[31\]
rlabel metal1 13570 21590 13570 21590 0 top8227.internalDataflow.addressLowBusModule.busInputs\[32\]
rlabel metal2 9430 25058 9430 25058 0 top8227.internalDataflow.addressLowBusModule.busInputs\[33\]
rlabel metal1 6256 24242 6256 24242 0 top8227.internalDataflow.addressLowBusModule.busInputs\[34\]
rlabel metal1 4462 25228 4462 25228 0 top8227.internalDataflow.addressLowBusModule.busInputs\[35\]
rlabel metal1 5566 26010 5566 26010 0 top8227.internalDataflow.addressLowBusModule.busInputs\[36\]
rlabel metal2 4370 26180 4370 26180 0 top8227.internalDataflow.addressLowBusModule.busInputs\[37\]
rlabel metal1 3956 24718 3956 24718 0 top8227.internalDataflow.addressLowBusModule.busInputs\[38\]
rlabel metal1 9246 21862 9246 21862 0 top8227.internalDataflow.addressLowBusModule.busInputs\[39\]
rlabel metal1 15870 7786 15870 7786 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[0\]
rlabel metal1 13156 6970 13156 6970 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[1\]
rlabel metal2 19366 6766 19366 6766 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[2\]
rlabel metal1 15364 8534 15364 8534 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[3\]
rlabel metal1 15548 9690 15548 9690 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[6\]
rlabel metal2 12650 19380 12650 19380 0 top8227.internalDataflow.stackBusModule.busInputs\[32\]
rlabel metal1 8574 19890 8574 19890 0 top8227.internalDataflow.stackBusModule.busInputs\[33\]
rlabel metal1 5842 19380 5842 19380 0 top8227.internalDataflow.stackBusModule.busInputs\[34\]
rlabel metal1 4278 19822 4278 19822 0 top8227.internalDataflow.stackBusModule.busInputs\[35\]
rlabel metal1 7360 18598 7360 18598 0 top8227.internalDataflow.stackBusModule.busInputs\[36\]
rlabel metal2 5290 18700 5290 18700 0 top8227.internalDataflow.stackBusModule.busInputs\[37\]
rlabel metal1 5198 19278 5198 19278 0 top8227.internalDataflow.stackBusModule.busInputs\[38\]
rlabel metal1 10488 19482 10488 19482 0 top8227.internalDataflow.stackBusModule.busInputs\[39\]
rlabel metal1 13064 20978 13064 20978 0 top8227.internalDataflow.stackBusModule.busInputs\[40\]
rlabel metal2 8602 21794 8602 21794 0 top8227.internalDataflow.stackBusModule.busInputs\[41\]
rlabel metal1 5152 22542 5152 22542 0 top8227.internalDataflow.stackBusModule.busInputs\[42\]
rlabel metal1 5796 21998 5796 21998 0 top8227.internalDataflow.stackBusModule.busInputs\[43\]
rlabel metal1 5934 20876 5934 20876 0 top8227.internalDataflow.stackBusModule.busInputs\[44\]
rlabel metal2 3634 20332 3634 20332 0 top8227.internalDataflow.stackBusModule.busInputs\[45\]
rlabel metal1 4324 23154 4324 23154 0 top8227.internalDataflow.stackBusModule.busInputs\[46\]
rlabel metal2 10626 20706 10626 20706 0 top8227.internalDataflow.stackBusModule.busInputs\[47\]
rlabel metal1 18492 5338 18492 5338 0 top8227.negEdgeDetector.q1
rlabel metal1 24380 3094 24380 3094 0 top8227.pulse_slower.currentEnableState\[0\]
rlabel metal2 24334 3196 24334 3196 0 top8227.pulse_slower.currentEnableState\[1\]
rlabel metal1 23230 2414 23230 2414 0 top8227.pulse_slower.nextEnableState\[0\]
rlabel metal1 26312 3162 26312 3162 0 top8227.pulse_slower.nextEnableState\[1\]
<< properties >>
string FIXED_BBOX 0 0 41757 43901
<< end >>

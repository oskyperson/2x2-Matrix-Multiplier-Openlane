* NGSPICE file created from matrix_multiplier.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

.subckt matrix_multiplier VGND VPWR cs hz100 miso mosi ready spi_clk
X_3155_ net127 net116 VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__and2_1
X_3086_ net585 net73 net25 VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__mux2_1
XFILLER_54_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2106_ net240 net242 net249 VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__and3_1
X_2037_ _0837_ _0839_ _0828_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_37_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2939_ net460 net87 net40 VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold340 matmult_inst.alu_inst.adder_inst.r3.fa1.a VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold351 matmult_inst.alu_inst.adder_inst.r0.fa2.a VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_12_hz100 clknet_2_3__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_12_hz100
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_79_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_hz100 clknet_2_0__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_27_hz100
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_48_Left_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2724_ _1438_ _1465_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__xor2_1
X_2655_ _1398_ _1399_ _1387_ VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__a21o_1
X_2586_ _1332_ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__inv_2
Xfanout127 _0546_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__buf_2
Xfanout116 net126 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__buf_2
XFILLER_67_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3207_ net131 net120 VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__and2_1
X_3138_ net129 net119 VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__and2_1
X_3069_ net393 net71 net28 VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__mux2_1
XFILLER_23_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold170 matmult_inst.mem_inst.matrixB0\[5\] VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 matmult_inst.alu_inst.out\[13\] VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 matmult_inst.mem_inst.matrixA1\[0\] VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2440_ net228 net226 net208 net209 VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__nand4_2
X_2371_ _1155_ net588 _1152_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2707_ _1412_ _1449_ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__xnor2_1
X_2638_ net222 net202 _1347_ _1349_ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__a22oi_1
X_2569_ net209 net220 net218 net212 VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__a22o_1
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1940_ matmult_inst.spi_inst.tx_reg_sys\[6\] matmult_inst.spi_inst.miso_shifter\[5\]
+ net276 VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__mux2_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1871_ net271 net263 matmult_inst.mem_inst.mem3\[0\] VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__and3_1
X_3610_ clknet_leaf_19_hz100 _0470_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA3\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_3541_ clknet_leaf_26_hz100 _0401_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA0\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3472_ clknet_leaf_8_hz100 _0332_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem0\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_2423_ _1168_ _1174_ net161 VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__o21ai_1
X_2354_ _0791_ _1142_ net199 VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__o21ba_1
X_2285_ _1057_ _1079_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__nand2_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire111 _1107_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_1
Xwire100 net102 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2070_ _0853_ _0854_ _0855_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__o21ai_2
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2972_ net320 net73 net37 VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__mux2_1
X_1923_ _0766_ _0784_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__nor2_1
X_1854_ net267 net260 matmult_inst.mem_inst.matrixA3\[2\] VGND VGND VPWR VPWR _0727_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_12_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1785_ matmult_inst.mem_inst.matrixB2\[8\] net191 net183 matmult_inst.mem_inst.matrixB1\[8\]
+ _0663_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__a221o_1
X_3524_ clknet_leaf_24_hz100 _0384_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem3\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3455_ clknet_leaf_30_hz100 _0315_ VGND VGND VPWR VPWR matmult_inst.alu_inst.a0_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2406_ _1156_ net579 net64 VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__mux2_1
X_3386_ clknet_leaf_29_hz100 _0248_ VGND VGND VPWR VPWR matmult_inst.alu_inst.col0\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2337_ net636 _1129_ net159 VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__mux2_1
XFILLER_57_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2268_ _1042_ _1063_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2199_ _0960_ _0962_ _0995_ _0959_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__a211o_1
XFILLER_52_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold30 matmult_inst.mem_inst.matrixB3\[15\] VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold41 matmult_inst.spi_inst.mosi_data_sync\[6\] VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 matmult_inst.mem_inst.matrixB1\[6\] VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 matmult_inst.alu_inst.out\[6\] VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 matmult_inst.mem_inst.matrixB0\[17\] VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold96 matmult_inst.mem_inst.matrixA3\[2\] VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 matmult_inst.alu_inst.row1\[5\] VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3240_ clknet_leaf_26_hz100 net451 VGND VGND VPWR VPWR matmult_inst.fsm_inst.alu_result\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_3171_ net136 net124 VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__and2_1
XFILLER_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2122_ _0919_ _0921_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__xor2_1
XFILLER_81_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2053_ net241 net254 net252 net243 VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__a22o_1
XFILLER_19_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2955_ net507 net71 net40 VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__mux2_1
X_1906_ _0542_ _0544_ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__or2_1
X_2886_ _0541_ _0775_ VGND VGND VPWR VPWR _1573_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_60_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1837_ net635 _0711_ net91 VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__mux2_1
X_1768_ net287 _0646_ _0648_ net279 VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__a22o_1
X_3507_ clknet_leaf_18_hz100 _0367_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem2\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1699_ matmult_inst.mem_inst.matrixB2\[16\] net191 net183 matmult_inst.mem_inst.matrixB1\[16\]
+ _0585_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__a221o_1
X_3438_ clknet_leaf_7_hz100 _0298_ VGND VGND VPWR VPWR matmult_inst.alu_inst.out\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3369_ clknet_leaf_25_hz100 _0004_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.rx_ready_edge
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_68_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2740_ net644 net160 _1475_ _1479_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__o22a_1
X_2671_ _1413_ _1414_ VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__nor2_1
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1622_ _0538_ _0539_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__or2_2
X_3223_ clknet_leaf_24_hz100 _0001_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.sel\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3154_ net127 net116 VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__and2_1
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3085_ net546 net74 net25 VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__mux2_1
X_2105_ net240 net250 net249 net242 VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__a22oi_2
X_2036_ net239 net258 net255 net241 VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__nand4_1
X_2938_ net277 net186 net88 VGND VGND VPWR VPWR _1585_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2869_ net220 net302 net93 VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__mux2_1
Xhold352 matmult_inst.alu_inst.adder_inst.r0.fa0.a VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold330 matmult_inst.alu_inst.adder_inst.r2.fa0.b VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 matmult_inst.spi_inst.tx_reg_sys\[4\] VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_8_hz100 clknet_2_3__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_8_hz100
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire19 _1536_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_62_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2723_ _1463_ _1464_ VGND VGND VPWR VPWR _1465_ sky130_fd_sc_hd__nor2_1
X_2654_ _1388_ _1395_ _1396_ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__or3_1
X_2585_ _1328_ _1329_ _1330_ net106 VGND VGND VPWR VPWR _1332_ sky130_fd_sc_hd__a22oi_2
Xfanout128 _0546_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__buf_1
Xfanout117 _0553_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3206_ net292 VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__inv_2
X_3137_ net129 net119 VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__and2_1
X_3068_ net512 net72 net27 VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__mux2_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2019_ net259 net243 net244 net256 VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold160 matmult_inst.mem_inst.matrixA0\[1\] VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 matmult_inst.mem_inst.mem2\[4\] VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 matmult_inst.alu_inst.out\[11\] VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 _0136_ VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2370_ _0731_ net167 VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__and2_2
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2706_ _1447_ _1448_ VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2637_ net631 _1382_ net159 VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__mux2_1
X_2568_ _1313_ _1314_ VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__nor2_1
X_2499_ net218 net215 VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__nand2_1
XFILLER_55_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Left_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_11_hz100 clknet_2_3__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_11_hz100
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_11_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_26_hz100 clknet_2_0__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_26_hz100
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_76_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1870_ net637 _0741_ net92 VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__mux2_1
X_3540_ clknet_leaf_17_hz100 _0400_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA0\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3471_ clknet_leaf_18_hz100 _0331_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem0\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2422_ _1168_ _1174_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__and2_1
X_2353_ net177 _0775_ net267 net166 VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__o211a_1
X_2284_ _1077_ _1078_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1999_ matmult_inst.fsm_inst.alu_result\[10\] net114 VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__and2_1
X_3669_ clknet_leaf_28_hz100 _0529_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.state\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_69_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire156 _0540_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__buf_1
XFILLER_50_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2971_ net584 net74 net37 VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__mux2_1
X_1922_ matmult_inst.fsm_inst.rx_ready_edge_delay _0537_ _0551_ _0771_ VGND VGND VPWR
+ VPWR _0790_ sky130_fd_sc_hd__nor4_1
X_1853_ matmult_inst.mem_inst.matrixB2\[2\] net186 net178 matmult_inst.mem_inst.matrixB1\[2\]
+ _0725_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_12_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1784_ net273 net265 matmult_inst.mem_inst.matrixB3\[8\] VGND VGND VPWR VPWR _0663_
+ sky130_fd_sc_hd__and3_1
X_3523_ clknet_leaf_24_hz100 _0383_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem3\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3454_ clknet_leaf_30_hz100 _0314_ VGND VGND VPWR VPWR matmult_inst.alu_inst.a0_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_2405_ _1155_ net386 _1165_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__mux2_1
X_3385_ clknet_leaf_29_hz100 _0247_ VGND VGND VPWR VPWR matmult_inst.alu_inst.col0\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2336_ _1125_ _1128_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__xnor2_1
X_2267_ _1058_ _1060_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__xnor2_1
X_2198_ _0991_ _0992_ _0994_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__a21o_1
XFILLER_65_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold20 matmult_inst.mem_inst.matrixB3\[2\] VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 matmult_inst.mem_inst.matrixB3\[0\] VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold53 _0129_ VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 matmult_inst.mem_inst.matrixB0\[7\] VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 _0165_ VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 matmult_inst.mem_inst.mem1\[15\] VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold86 matmult_inst.alu_inst.out\[3\] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 matmult_inst.alu_inst.out\[9\] VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3170_ net136 net125 VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__and2_1
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2121_ _0883_ _0920_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__nand2_1
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2052_ net241 net243 net254 net252 VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__and4_1
XFILLER_81_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2954_ net433 net72 net39 VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__mux2_1
X_1905_ _0542_ _0544_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__nor2_1
X_2885_ net152 _1569_ VGND VGND VPWR VPWR _1572_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_60_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1836_ matmult_inst.mem_inst.matrixA0\[4\] net169 _0709_ _0710_ VGND VGND VPWR VPWR
+ _0711_ sky130_fd_sc_hd__a211o_1
X_1767_ matmult_inst.mem_inst.mem2\[10\] net188 net180 matmult_inst.mem_inst.mem1\[10\]
+ _0647_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__a221o_1
X_3506_ clknet_leaf_24_hz100 _0366_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem2\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1698_ net272 net264 matmult_inst.mem_inst.matrixB3\[16\] VGND VGND VPWR VPWR _0585_
+ sky130_fd_sc_hd__and3_1
X_3437_ clknet_leaf_7_hz100 _0297_ VGND VGND VPWR VPWR matmult_inst.alu_inst.out\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_3368_ clknet_leaf_30_hz100 _0232_ VGND VGND VPWR VPWR matmult_inst.alu_inst.row0\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2319_ _1066_ _1089_ _1091_ _1088_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__a31o_1
XFILLER_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3299_ clknet_leaf_25_hz100 _0169_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB3\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_68_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2670_ net205 net217 net216 net207 VGND VGND VPWR VPWR _1414_ sky130_fd_sc_hd__a22oi_1
X_1621_ _0538_ _0539_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__nor2_1
X_3222_ clknet_leaf_25_hz100 _0000_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.sel\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3153_ net127 net116 VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2104_ _0902_ _0903_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__or2_1
X_3084_ net396 net75 net25 VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__mux2_1
X_2035_ net238 net258 net255 net241 VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2937_ net447 net70 net42 VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2868_ net221 net513 net93 VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__mux2_1
Xhold320 matmult_inst.alu_inst.adder_inst.r3.fa2.b VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__dlygate4sd3_1
X_2799_ _1511_ _1513_ VGND VGND VPWR VPWR _1514_ sky130_fd_sc_hd__xnor2_1
X_1819_ net281 _0692_ _0694_ net285 VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__a22o_1
Xhold331 matmult_inst.spi_inst.rx_done2 VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 matmult_inst.spi_inst.tx_reg_sys\[15\] VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 matmult_inst.alu_inst.adder_inst.r3.fa1.b VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2722_ _1460_ _1461_ _1462_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__a21oi_1
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2653_ _1395_ _1396_ _1388_ VGND VGND VPWR VPWR _1398_ sky130_fd_sc_hd__o21ai_1
X_2584_ net106 _1328_ _1329_ _1330_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__and4_1
Xfanout118 net121 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
Xfanout129 net132 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
X_3205_ net133 net122 VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__and2_1
X_3136_ net129 net119 VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__and2_1
X_3067_ net395 net73 net27 VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__mux2_1
X_2018_ net500 net175 _0823_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__a21o_1
XFILLER_23_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold161 matmult_inst.mem_inst.matrixB1\[0\] VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 matmult_inst.mem_inst.mem2\[9\] VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _0134_ VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 matmult_inst.alu_inst.out\[10\] VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 matmult_inst.mem_inst.mem2\[14\] VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2705_ net219 net217 net201 net203 VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__and4_1
X_2636_ _1379_ _1381_ VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_7_hz100 clknet_2_3__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_7_hz100
+ sky130_fd_sc_hd__clkbuf_8
X_2567_ _1307_ _1311_ net157 VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__nor3_1
X_2498_ _1245_ _1246_ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__or2_1
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3119_ matmult_inst.fsm_inst.state\[2\] _0762_ net151 _0758_ VGND VGND VPWR VPWR
+ _1601_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_81_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap7 _1560_ VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3470_ clknet_leaf_25_hz100 _0330_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem0\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2421_ _1172_ _1173_ VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__nor2_1
X_2352_ matmult_inst.fsm_inst.tx_start_send net198 _0555_ _1140_ VGND VGND VPWR VPWR
+ _1141_ sky130_fd_sc_hd__a31o_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2283_ _1044_ _1051_ _1053_ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__o21a_1
XFILLER_20_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1998_ net521 net78 net56 VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__mux2_1
X_3668_ clknet_leaf_27_hz100 _0528_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.state\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_2619_ _1313_ _1363_ _1364_ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__o21a_1
X_3599_ clknet_leaf_7_hz100 _0459_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA3\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout290 net291 VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__clkbuf_4
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2970_ net563 net75 net37 VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__mux2_1
X_1921_ matmult_inst.fsm_inst.rx_ready_edge_delay matmult_inst.fsm_inst.rx_ready_edge
+ net154 net165 VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__and4b_1
XFILLER_42_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1852_ net267 net260 matmult_inst.mem_inst.matrixB3\[2\] VGND VGND VPWR VPWR _0725_
+ sky130_fd_sc_hd__and3_1
X_1783_ matmult_inst.mem_inst.matrixA0\[8\] net169 _0661_ net196 _0565_ VGND VGND
+ VPWR VPWR _0662_ sky130_fd_sc_hd__a221o_1
X_3522_ clknet_leaf_17_hz100 _0382_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem3\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3453_ clknet_leaf_29_hz100 _0313_ VGND VGND VPWR VPWR matmult_inst.alu_inst.a0_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_2404_ _1154_ net547 _1165_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__mux2_1
X_3384_ clknet_leaf_29_hz100 _0246_ VGND VGND VPWR VPWR matmult_inst.alu_inst.col0\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2335_ _1123_ _1126_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_10_hz100 clknet_2_3__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_10_hz100
+ sky130_fd_sc_hd__clkbuf_8
X_2266_ _1059_ _1060_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__nor2_1
X_2197_ _0991_ _0992_ _0994_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_25_hz100 clknet_2_2__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_25_hz100
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold32 matmult_inst.mem_inst.matrixA3\[6\] VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 matmult_inst.mem_inst.mem3\[17\] VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 matmult_inst.mem_inst.mem3\[7\] VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 matmult_inst.mem_inst.matrixA3\[1\] VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold54 matmult_inst.mem_inst.matrixB3\[13\] VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 matmult_inst.mem_inst.mem3\[5\] VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold76 matmult_inst.mem_inst.mem2\[10\] VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 _0126_ VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 _0132_ VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2120_ _0867_ net54 _0885_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__o21bai_1
X_2051_ net244 net250 VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_17_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2953_ net488 net73 net39 VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__mux2_1
XFILLER_62_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1904_ matmult_inst.fsm_inst.rx_ready_edge_delay _0771_ _0772_ net154 VGND VGND VPWR
+ VPWR _0773_ sky130_fd_sc_hd__o211a_1
X_2884_ _1136_ _1568_ _1570_ VGND VGND VPWR VPWR _1571_ sky130_fd_sc_hd__or3b_2
XFILLER_30_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1835_ net195 _0704_ _0708_ net288 VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__a22o_1
X_1766_ net269 net262 matmult_inst.mem_inst.mem3\[10\] VGND VGND VPWR VPWR _0647_
+ sky130_fd_sc_hd__and3_1
X_3505_ clknet_leaf_24_hz100 _0365_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem2\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1697_ matmult_inst.mem_inst.matrixA2\[16\] net191 net183 matmult_inst.mem_inst.matrixA1\[16\]
+ _0583_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__a221o_1
X_3436_ clknet_leaf_1_hz100 _0296_ VGND VGND VPWR VPWR matmult_inst.alu_inst.out\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3367_ clknet_leaf_30_hz100 _0231_ VGND VGND VPWR VPWR matmult_inst.alu_inst.row0\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_2318_ _1109_ _1111_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__nand2_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3298_ clknet_leaf_17_hz100 _0168_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB3\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_68_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2249_ _1012_ _1014_ _1013_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__a21bo_1
XFILLER_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1620_ matmult_inst.fsm_inst.state\[1\] matmult_inst.fsm_inst.state\[0\] VGND VGND
+ VPWR VPWR _0539_ sky130_fd_sc_hd__nand2_1
X_3221_ clknet_leaf_11_hz100 _0122_ _0023_ VGND VGND VPWR VPWR matmult_inst.spi_inst.rx_done_sys
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3152_ net136 net116 VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__and2_1
X_2103_ net238 net253 net251 net236 VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__and4_1
X_3083_ net516 net76 net25 VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__mux2_1
XFILLER_54_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2034_ net238 net257 net255 net240 VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__a22o_1
XFILLER_10_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2936_ net356 net71 net42 VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2867_ net222 net426 net93 VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__mux2_1
XFILLER_30_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1818_ matmult_inst.mem_inst.matrixB2\[5\] net189 net181 matmult_inst.mem_inst.matrixB1\[5\]
+ _0693_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__a221o_1
Xhold310 matmult_inst.alu_inst.b0_reg\[0\] VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__dlygate4sd3_1
X_2798_ _1504_ _1512_ VGND VGND VPWR VPWR _1513_ sky130_fd_sc_hd__or2_1
X_1749_ net278 matmult_inst.mem_inst.mem0\[11\] matmult_inst.mem_inst.matrixB0\[11\]
+ net283 VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__a22o_1
Xhold321 matmult_inst.alu_inst.adder_inst.r3.fa0.a VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 matmult_inst.spi_inst.tx_reg_sys\[1\] VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 matmult_inst.spi_inst.tx_reg_sys\[14\] VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 matmult_inst.alu_inst.adder_inst.r1.fa1.a VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__dlygate4sd3_1
X_3419_ clknet_leaf_4_hz100 _0279_ VGND VGND VPWR VPWR matmult_inst.alu_inst.a1_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_28_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2721_ _1460_ _1461_ _1462_ VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__and3_1
X_2652_ _1389_ _1393_ _1394_ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__nand3_1
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2583_ _1234_ _1273_ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__nand2b_1
Xfanout119 net121 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_2
X_3204_ net289 VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__inv_2
X_3135_ net134 net124 VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__and2_1
XFILLER_27_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3066_ net548 net74 net27 VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__mux2_1
X_2017_ net259 net244 net162 VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__and3_1
X_2919_ net277 net178 net88 VGND VGND VPWR VPWR _1584_ sky130_fd_sc_hd__and3_1
XFILLER_50_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold151 matmult_inst.mem_inst.matrixA2\[13\] VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 matmult_inst.alu_inst.row1\[1\] VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 matmult_inst.mem_inst.mem0\[17\] VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 matmult_inst.mem_inst.mem2\[1\] VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 matmult_inst.alu_inst.col0\[3\] VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _0133_ VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2704_ net219 net201 _1446_ VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__a21boi_1
X_2635_ _1339_ _1380_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__nand2_1
X_2566_ _1311_ _1312_ _1307_ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__o21a_1
X_2497_ net207 net224 net209 net223 VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__and4_1
X_3118_ net199 _1599_ _1600_ _1595_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__a22o_1
X_3049_ net423 net72 net29 VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2420_ net228 net211 _1170_ _1171_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__o2bb2a_1
X_2351_ _1139_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__inv_2
X_2282_ _1075_ _1076_ VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__and2b_1
XFILLER_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1997_ matmult_inst.fsm_inst.alu_result\[9\] net114 VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__and2_1
XFILLER_20_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3667_ clknet_leaf_27_hz100 net94 VGND VGND VPWR VPWR matmult_inst.alu_inst.state\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2618_ _1317_ _1318_ _1316_ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__a21boi_1
X_3598_ clknet_leaf_9_hz100 _0458_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA3\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2549_ _1279_ _1280_ net61 VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__nand3_1
XFILLER_28_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout291 net3 VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__clkbuf_2
Xfanout280 net281 VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_6_hz100 clknet_2_1__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_6_hz100
+ sky130_fd_sc_hd__clkbuf_8
X_1920_ net197 net166 net176 _0788_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__a31o_1
X_1851_ net277 matmult_inst.mem_inst.mem0\[2\] matmult_inst.mem_inst.matrixB0\[2\]
+ net282 VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__a22o_1
X_3521_ clknet_leaf_13_hz100 _0381_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem2\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_1782_ net280 matmult_inst.mem_inst.mem0\[8\] matmult_inst.mem_inst.matrixB0\[8\]
+ net285 VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__a22o_1
X_3452_ clknet_leaf_29_hz100 _0312_ VGND VGND VPWR VPWR matmult_inst.alu_inst.a0_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3383_ clknet_leaf_29_hz100 _0245_ VGND VGND VPWR VPWR matmult_inst.alu_inst.col0\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_2403_ _1153_ net448 net63 VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__mux2_1
X_2334_ _1109_ _1124_ _1126_ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_4_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2265_ _1059_ _1060_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__nand2_1
X_2196_ _0937_ _0993_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__nand2b_1
XFILLER_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold22 matmult_inst.mem_inst.matrixB3\[10\] VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 matmult_inst.alu_inst.out\[1\] VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 matmult_inst.mem_inst.matrixA3\[11\] VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 matmult_inst.mem_inst.matrixA3\[3\] VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 matmult_inst.mem_inst.matrixA3\[16\] VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold77 matmult_inst.mem_inst.mem3\[1\] VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 matmult_inst.mem_inst.matrixB0\[16\] VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 matmult_inst.mem_inst.matrixA0\[17\] VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 matmult_inst.mem_inst.mem3\[4\] VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2050_ _0838_ _0849_ _0850_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_17_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2952_ net545 net74 net39 VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__mux2_1
X_1903_ matmult_inst.fsm_inst.rx_ready_edge_delay matmult_inst.fsm_inst.rx_ready_edge
+ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__nand2b_1
XFILLER_30_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2883_ _0552_ net153 _1569_ net197 VGND VGND VPWR VPWR _1570_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_60_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1834_ net281 _0703_ _0706_ net285 VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__a22o_1
X_1765_ matmult_inst.mem_inst.matrixA3\[10\] _0535_ _0645_ VGND VGND VPWR VPWR _0646_
+ sky130_fd_sc_hd__a21o_1
X_3504_ clknet_leaf_16_hz100 _0364_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem2\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1696_ net272 net264 matmult_inst.mem_inst.matrixA3\[16\] VGND VGND VPWR VPWR _0583_
+ sky130_fd_sc_hd__and3_1
X_3435_ clknet_leaf_7_hz100 _0295_ VGND VGND VPWR VPWR matmult_inst.alu_inst.out\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3366_ clknet_leaf_30_hz100 _0230_ VGND VGND VPWR VPWR matmult_inst.alu_inst.row0\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3297_ clknet_leaf_17_hz100 _0167_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB3\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2317_ _1110_ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__inv_2
X_2248_ net250 net233 VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_68_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2179_ net253 net251 net232 net234 VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__nand4_1
XFILLER_25_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_24_hz100 clknet_2_2__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_24_hz100
+ sky130_fd_sc_hd__clkbuf_8
X_3220_ net290 VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__inv_2
X_3151_ net131 net120 VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__and2_1
XFILLER_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2102_ net238 net252 net236 net253 VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__a22oi_1
X_3082_ net480 _0814_ net25 VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__mux2_1
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2033_ _0834_ _0835_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__nor2_1
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2935_ net369 net72 net41 VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__mux2_1
X_2866_ net225 net588 net93 VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1817_ net271 net263 matmult_inst.mem_inst.matrixB3\[5\] VGND VGND VPWR VPWR _0693_
+ sky130_fd_sc_hd__and3_1
X_2797_ _1492_ _1497_ _1500_ _1503_ _1498_ VGND VGND VPWR VPWR _1512_ sky130_fd_sc_hd__o311a_1
Xhold311 matmult_inst.alu_inst.adder_inst.r1.fa0.b VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold300 matmult_inst.mem_inst.matrixB1\[9\] VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold333 matmult_inst.alu_inst.adder_inst.r3.fa3.b VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold322 matmult_inst.alu_inst.adder_inst.r1.fa3.b VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__dlygate4sd3_1
X_1748_ net630 net91 _0630_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__o21a_1
Xhold344 matmult_inst.spi_inst.tx_reg_sys\[10\] VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__dlygate4sd3_1
X_1679_ net282 net277 VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__nor2_1
Xhold355 matmult_inst.alu_inst.adder_inst.r0.fa3.b VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__dlygate4sd3_1
X_3418_ clknet_leaf_2_hz100 _0278_ VGND VGND VPWR VPWR matmult_inst.alu_inst.a1_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3349_ clknet_leaf_3_hz100 _0214_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r2.fa0.b
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2720_ _1412_ _1448_ _1447_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__o21ba_1
X_2651_ _1389_ _1393_ _1394_ VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__and3_1
XFILLER_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2582_ _1270_ _1326_ net105 VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__nand3_1
XFILLER_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3203_ net289 VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__inv_2
XFILLER_79_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3134_ net132 net120 VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__and2_1
X_3065_ net418 net75 net27 VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__mux2_1
X_2016_ net174 VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__inv_2
XFILLER_23_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2918_ net434 net70 net44 VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__mux2_1
XFILLER_12_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2849_ _1554_ _1555_ VGND VGND VPWR VPWR _1556_ sky130_fd_sc_hd__xnor2_1
Xhold152 matmult_inst.mem_inst.mem1\[1\] VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 matmult_inst.alu_inst.out\[2\] VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 matmult_inst.mem_inst.matrixA1\[16\] VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 matmult_inst.spi_inst.mosi_data_sync\[0\] VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 matmult_inst.mem_inst.matrixA2\[12\] VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 matmult_inst.mem_inst.matrixB0\[9\] VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 matmult_inst.mem_inst.matrixA0\[8\] VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2703_ net218 net203 VGND VGND VPWR VPWR _1446_ sky130_fd_sc_hd__nand2_1
X_2634_ _1302_ _1303_ _1304_ _1340_ VGND VGND VPWR VPWR _1380_ sky130_fd_sc_hd__a211o_1
X_2565_ _1308_ _1309_ _1310_ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__a21oi_1
X_2496_ net207 net224 net209 net223 VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__a22oi_1
X_3117_ net199 _0766_ _0554_ VGND VGND VPWR VPWR _1600_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_27_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3048_ net341 net73 net29 VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_45_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout91 net92 VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_4
Xfanout80 _0811_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_2
XFILLER_80_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2350_ _0769_ _1136_ _1138_ _0781_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__and4bb_1
X_2281_ _1041_ _1074_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_63_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_72_Left_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1996_ net319 net79 net56 VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__mux2_1
X_3666_ clknet_leaf_27_hz100 net161 VGND VGND VPWR VPWR matmult_inst.alu_inst.state\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2617_ _1307_ _1311_ net157 _1319_ _1320_ VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__o32a_1
X_3597_ clknet_leaf_25_hz100 _0457_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA3\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_81_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2548_ _1289_ _1295_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__xor2_1
X_2479_ _1227_ _1228_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__or2_1
XFILLER_75_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload0 clknet_2_0__leaf_hz100 VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__inv_8
XFILLER_50_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout270 matmult_inst.addr\[0\] VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__clkbuf_2
Xfanout281 matmult_inst.fsm_inst.sel\[2\] VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__buf_2
Xfanout292 net293 VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__buf_2
XFILLER_75_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1850_ matmult_inst.mem_inst.mem2\[2\] net186 net178 matmult_inst.mem_inst.mem1\[2\]
+ _0722_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__a221o_1
X_1781_ net639 net91 _0652_ _0660_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_12_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3520_ clknet_leaf_19_hz100 _0380_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem2\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_3451_ clknet_leaf_29_hz100 _0311_ VGND VGND VPWR VPWR matmult_inst.alu_inst.a0_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2402_ _0766_ _1164_ _1162_ VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__o21ai_2
X_3382_ clknet_leaf_28_hz100 _0244_ VGND VGND VPWR VPWR matmult_inst.alu_inst.col0\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2333_ _1100_ _1122_ _1121_ VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_4_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2264_ _1022_ _1024_ _1021_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__a21bo_1
X_2195_ _0933_ _0934_ _0936_ net68 VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__a31o_1
XFILLER_80_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1979_ matmult_inst.fsm_inst.rx_data\[0\] _0786_ net113 matmult_inst.fsm_inst.alu_result\[0\]
+ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__a22o_1
XFILLER_20_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3649_ clknet_leaf_17_hz100 _0509_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB2\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold12 _0124_ VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 matmult_inst.mem_inst.matrixA3\[4\] VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 matmult_inst.mem_inst.mem3\[11\] VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 matmult_inst.mem_inst.matrixA3\[0\] VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold34 matmult_inst.mem_inst.matrixA3\[5\] VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 matmult_inst.mem_inst.matrixB2\[11\] VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 matmult_inst.mem_inst.mem3\[6\] VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 matmult_inst.mem_inst.matrixA2\[4\] VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2951_ net549 net75 net39 VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__mux2_1
XFILLER_15_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1902_ matmult_inst.fsm_inst.count\[2\] _1605_ _0770_ VGND VGND VPWR VPWR _0771_
+ sky130_fd_sc_hd__or3b_2
X_2882_ matmult_inst.fsm_inst.count\[2\] _1605_ net177 _0766_ VGND VGND VPWR VPWR
+ _1569_ sky130_fd_sc_hd__a31o_1
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1833_ matmult_inst.mem_inst.matrixA2\[4\] net190 net182 matmult_inst.mem_inst.matrixA1\[4\]
+ _0707_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__a221o_1
X_1764_ matmult_inst.mem_inst.matrixA2\[10\] net188 net180 matmult_inst.mem_inst.matrixA1\[10\]
+ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__a22o_1
X_3503_ clknet_leaf_13_hz100 _0363_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem1\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_1695_ matmult_inst.mem_inst.matrixA0\[16\] net169 _0581_ net196 net115 VGND VGND
+ VPWR VPWR _0582_ sky130_fd_sc_hd__a221o_1
X_3434_ clknet_leaf_7_hz100 _0294_ VGND VGND VPWR VPWR matmult_inst.alu_inst.out\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3365_ clknet_leaf_29_hz100 _0229_ VGND VGND VPWR VPWR matmult_inst.alu_inst.row0\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_2316_ _1080_ _1094_ _1108_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__and3_1
X_3296_ clknet_leaf_9_hz100 net583 _0077_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.rx_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2247_ _1008_ _1016_ _1010_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_68_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2178_ net253 net232 net234 net251 VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_51_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_5_hz100 clknet_2_1__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_5_hz100
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3150_ net129 net119 VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__and2_1
XFILLER_39_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3081_ net594 _0813_ net26 VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__mux2_1
X_2101_ _0891_ _0898_ _0899_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__and3_1
X_2032_ net243 net254 net244 net252 VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2934_ net555 _0818_ net41 VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__mux2_1
X_2865_ net226 net554 net94 VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__mux2_1
XFILLER_30_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1816_ matmult_inst.mem_inst.mem2\[5\] net190 net182 matmult_inst.mem_inst.mem1\[5\]
+ _0691_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__a221o_1
Xhold301 matmult_inst.alu_inst.col0\[2\] VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2796_ _1509_ _1510_ VGND VGND VPWR VPWR _1511_ sky130_fd_sc_hd__and2b_1
Xhold323 matmult_inst.spi_inst.tx_reg_sys\[8\] VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__dlygate4sd3_1
X_1747_ net283 _0624_ _0629_ _0622_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__a211o_1
Xhold312 matmult_inst.mem_inst.matrixA2\[14\] VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 matmult_inst.spi_inst.tx_reg_sys\[16\] VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__dlygate4sd3_1
X_1678_ net272 net264 VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__nor2_1
Xhold356 matmult_inst.alu_inst.adder_inst.r0.fa1.b VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 matmult_inst.spi_inst.tx_reg_sys\[9\] VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__dlygate4sd3_1
X_3417_ clknet_leaf_4_hz100 _0277_ VGND VGND VPWR VPWR matmult_inst.alu_inst.a1_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3348_ clknet_leaf_2_hz100 _0213_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r1.fa3.b
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3279_ net292 _0021_ _0060_ VGND VGND VPWR VPWR matmult_inst.spi_inst.miso_shifter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2650_ _1393_ _1394_ _1389_ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2581_ _1326_ _1327_ _1270_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__a21o_1
X_3202_ net289 VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_78_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3133_ net132 net120 VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__and2_1
X_3064_ net439 net76 net27 VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__mux2_1
X_2015_ matmult_inst.alu_inst.state\[1\] matmult_inst.alu_inst.state\[0\] VGND VGND
+ VPWR VPWR _0822_ sky130_fd_sc_hd__nand2b_1
XFILLER_50_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2917_ net362 net71 net44 VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__mux2_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2848_ _1547_ _1550_ _1548_ VGND VGND VPWR VPWR _1555_ sky130_fd_sc_hd__o21ai_1
X_2779_ net380 _1496_ net163 VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__mux2_1
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold120 matmult_inst.mem_inst.matrixA0\[15\] VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 matmult_inst.mem_inst.matrixA1\[3\] VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 _0125_ VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 matmult_inst.mem_inst.mem1\[17\] VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 _0159_ VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 matmult_inst.mem_inst.matrixB1\[10\] VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 matmult_inst.mem_inst.matrixB2\[17\] VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 matmult_inst.mem_inst.matrixA1\[5\] VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_hz100 clknet_2_2__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_23_hz100
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2702_ _1443_ _1444_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_30_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2633_ _1376_ _1378_ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__nand2_1
X_2564_ _1308_ _1309_ _1310_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__and3_1
X_2495_ _1239_ _1240_ _1242_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__and3_1
X_3116_ _1597_ _1599_ net200 VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3047_ net420 net74 net29 VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout92 matmult_inst.fsm_inst.load VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_4
Xfanout81 _0810_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_2
Xfanout70 _0821_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_2
XFILLER_80_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2280_ _1041_ _1074_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__and2_1
XFILLER_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1995_ matmult_inst.fsm_inst.alu_result\[8\] net113 VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__and2_1
XFILLER_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3665_ clknet_leaf_14_hz100 _0525_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB2\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_2616_ _1270_ net104 VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__nand2_1
X_3596_ clknet_leaf_23_hz100 _0456_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA3\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2547_ _1293_ _1294_ VGND VGND VPWR VPWR _1295_ sky130_fd_sc_hd__or2_1
X_2478_ _1211_ net51 VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__and2_1
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload1 clknet_2_1__leaf_hz100 VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__inv_6
Xwire149 _0857_ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout260 net262 VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__buf_2
Xfanout282 net284 VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__buf_2
Xfanout271 net274 VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__buf_2
Xfanout293 net3 VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_57_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1780_ net288 _0654_ _0659_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_12_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3450_ clknet_leaf_29_hz100 _0310_ VGND VGND VPWR VPWR matmult_inst.alu_inst.a0_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2401_ matmult_inst.fsm_inst.count\[1\] _1604_ _0544_ VGND VGND VPWR VPWR _1164_
+ sky130_fd_sc_hd__a21oi_1
X_3381_ clknet_leaf_28_hz100 _0243_ VGND VGND VPWR VPWR matmult_inst.alu_inst.col0\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2332_ _1109_ _1124_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__nand2_1
XFILLER_69_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2263_ net52 VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__inv_2
X_2194_ _0973_ _0974_ net67 VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__a21o_1
XFILLER_80_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1978_ net282 net198 net88 VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__and3_1
X_3648_ clknet_leaf_17_hz100 _0508_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB2\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3579_ clknet_leaf_25_hz100 _0439_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA2\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold13 matmult_inst.mem_inst.matrixA3\[17\] VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 matmult_inst.mem_inst.matrixB3\[12\] VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 matmult_inst.mem_inst.mem3\[9\] VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 matmult_inst.mem_inst.matrixB3\[4\] VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold57 matmult_inst.mem_inst.matrixB3\[11\] VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 matmult_inst.mem_inst.mem0\[16\] VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 matmult_inst.mem_inst.matrixB2\[16\] VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2950_ net417 net76 net39 VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__mux2_1
X_2881_ _0541_ _1567_ VGND VGND VPWR VPWR _1568_ sky130_fd_sc_hd__nor2_1
X_1901_ matmult_inst.fsm_inst.count\[1\] matmult_inst.fsm_inst.count\[0\] VGND VGND
+ VPWR VPWR _0770_ sky130_fd_sc_hd__nor2_1
X_1832_ net271 net263 matmult_inst.mem_inst.matrixA3\[4\] VGND VGND VPWR VPWR _0707_
+ sky130_fd_sc_hd__and3_1
X_1763_ matmult_inst.mem_inst.matrixB2\[10\] net188 net180 matmult_inst.mem_inst.matrixB1\[10\]
+ _0643_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__a221o_1
X_3502_ clknet_leaf_15_hz100 _0362_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem1\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_1694_ net280 matmult_inst.mem_inst.mem0\[16\] matmult_inst.mem_inst.matrixB0\[16\]
+ net286 VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__a22o_1
X_3433_ clknet_leaf_1_hz100 _0293_ VGND VGND VPWR VPWR matmult_inst.alu_inst.out\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3364_ clknet_leaf_28_hz100 _0228_ VGND VGND VPWR VPWR matmult_inst.alu_inst.row0\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2315_ _1080_ _1094_ _1108_ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__a21o_1
X_3295_ clknet_leaf_9_hz100 net336 _0076_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.rx_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2246_ _1039_ _1041_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_68_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2177_ _0941_ _0942_ _0940_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__o21bai_1
XFILLER_53_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3080_ net378 _0812_ net26 VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__mux2_1
X_2100_ _0898_ _0899_ _0891_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__a21oi_1
X_2031_ net243 net254 net244 net252 VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_65_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2933_ net608 net74 net41 VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2864_ net228 net576 net94 VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__mux2_1
XFILLER_30_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2795_ matmult_inst.alu_inst.adder_inst.r1.fa2.b matmult_inst.alu_inst.adder_inst.r1.fa2.a
+ VGND VGND VPWR VPWR _1510_ sky130_fd_sc_hd__nand2_1
X_1815_ net274 net266 matmult_inst.mem_inst.mem3\[5\] VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__and3_1
X_1746_ net287 _0626_ _0628_ net278 VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__a22o_1
Xhold302 matmult_inst.mem_inst.mem0\[1\] VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold313 matmult_inst.alu_inst.adder_inst.r3.fa2.a VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 matmult_inst.spi_inst.tx_reg_sys\[11\] VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 matmult_inst.spi_inst.tx_reg_sys\[7\] VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__dlygate4sd3_1
X_1677_ net115 VGND VGND VPWR VPWR matmult_inst.fsm_inst.load sky130_fd_sc_hd__inv_2
Xhold357 matmult_inst.alu_inst.adder_inst.r0.fa1.a VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 matmult_inst.alu_inst.adder_inst.r1.fa0.a VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__dlygate4sd3_1
X_3416_ clknet_leaf_6_hz100 _0276_ VGND VGND VPWR VPWR matmult_inst.alu_inst.a1_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3347_ clknet_leaf_2_hz100 _0212_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r1.fa2.b
+ sky130_fd_sc_hd__dfxtp_1
X_3278_ net292 _0020_ _0059_ VGND VGND VPWR VPWR matmult_inst.spi_inst.miso_shifter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2229_ _1021_ _1022_ _1024_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__a21o_1
XFILLER_53_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2580_ net139 _1293_ _1294_ net138 _1288_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__o311ai_2
X_3201_ net289 VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__inv_2
XFILLER_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3132_ net129 net118 VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_78_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3063_ net404 net77 net27 VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__mux2_1
X_2014_ net322 net70 net56 VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_4_hz100 clknet_2_1__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_4_hz100
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_23_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2916_ net409 net72 net43 VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__mux2_1
X_2847_ _1552_ _1553_ VGND VGND VPWR VPWR _1554_ sky130_fd_sc_hd__nand2_1
Xhold110 matmult_inst.mem_inst.matrixB0\[10\] VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__dlygate4sd3_1
X_2778_ _1494_ _1495_ VGND VGND VPWR VPWR _1496_ sky130_fd_sc_hd__xnor2_1
Xhold132 matmult_inst.alu_inst.row0\[3\] VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 matmult_inst.alu_inst.col0\[5\] VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__dlygate4sd3_1
X_1729_ net269 net262 matmult_inst.mem_inst.matrixA3\[13\] VGND VGND VPWR VPWR _0613_
+ sky130_fd_sc_hd__and3_1
Xhold121 matmult_inst.mem_inst.matrixB3\[1\] VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 matmult_inst.mem_inst.mem0\[11\] VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 matmult_inst.mem_inst.matrixB1\[3\] VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 matmult_inst.alu_inst.col1\[0\] VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 matmult_inst.mem_inst.matrixA1\[15\] VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 matmult_inst.mem_inst.mem0\[13\] VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2701_ _1441_ _1442_ VGND VGND VPWR VPWR _1444_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_30_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2632_ net14 VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__inv_2
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2563_ net207 net221 VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__nand2_1
X_2494_ _1239_ _1240_ _1242_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__a21oi_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3115_ _1595_ _1598_ VGND VGND VPWR VPWR _1599_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_38_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3046_ net376 net75 net29 VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__mux2_1
XFILLER_63_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout71 _0820_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_2
Xfanout82 _0809_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_2
Xfanout93 net94 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1994_ net353 net80 net56 VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__mux2_1
XFILLER_20_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3664_ clknet_leaf_14_hz100 _0524_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB2\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_2615_ _1355_ net137 VGND VGND VPWR VPWR _1361_ sky130_fd_sc_hd__xnor2_1
X_3595_ clknet_leaf_24_hz100 _0455_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA3\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_22_hz100 clknet_2_2__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_22_hz100
+ sky130_fd_sc_hd__clkbuf_8
X_2546_ _1290_ _1291_ _1292_ VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__and3_1
X_2477_ _1211_ _1226_ VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__nor2_1
XFILLER_18_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3029_ net606 net73 net31 VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__mux2_1
XFILLER_34_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload2 clknet_2_2__leaf_hz100 VGND VGND VPWR VPWR clkload2/X sky130_fd_sc_hd__clkbuf_8
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout250 matmult_inst.alu_inst.a1_reg\[4\] VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkbuf_4
Xfanout261 net262 VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__clkbuf_2
Xfanout283 net284 VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__clkbuf_4
Xfanout272 net274 VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__clkbuf_2
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2400_ _1160_ net533 net65 VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__mux2_1
X_3380_ clknet_leaf_27_hz100 _0242_ VGND VGND VPWR VPWR matmult_inst.alu_inst.col0\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2331_ _1066_ _1089_ _1091_ _1110_ _1088_ VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__a311o_1
X_2262_ _1043_ _1056_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__xor2_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2193_ _0973_ _0974_ net67 VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__nand3_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1977_ _0786_ net114 VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__or2_1
X_3647_ clknet_leaf_13_hz100 _0507_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB1\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_3578_ clknet_leaf_23_hz100 _0438_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA2\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2529_ _1212_ _1238_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__nand2_1
Xhold14 matmult_inst.alu_inst.out\[16\] VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold47 matmult_inst.mem_inst.matrixA3\[14\] VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 matmult_inst.mem_inst.matrixB3\[5\] VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 matmult_inst.mem_inst.matrixB3\[8\] VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 matmult_inst.mem_inst.matrixB3\[3\] VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 matmult_inst.mem_inst.matrixB1\[16\] VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2880_ matmult_inst.fsm_inst.tx_ready _0564_ _0798_ matmult_inst.fsm_inst.load_delay
+ VGND VGND VPWR VPWR _1567_ sky130_fd_sc_hd__o22a_1
X_1900_ _0537_ _0549_ _0768_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_25_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1831_ matmult_inst.mem_inst.matrixB2\[4\] net190 net182 matmult_inst.mem_inst.matrixB1\[4\]
+ _0705_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__a221o_1
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1762_ net268 net261 matmult_inst.mem_inst.matrixB3\[10\] VGND VGND VPWR VPWR _0643_
+ sky130_fd_sc_hd__and3_1
X_3501_ clknet_leaf_22_hz100 _0361_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem1\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_1693_ net622 net91 _0580_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__o21a_1
X_3432_ clknet_leaf_26_hz100 _0292_ VGND VGND VPWR VPWR matmult_inst.alu_inst.out\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3363_ clknet_leaf_28_hz100 _0227_ VGND VGND VPWR VPWR matmult_inst.alu_inst.row0\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2314_ _1101_ net111 VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__xnor2_1
X_3294_ clknet_leaf_5_hz100 net572 _0075_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.rx_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2245_ net251 net231 _1040_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__and3_1
XFILLER_38_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2176_ _0970_ _0971_ _0972_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_68_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_69_Left_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2030_ _0832_ _0833_ net510 net175 VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_65_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap90 _0768_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
X_2932_ net406 net75 net41 VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2863_ net602 _0796_ _1565_ _1566_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__a22o_1
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2794_ matmult_inst.alu_inst.adder_inst.r1.fa2.b matmult_inst.alu_inst.adder_inst.r1.fa2.a
+ VGND VGND VPWR VPWR _1509_ sky130_fd_sc_hd__nor2_1
X_1814_ net620 _0690_ net91 VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__mux2_1
X_1745_ matmult_inst.mem_inst.mem3\[12\] net198 _0627_ VGND VGND VPWR VPWR _0628_
+ sky130_fd_sc_hd__a21o_1
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold314 matmult_inst.mem_inst.mem1\[13\] VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 matmult_inst.alu_inst.adder_inst.r2.fa2.b VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold303 matmult_inst.mem_inst.matrixB1\[7\] VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 matmult_inst.fsm_inst.count\[3\] VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__dlygate4sd3_1
X_1676_ matmult_inst.spi_inst.current_state _0541_ _0564_ VGND VGND VPWR VPWR _0565_
+ sky130_fd_sc_hd__or3_2
Xhold347 matmult_inst.alu_inst.adder_inst.r1.fa2.a VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 matmult_inst.spi_inst.tx_reg_sys\[12\] VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__dlygate4sd3_1
X_3415_ clknet_leaf_6_hz100 _0275_ VGND VGND VPWR VPWR matmult_inst.alu_inst.a1_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3346_ clknet_leaf_6_hz100 _0211_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r1.fa1.b
+ sky130_fd_sc_hd__dfxtp_1
X_3277_ net292 _0019_ _0058_ VGND VGND VPWR VPWR matmult_inst.spi_inst.miso_shifter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2228_ _1021_ _1022_ _1024_ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__nand3_1
XFILLER_38_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2159_ _0937_ _0938_ net68 VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_36_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3200_ net289 VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__inv_2
X_3131_ net130 net118 VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_78_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3062_ net457 net78 net28 VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__mux2_1
X_2013_ matmult_inst.fsm_inst.alu_result\[17\] net113 VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__and2_1
XFILLER_35_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2915_ net558 net73 net43 VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__mux2_1
X_2846_ matmult_inst.alu_inst.adder_inst.r3.fa2.b matmult_inst.alu_inst.adder_inst.r3.fa2.a
+ VGND VGND VPWR VPWR _1553_ sky130_fd_sc_hd__nand2_1
X_2777_ _1486_ _1490_ _1487_ VGND VGND VPWR VPWR _1495_ sky130_fd_sc_hd__o21ai_1
Xhold100 matmult_inst.mem_inst.mem2\[7\] VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold122 matmult_inst.mem_inst.matrixB2\[12\] VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__dlygate4sd3_1
X_1728_ matmult_inst.mem_inst.matrixA0\[13\] net168 _0611_ net195 net115 VGND VGND
+ VPWR VPWR _0612_ sky130_fd_sc_hd__a221o_1
Xhold111 matmult_inst.mem_inst.mem2\[6\] VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 matmult_inst.mem_inst.mem2\[8\] VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 matmult_inst.mem_inst.matrixA0\[4\] VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__dlygate4sd3_1
X_1659_ matmult_inst.cs _0556_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__or2_4
Xhold166 matmult_inst.mem_inst.mem2\[0\] VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 matmult_inst.mem_inst.matrixA1\[7\] VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 matmult_inst.mem_inst.matrixA2\[9\] VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 matmult_inst.mem_inst.mem0\[12\] VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 matmult_inst.alu_inst.row1\[4\] VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3329_ _0104_ _0197_ _0103_ VGND VGND VPWR VPWR matmult_inst.spi_inst.mosi_data_spi\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2700_ _1441_ _1442_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__and2_1
X_2631_ _1373_ _1374_ _1336_ VGND VGND VPWR VPWR _1377_ sky130_fd_sc_hd__a21oi_1
X_2562_ net205 net224 net222 net203 VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__nand4_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2493_ _1214_ _1215_ _1241_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__o21a_1
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3114_ matmult_inst.fsm_inst.state\[1\] matmult_inst.fsm_inst.state\[0\] net199 matmult_inst.fsm_inst.state\[4\]
+ VGND VGND VPWR VPWR _1598_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_38_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3045_ net349 net76 net29 VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__mux2_1
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2829_ _1537_ _1538_ VGND VGND VPWR VPWR _1539_ sky130_fd_sc_hd__nand2_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout72 _0819_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_2
Xfanout83 _0808_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
XFILLER_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout94 _0527_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_2
XFILLER_10_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_3_hz100 clknet_2_1__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_3_hz100
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_32_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1993_ matmult_inst.fsm_inst.rx_data\[7\] _0786_ net113 matmult_inst.fsm_inst.alu_result\[7\]
+ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__a22o_1
XFILLER_20_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3663_ clknet_leaf_21_hz100 _0523_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB2\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload20 clknet_leaf_25_hz100 VGND VGND VPWR VPWR clkload20/Y sky130_fd_sc_hd__clkinv_2
XPHY_EDGE_ROW_41_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2614_ _1356_ _1359_ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__xnor2_1
X_3594_ clknet_leaf_17_hz100 _0454_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA3\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2545_ _1290_ _1291_ _1292_ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__a21oi_1
X_2476_ _1219_ net107 VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__xnor2_1
XFILLER_28_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_50_Left_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3028_ net445 net74 net31 VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__mux2_1
XFILLER_34_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload3 clknet_leaf_27_hz100 VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__clkinv_8
XFILLER_50_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout240 matmult_inst.alu_inst.b1_reg\[2\] VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__buf_2
Xfanout262 matmult_inst.addr\[1\] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__buf_2
Xfanout273 net274 VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout251 matmult_inst.alu_inst.a1_reg\[3\] VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__buf_2
Xfanout284 matmult_inst.fsm_inst.sel\[1\] VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__clkbuf_2
XFILLER_75_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2330_ _1100_ _1121_ _1122_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__and3_1
X_2261_ _1054_ _1055_ _1043_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__a21o_1
X_2192_ _0983_ _0989_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__xnor2_1
XFILLER_65_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1976_ _0547_ _0778_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__nor2_1
XFILLER_20_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3646_ clknet_leaf_14_hz100 _0506_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB1\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_3577_ clknet_leaf_24_hz100 _0437_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA2\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2528_ _1273_ _1274_ _1234_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_3_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold26 matmult_inst.mem_inst.mem3\[14\] VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ _1188_ _1209_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__xnor2_1
Xhold15 _0139_ VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 matmult_inst.mem_inst.matrixA3\[8\] VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 matmult_inst.alu_inst.out\[12\] VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 matmult_inst.mem_inst.matrixB3\[7\] VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_7_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_hz100 clknet_2_2__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_21_hz100
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_30_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1830_ net271 net263 matmult_inst.mem_inst.matrixB3\[4\] VGND VGND VPWR VPWR _0705_
+ sky130_fd_sc_hd__and3_1
X_1761_ matmult_inst.mem_inst.matrixA0\[10\] net168 _0641_ net194 net115 VGND VGND
+ VPWR VPWR _0642_ sky130_fd_sc_hd__a221o_1
X_3500_ clknet_leaf_20_hz100 _0360_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem1\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_1692_ net286 _0574_ _0579_ _0570_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__a211o_1
X_3431_ clknet_leaf_1_hz100 _0291_ VGND VGND VPWR VPWR matmult_inst.alu_inst.out\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3362_ clknet_leaf_27_hz100 _0226_ VGND VGND VPWR VPWR matmult_inst.alu_inst.row0\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2313_ _1069_ _1106_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__xnor2_1
X_3293_ clknet_leaf_6_hz100 net523 _0074_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.rx_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2244_ net253 net232 _1003_ _1005_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__a22o_1
X_2175_ _0970_ _0971_ _0972_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__a21o_1
XFILLER_25_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1959_ net305 net57 net22 matmult_inst.fsm_inst.alu_result\[1\] VGND VGND VPWR VPWR
+ _0124_ sky130_fd_sc_hd__a22o_1
X_3629_ clknet_leaf_15_hz100 _0489_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB0\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2931_ net591 net76 net41 VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2862_ matmult_inst.alu_inst.adder_inst.fa.b matmult_inst.alu_inst.adder_inst.fa.a
+ net163 VGND VGND VPWR VPWR _1566_ sky130_fd_sc_hd__o21a_1
X_1813_ matmult_inst.mem_inst.matrixA0\[6\] net169 _0688_ _0689_ VGND VGND VPWR VPWR
+ _0690_ sky130_fd_sc_hd__a211o_1
X_2793_ net520 _1508_ net164 VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__mux2_1
X_1744_ matmult_inst.mem_inst.mem2\[12\] net188 net180 matmult_inst.mem_inst.mem1\[12\]
+ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__a22o_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold304 matmult_inst.mem_inst.mem1\[2\] VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 matmult_inst.spi_inst.tx_reg_sys\[6\] VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 matmult_inst.mem_inst.matrixB2\[7\] VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__dlygate4sd3_1
X_1675_ matmult_inst.fsm_inst.count\[1\] _1604_ _0544_ VGND VGND VPWR VPWR _0564_
+ sky130_fd_sc_hd__or3_2
Xhold348 matmult_inst.spi_inst.tx_reg_sys\[13\] VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 matmult_inst.alu_inst.adder_inst.r2.fa1.a VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__dlygate4sd3_1
X_3414_ clknet_leaf_2_hz100 _0274_ VGND VGND VPWR VPWR matmult_inst.alu_inst.a1_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold359 matmult_inst.fsm_inst.rx_valid_delay VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3345_ clknet_leaf_2_hz100 _0210_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r1.fa0.b
+ sky130_fd_sc_hd__dfxtp_1
X_3276_ net292 _0018_ _0057_ VGND VGND VPWR VPWR matmult_inst.spi_inst.miso_shifter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2227_ net255 net231 _1023_ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__and3_1
XFILLER_38_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2158_ _0937_ _0938_ net68 VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2089_ _0874_ _0881_ _0849_ _0873_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_36_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3130_ net130 net118 VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_78_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3061_ net557 net79 net28 VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2012_ net303 net71 net56 VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2914_ net481 net74 net43 VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__mux2_1
XFILLER_31_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2845_ matmult_inst.alu_inst.adder_inst.r3.fa2.b matmult_inst.alu_inst.adder_inst.r3.fa2.a
+ VGND VGND VPWR VPWR _1552_ sky130_fd_sc_hd__or2_1
XFILLER_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold101 matmult_inst.mem_inst.matrixB0\[14\] VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__dlygate4sd3_1
X_2776_ _1492_ _1493_ VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__nand2b_1
Xhold112 matmult_inst.mem_inst.mem1\[12\] VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 matmult_inst.mem_inst.mem2\[11\] VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 matmult_inst.mem_inst.matrixA1\[10\] VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__dlygate4sd3_1
X_1727_ net278 matmult_inst.mem_inst.mem0\[13\] matmult_inst.mem_inst.matrixB0\[13\]
+ net283 VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__a22o_1
Xhold145 matmult_inst.mem_inst.matrixB0\[11\] VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 matmult_inst.mem_inst.mem0\[2\] VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 matmult_inst.alu_inst.out\[15\] VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__dlygate4sd3_1
X_1658_ net296 matmult_inst.spi_inst.rx_done_sys VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__or2_1
Xhold178 matmult_inst.mem_inst.matrixB2\[14\] VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 matmult_inst.mem_inst.mem0\[7\] VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__dlygate4sd3_1
X_3328_ _0102_ _0196_ _0101_ VGND VGND VPWR VPWR matmult_inst.spi_inst.mosi_data_spi\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3259_ clknet_leaf_10_hz100 _0148_ _0040_ VGND VGND VPWR VPWR matmult_inst.spi_inst.tx_reg_sys\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2630_ _1336_ _1373_ _1374_ VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__nand3_1
X_2561_ net205 net222 net203 net224 VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__a22o_1
X_2492_ _1214_ _1215_ _1191_ VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__a21o_1
XFILLER_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3113_ net200 _1597_ _0538_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__a21bo_1
XFILLER_67_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3044_ net473 net77 net29 VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2828_ matmult_inst.alu_inst.adder_inst.r2.fa3.b matmult_inst.alu_inst.adder_inst.r2.fa3.a
+ VGND VGND VPWR VPWR _1538_ sky130_fd_sc_hd__nand2_1
X_2759_ matmult_inst.alu_inst.adder_inst.r0.fa0.b matmult_inst.alu_inst.adder_inst.r0.fa0.a
+ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__nand2_1
XFILLER_48_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout40 _1585_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_4
Xfanout73 _0818_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_2
Xfanout84 _0807_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_2
Xfanout95 net97 VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1992_ net313 net81 net56 VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__mux2_1
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3662_ clknet_leaf_19_hz100 _0522_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB2\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload10 clknet_leaf_4_hz100 VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__inv_8
X_2613_ net219 _1358_ _1357_ VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__a21bo_1
Xclkload21 clknet_leaf_7_hz100 VGND VGND VPWR VPWR clkload21/X sky130_fd_sc_hd__clkbuf_4
X_3593_ clknet_leaf_14_hz100 _0453_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA2\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_2544_ net216 net215 VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__nand2_1
X_2475_ _1190_ _1224_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3027_ net479 net75 net31 VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__mux2_1
XFILLER_63_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload4 clknet_leaf_28_hz100 VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__inv_8
XFILLER_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout230 matmult_inst.alu_inst.b1_reg\[7\] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__buf_2
Xfanout241 matmult_inst.alu_inst.b1_reg\[2\] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_2
Xfanout274 matmult_inst.addr\[0\] VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__clkbuf_2
Xfanout263 net266 VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__buf_2
Xfanout252 matmult_inst.alu_inst.a1_reg\[3\] VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__clkbuf_2
Xfanout285 matmult_inst.fsm_inst.sel\[1\] VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__clkbuf_4
XFILLER_46_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2260_ _1054_ _1055_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__nand2_1
XFILLER_37_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2191_ _0987_ _0988_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__nand2_1
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1975_ net602 net57 net22 matmult_inst.fsm_inst.alu_result\[17\] VGND VGND VPWR VPWR
+ _0140_ sky130_fd_sc_hd__a22o_1
X_3645_ clknet_leaf_21_hz100 _0505_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB1\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3576_ clknet_leaf_17_hz100 _0436_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA2\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2527_ _1234_ _1273_ net106 VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__nand3_1
X_2458_ _1207_ _1208_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_3_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold27 matmult_inst.mem_inst.mem3\[10\] VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 matmult_inst.mem_inst.matrixB3\[14\] VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 matmult_inst.mem_inst.matrixA3\[7\] VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 _0135_ VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__dlygate4sd3_1
X_2389_ _1159_ net388 _1161_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__mux2_1
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_2_hz100 clknet_2_1__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_2_hz100
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_51_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1760_ net278 matmult_inst.mem_inst.mem0\[10\] matmult_inst.mem_inst.matrixB0\[10\]
+ net284 VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__a22o_1
X_1691_ net288 _0576_ _0578_ net280 VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__a22o_1
X_3430_ clknet_leaf_1_hz100 _0290_ VGND VGND VPWR VPWR matmult_inst.alu_inst.out\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3361_ clknet_leaf_27_hz100 _0225_ VGND VGND VPWR VPWR matmult_inst.alu_inst.row0\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2312_ _1104_ _1105_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__or2_1
X_3292_ clknet_leaf_5_hz100 net593 _0073_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.rx_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2243_ _1038_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__inv_2
X_2174_ _0912_ _0929_ _0930_ _0932_ _0894_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__a32o_1
XFILLER_65_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1958_ net569 net57 net22 net530 VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__a22o_1
X_1889_ _0551_ _0757_ _0756_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__o21ai_1
X_3628_ clknet_leaf_15_hz100 _0488_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB0\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_3559_ clknet_leaf_24_hz100 _0419_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA1\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2930_ net504 net77 net41 VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2861_ matmult_inst.alu_inst.adder_inst.fa.b matmult_inst.alu_inst.adder_inst.fa.a
+ _1563_ VGND VGND VPWR VPWR _1565_ sky130_fd_sc_hd__a21o_1
XFILLER_30_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1812_ net280 _0682_ _0687_ net286 VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__a22o_1
X_2792_ _1506_ _1507_ VGND VGND VPWR VPWR _1508_ sky130_fd_sc_hd__xnor2_1
X_1743_ matmult_inst.mem_inst.matrixA2\[12\] net188 net180 matmult_inst.mem_inst.matrixA1\[12\]
+ _0625_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__a221o_1
X_1674_ matmult_inst.fsm_inst.rx_data\[0\] net468 matmult_inst.spi_inst.rx_done_sys
+ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__mux2_1
XFILLER_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold305 matmult_inst.mem_inst.mem1\[3\] VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 matmult_inst.mem_inst.mem1\[6\] VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__dlygate4sd3_1
X_3413_ clknet_leaf_26_hz100 net164 VGND VGND VPWR VPWR matmult_inst.alu_inst.complete
+ sky130_fd_sc_hd__dfxtp_1
Xhold349 matmult_inst.spi_inst.tx_reg_sys\[2\] VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 matmult_inst.spi_inst.tx_reg_sys\[3\] VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold327 matmult_inst.spi_inst.tx_reg_sys\[5\] VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__dlygate4sd3_1
X_3344_ clknet_leaf_6_hz100 _0209_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r0.fa3.b
+ sky130_fd_sc_hd__dfxtp_1
X_3275_ net291 _0017_ _0056_ VGND VGND VPWR VPWR matmult_inst.spi_inst.miso_shifter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2226_ _0892_ _0966_ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__nand2_1
XFILLER_38_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2157_ _0947_ net146 VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__xnor2_1
XFILLER_26_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2088_ net162 _0886_ _0887_ _0888_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_10_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_20_hz100 clknet_2_2__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_20_hz100
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_76_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3060_ net358 net80 net28 VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__mux2_1
X_2011_ matmult_inst.fsm_inst.alu_result\[16\] net113 VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__and2_1
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2913_ net482 _0816_ net43 VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2844_ net486 net9 net164 VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__mux2_1
X_2775_ matmult_inst.alu_inst.adder_inst.r0.fa3.b matmult_inst.alu_inst.adder_inst.r0.fa3.a
+ VGND VGND VPWR VPWR _1493_ sky130_fd_sc_hd__nand2_1
Xhold102 matmult_inst.mem_inst.matrixB1\[12\] VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 matmult_inst.mem_inst.matrixB0\[12\] VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 matmult_inst.mem_inst.matrixA0\[3\] VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__dlygate4sd3_1
X_1726_ net626 net92 _0610_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__o21a_1
Xhold135 matmult_inst.mem_inst.matrixA0\[6\] VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__dlygate4sd3_1
X_1657_ matmult_inst.spi_inst.rx_bit_count\[2\] net1 _0558_ matmult_inst.spi_inst.rx_done_spi
+ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__a31o_1
Xhold168 matmult_inst.mem_inst.matrixB2\[2\] VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 _0138_ VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 matmult_inst.alu_inst.adder_inst.r0.fa3.a VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 matmult_inst.mem_inst.matrixA3\[10\] VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__dlygate4sd3_1
X_3327_ _0100_ _0195_ _0099_ VGND VGND VPWR VPWR matmult_inst.spi_inst.mosi_data_spi\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3258_ clknet_leaf_10_hz100 _0147_ _0039_ VGND VGND VPWR VPWR matmult_inst.spi_inst.tx_reg_sys\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_3189_ net134 net123 VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__and2_1
XFILLER_66_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2209_ _1002_ _1004_ _1005_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_49_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2560_ _1283_ _1284_ net170 VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__o21ba_1
X_2491_ _1237_ _1238_ _1212_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__a21o_1
XFILLER_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3112_ net199 net166 _1595_ VGND VGND VPWR VPWR _1597_ sky130_fd_sc_hd__and3_1
XFILLER_55_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3043_ net333 net78 net30 VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2827_ matmult_inst.alu_inst.adder_inst.r2.fa3.b matmult_inst.alu_inst.adder_inst.r2.fa3.a
+ VGND VGND VPWR VPWR _1537_ sky130_fd_sc_hd__or2_1
X_2758_ net230 net577 net95 VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__mux2_1
X_1709_ matmult_inst.mem_inst.matrixA2\[15\] net188 net180 matmult_inst.mem_inst.matrixA1\[15\]
+ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__a22o_1
X_2689_ _1404_ net13 _1431_ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__nand3_1
XFILLER_48_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout30 _1590_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_4
Xfanout41 _1584_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_4
Xfanout74 _0817_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout85 _0806_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
Xfanout96 net100 VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1991_ matmult_inst.fsm_inst.rx_data\[6\] _0786_ net113 matmult_inst.fsm_inst.alu_result\[6\]
+ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__a22o_1
XFILLER_60_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3661_ clknet_leaf_18_hz100 _0521_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB2\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_2612_ net207 net209 net217 VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__and3_1
X_3592_ clknet_leaf_14_hz100 _0452_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA2\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload11 clknet_leaf_5_hz100 VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__inv_8
Xclkload22 clknet_leaf_9_hz100 VGND VGND VPWR VPWR clkload22/Y sky130_fd_sc_hd__inv_8
X_2543_ net212 net220 net218 net213 VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__nand4_1
X_2474_ net206 _1223_ _1222_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__a21bo_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3026_ net535 net76 net31 VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__mux2_1
XFILLER_55_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload5 clknet_leaf_29_hz100 VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__clkinvlp_4
Xwire109 net110 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout220 matmult_inst.alu_inst.a0_reg\[5\] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__buf_2
Xfanout231 matmult_inst.alu_inst.b1_reg\[7\] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_2
Xfanout264 net266 VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__buf_2
Xfanout242 matmult_inst.alu_inst.b1_reg\[1\] VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__buf_2
XFILLER_59_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout253 matmult_inst.alu_inst.a1_reg\[2\] VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__buf_2
Xfanout286 matmult_inst.fsm_inst.sel\[1\] VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__buf_2
Xfanout275 net276 VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__clkbuf_4
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2190_ _0984_ _0985_ _0986_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__nand3_1
XFILLER_37_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1974_ net308 net57 net21 matmult_inst.fsm_inst.alu_result\[16\] VGND VGND VPWR VPWR
+ _0139_ sky130_fd_sc_hd__a22o_1
XFILLER_60_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3644_ clknet_leaf_20_hz100 _0504_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB1\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_3575_ clknet_leaf_14_hz100 _0435_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA1\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_2526_ net141 net140 _1271_ _1270_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__o211ai_1
X_2457_ _1203_ _1204_ _1206_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__nand3_1
Xhold28 matmult_inst.mem_inst.matrixB3\[17\] VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 matmult_inst.mem_inst.mem3\[8\] VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2388_ _1158_ net379 _1161_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__mux2_1
Xhold39 matmult_inst.mem_inst.matrixA3\[9\] VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_71_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3009_ net528 _0817_ net33 VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1690_ matmult_inst.mem_inst.mem2\[17\] net192 net184 matmult_inst.mem_inst.mem1\[17\]
+ _0577_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__a221o_1
X_3360_ clknet_leaf_24_hz100 _0224_ VGND VGND VPWR VPWR matmult_inst.addr\[1\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_29_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2311_ net248 net246 net230 net233 VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__and4_1
X_3291_ clknet_leaf_5_hz100 net499 _0072_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.rx_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2242_ net251 net231 _1003_ _1005_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__a22o_1
X_2173_ _0927_ _0968_ _0969_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__nand3_1
XFILLER_65_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1957_ net58 _0799_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__nor2_1
X_1888_ matmult_inst.fsm_inst.state\[2\] net200 VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__nand2b_1
X_3627_ clknet_leaf_20_hz100 _0487_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB0\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_3558_ clknet_leaf_17_hz100 _0418_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA1\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2509_ _1243_ _1244_ net62 VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__o21ai_1
X_3489_ clknet_leaf_18_hz100 _0349_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem1\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_56_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2860_ net308 _1564_ net163 VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1811_ net196 _0683_ _0685_ net288 VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__a22o_1
X_2791_ _1497_ _1501_ _1498_ VGND VGND VPWR VPWR _1507_ sky130_fd_sc_hd__o21ai_1
X_1742_ net268 net261 matmult_inst.mem_inst.matrixA3\[12\] VGND VGND VPWR VPWR _0625_
+ sky130_fd_sc_hd__and3_1
Xhold306 matmult_inst.alu_inst.col0\[0\] VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold317 matmult_inst.alu_inst.adder_inst.r2.fa3.a VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__dlygate4sd3_1
X_1673_ matmult_inst.fsm_inst.rx_data\[1\] net565 matmult_inst.spi_inst.rx_done_sys
+ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__mux2_1
X_3412_ clknet_leaf_1_hz100 _0273_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.fa.a
+ sky130_fd_sc_hd__dfxtp_1
Xhold339 matmult_inst.spi_inst.tx_reg_sys\[0\] VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 matmult_inst.spi_inst.tx_reg_sys\[17\] VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_2_1__f_hz100 clknet_0_hz100 VGND VGND VPWR VPWR clknet_2_1__leaf_hz100 sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_1_hz100 clknet_2_1__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_1_hz100
+ sky130_fd_sc_hd__clkbuf_8
X_3343_ clknet_leaf_6_hz100 _0208_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r0.fa2.b
+ sky130_fd_sc_hd__dfxtp_1
X_3274_ net291 _0016_ _0055_ VGND VGND VPWR VPWR matmult_inst.spi_inst.miso_shifter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2225_ _0981_ _1019_ _1020_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__nand3_1
X_2156_ _0950_ _0951_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__xnor2_1
XFILLER_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2087_ matmult_inst.alu_inst.adder_inst.r1.fa1.b _0822_ VGND VGND VPWR VPWR _0888_
+ sky130_fd_sc_hd__and2_1
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2989_ net402 net75 net35 VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__mux2_1
XFILLER_16_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2010_ net324 net72 net55 VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__mux2_1
XFILLER_35_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2912_ net470 net76 net43 VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2843_ _1549_ net10 VGND VGND VPWR VPWR _1551_ sky130_fd_sc_hd__xnor2_1
X_2774_ matmult_inst.alu_inst.adder_inst.r0.fa3.b matmult_inst.alu_inst.adder_inst.r0.fa3.a
+ VGND VGND VPWR VPWR _1492_ sky130_fd_sc_hd__nor2_1
X_1725_ net279 _0604_ _0609_ _0602_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__a211o_1
Xhold114 matmult_inst.mem_inst.matrixA1\[17\] VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 matmult_inst.mem_inst.matrixA0\[7\] VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 matmult_inst.mem_inst.mem1\[7\] VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__dlygate4sd3_1
X_1656_ _0534_ matmult_inst.spi_inst.mosi_data_spi\[0\] _0562_ VGND VGND VPWR VPWR
+ _0194_ sky130_fd_sc_hd__mux2_1
Xhold147 matmult_inst.mem_inst.matrixA2\[0\] VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 matmult_inst.mem_inst.matrixB1\[5\] VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 matmult_inst.mem_inst.mem0\[9\] VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 matmult_inst.mem_inst.matrixA2\[8\] VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__dlygate4sd3_1
X_3326_ _0098_ _0194_ _0097_ VGND VGND VPWR VPWR matmult_inst.spi_inst.mosi_data_spi\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3257_ clknet_leaf_7_hz100 _0146_ _0038_ VGND VGND VPWR VPWR matmult_inst.spi_inst.tx_reg_sys\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2208_ net250 net235 VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__and2_1
X_3188_ net131 net120 VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_49_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2139_ _0933_ _0934_ _0936_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__and3_1
XFILLER_41_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2490_ _1212_ _1237_ _1238_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__nand3_1
XFILLER_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3111_ _1595_ VGND VGND VPWR VPWR _1596_ sky130_fd_sc_hd__inv_2
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3042_ net331 net79 net30 VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__mux2_1
XFILLER_16_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2826_ net466 net19 net164 VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__mux2_1
X_2757_ net233 net399 net95 VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__mux2_1
X_1708_ matmult_inst.mem_inst.matrixB2\[15\] net188 net180 matmult_inst.mem_inst.matrixB1\[15\]
+ _0593_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__a221o_1
XFILLER_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2688_ _1404_ _1431_ net13 VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__a21oi_1
X_1639_ net1 _0556_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__and2_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3309_ clknet_leaf_22_hz100 _0179_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB3\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout31 _1589_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_4
Xfanout42 _1584_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout75 _0816_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_2
Xfanout86 _0805_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_2
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1990_ net330 net82 net56 VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__mux2_1
X_3660_ clknet_leaf_21_hz100 _0520_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB2\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_3591_ clknet_leaf_22_hz100 _0451_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA2\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_2611_ net207 net219 net217 net209 VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__a22o_1
Xclkload12 clknet_leaf_6_hz100 VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__bufinv_16
Xclkload23 clknet_leaf_10_hz100 VGND VGND VPWR VPWR clkload23/Y sky130_fd_sc_hd__bufinv_16
X_2542_ net212 net220 net218 net213 VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__a22o_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2473_ net229 _1220_ net171 VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__and3_1
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3025_ net589 net77 net31 VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__mux2_1
XFILLER_51_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload6 clknet_leaf_30_hz100 VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__inv_12
X_2809_ matmult_inst.alu_inst.adder_inst.r2.fa0.b matmult_inst.alu_inst.adder_inst.r2.fa0.a
+ VGND VGND VPWR VPWR _1522_ sky130_fd_sc_hd__nand2_1
XFILLER_3_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout221 matmult_inst.alu_inst.a0_reg\[4\] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__buf_2
Xfanout210 matmult_inst.alu_inst.b0_reg\[3\] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout232 net233 VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__buf_2
Xfanout243 matmult_inst.alu_inst.b1_reg\[1\] VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_2
Xfanout254 matmult_inst.alu_inst.a1_reg\[2\] VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__buf_2
Xfanout265 net266 VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout287 net288 VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__clkbuf_4
Xfanout276 matmult_inst.spi_inst.first_bit_sent VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__clkbuf_4
XFILLER_46_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1973_ net450 net58 net21 matmult_inst.fsm_inst.alu_result\[15\] VGND VGND VPWR VPWR
+ _0138_ sky130_fd_sc_hd__a22o_1
X_3643_ clknet_leaf_18_hz100 _0503_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB1\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_3574_ clknet_leaf_14_hz100 _0434_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA1\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_2525_ _1270_ _1271_ net140 net141 VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__a211o_1
X_2456_ _1203_ _1204_ _1206_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__a21o_1
Xhold29 matmult_inst.mem_inst.mem3\[3\] VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 matmult_inst.mem_inst.mem3\[16\] VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2387_ _1157_ net493 _1161_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__mux2_1
XFILLER_68_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3008_ net567 net75 net33 VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2310_ _1103_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__inv_2
X_3290_ clknet_leaf_9_hz100 net566 _0071_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.rx_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2241_ net525 _1037_ net162 VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__mux2_1
XFILLER_38_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2172_ _0968_ _0969_ _0927_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__a21o_1
XFILLER_65_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1956_ _0537_ _0759_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__nor2_1
X_1887_ _0538_ matmult_inst.fsm_inst.state\[1\] matmult_inst.fsm_inst.state\[0\] VGND
+ VGND VPWR VPWR _0756_ sky130_fd_sc_hd__or3b_1
X_3626_ clknet_leaf_18_hz100 _0486_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB0\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_3557_ clknet_leaf_13_hz100 _0417_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA0\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_2508_ _1243_ _1244_ net62 VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__or3_1
X_3488_ clknet_leaf_24_hz100 _0348_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem1\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2439_ net226 net208 VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__and2_1
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap61 _1296_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
XFILLER_15_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1810_ matmult_inst.mem_inst.matrixB2\[6\] net189 net181 matmult_inst.mem_inst.matrixB1\[6\]
+ _0686_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__a221o_1
XFILLER_62_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2790_ _1503_ _1505_ VGND VGND VPWR VPWR _1506_ sky130_fd_sc_hd__nand2_1
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1741_ matmult_inst.mem_inst.matrixB2\[12\] net188 net180 matmult_inst.mem_inst.matrixB1\[12\]
+ _0623_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__a221o_1
XFILLER_7_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold307 matmult_inst.alu_inst.adder_inst.r1.fa2.b VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__dlygate4sd3_1
X_1672_ matmult_inst.fsm_inst.rx_data\[2\] net498 matmult_inst.spi_inst.rx_done_sys
+ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__mux2_1
X_3411_ clknet_leaf_31_hz100 _0272_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r3.fa3.a
+ sky130_fd_sc_hd__dfxtp_1
Xhold329 matmult_inst.alu_inst.adder_inst.fa.b VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 matmult_inst.alu_inst.out\[7\] VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__dlygate4sd3_1
X_3342_ clknet_leaf_6_hz100 _0207_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r0.fa1.b
+ sky130_fd_sc_hd__dfxtp_1
X_3273_ net291 _0015_ _0054_ VGND VGND VPWR VPWR matmult_inst.spi_inst.miso_shifter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2224_ _0981_ _1020_ _1019_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__a21o_1
X_2155_ _0950_ _0952_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__or2_1
XFILLER_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2086_ _0883_ _0884_ _0885_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__a21o_1
XFILLER_34_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2988_ net385 _0815_ net35 VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__mux2_1
X_1939_ matmult_inst.spi_inst.tx_reg_sys\[5\] matmult_inst.spi_inst.miso_shifter\[4\]
+ net276 VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__mux2_1
X_3609_ clknet_leaf_22_hz100 _0469_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA3\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_57_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Left_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2911_ net421 net77 net43 VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__mux2_1
XFILLER_73_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2842_ _1542_ _1545_ _1543_ VGND VGND VPWR VPWR _1550_ sky130_fd_sc_hd__a21boi_1
XPHY_EDGE_ROW_75_Left_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2773_ net424 _1491_ net164 VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__mux2_1
X_1724_ net283 _0606_ _0608_ net287 VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__a22o_1
XFILLER_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold115 matmult_inst.mem_inst.mem0\[15\] VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 matmult_inst.mem_inst.matrixA3\[13\] VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 matmult_inst.mem_inst.mem1\[4\] VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 matmult_inst.mem_inst.matrixA1\[1\] VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 matmult_inst.mem_inst.matrixA0\[14\] VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 matmult_inst.mem_inst.matrixA1\[4\] VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__dlygate4sd3_1
X_1655_ matmult_inst.spi_inst.mosi_shifter\[0\] matmult_inst.spi_inst.mosi_data_spi\[1\]
+ _0562_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__mux2_1
X_3325_ clknet_leaf_9_hz100 net295 _0096_ VGND VGND VPWR VPWR matmult_inst.spi_inst.cs_sync_prev
+ sky130_fd_sc_hd__dfstp_1
X_3256_ clknet_leaf_7_hz100 _0145_ _0037_ VGND VGND VPWR VPWR matmult_inst.spi_inst.tx_reg_sys\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2207_ net253 net251 net231 net232 VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__and4_1
X_3187_ net128 net117 VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__and2_1
XFILLER_66_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2138_ _0933_ _0934_ _0936_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__a21oi_1
X_2069_ _0868_ _0869_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__nand2_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_0_hz100 clknet_2_1__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_0_hz100
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_30_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3110_ net127 _1594_ VGND VGND VPWR VPWR _1595_ sky130_fd_sc_hd__and2_1
XFILLER_67_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3041_ net332 net80 net30 VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__mux2_1
XFILLER_63_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2825_ _1534_ net45 VGND VGND VPWR VPWR _1536_ sky130_fd_sc_hd__xnor2_1
X_2756_ net234 net384 net95 VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__mux2_1
X_1707_ net268 net261 matmult_inst.mem_inst.matrixB3\[15\] VGND VGND VPWR VPWR _0593_
+ sky130_fd_sc_hd__and3_1
X_2687_ _1402_ _1403_ _1386_ VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__o21bai_1
X_1638_ matmult_inst.spi_inst.rx_bit_count\[2\] matmult_inst.spi_inst.rx_bit_count\[1\]
+ matmult_inst.spi_inst.rx_bit_count\[0\] matmult_inst.spi_inst.rx_bit_count\[3\]
+ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__a31o_1
X_3308_ clknet_leaf_23_hz100 _0178_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB3\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_3239_ clknet_leaf_26_hz100 net301 VGND VGND VPWR VPWR matmult_inst.fsm_inst.alu_result\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout21 _0800_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_2
XFILLER_80_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout43 _1583_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_4
Xfanout32 _1589_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout76 _0815_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_2
Xfanout87 _0804_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload24 clknet_leaf_11_hz100 VGND VGND VPWR VPWR clkload24/Y sky130_fd_sc_hd__inv_12
X_2610_ net212 net216 VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__nand2_1
X_3590_ clknet_leaf_19_hz100 _0450_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA2\[14\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload13 clknet_leaf_17_hz100 VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__clkinv_2
X_2541_ net139 _1288_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__and2b_1
X_2472_ net206 net229 _1220_ net171 VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__a22o_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3024_ net449 net78 net32 VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__mux2_1
Xclkload7 clknet_leaf_31_hz100 VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__inv_12
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2808_ matmult_inst.alu_inst.adder_inst.r2.fa0.b matmult_inst.alu_inst.adder_inst.r2.fa0.a
+ VGND VGND VPWR VPWR _1521_ sky130_fd_sc_hd__nor2_1
X_2739_ net218 matmult_inst.alu_inst.a0_reg\[7\] net201 net203 _1476_ VGND VGND VPWR
+ VPWR _1479_ sky130_fd_sc_hd__a41o_1
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout200 matmult_inst.fsm_inst.state\[3\] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__buf_2
Xfanout222 net223 VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_2
Xfanout211 net212 VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout244 matmult_inst.alu_inst.b1_reg\[0\] VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__buf_2
Xfanout233 matmult_inst.alu_inst.b1_reg\[6\] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__buf_2
Xfanout255 matmult_inst.alu_inst.a1_reg\[1\] VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__buf_2
Xfanout288 matmult_inst.fsm_inst.sel\[0\] VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__clkbuf_4
Xfanout277 net279 VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__buf_2
Xfanout266 matmult_inst.addr\[1\] VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkbuf_2
XFILLER_75_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1972_ net300 net58 net21 matmult_inst.fsm_inst.alu_result\[14\] VGND VGND VPWR VPWR
+ _0137_ sky130_fd_sc_hd__a22o_1
X_3642_ clknet_leaf_21_hz100 _0502_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB1\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3573_ clknet_leaf_22_hz100 _0433_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA1\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2524_ _1221_ _1251_ _1252_ _1247_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__a31oi_1
X_2455_ _1183_ _1205_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__nor2_1
Xhold19 matmult_inst.mem_inst.matrixB3\[6\] VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__dlygate4sd3_1
X_2386_ _1156_ net377 _1161_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3007_ net503 net76 net33 VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__mux2_1
XFILLER_36_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2240_ _1035_ _1036_ _0998_ _1033_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__o2bb2a_1
X_2171_ net147 _0955_ net145 _0946_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__o211ai_2
XFILLER_53_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1955_ matmult_inst.fsm_inst.count\[1\] matmult_inst.fsm_inst.load_delay net156 _0783_
+ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__and4_1
X_1886_ matmult_inst.fsm_inst.state\[2\] _0754_ _0753_ _0548_ VGND VGND VPWR VPWR
+ _0755_ sky130_fd_sc_hd__a211o_1
X_3625_ clknet_leaf_18_hz100 _0485_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB0\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_3556_ clknet_leaf_14_hz100 _0416_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA0\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_2507_ _1247_ _1255_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__xnor2_1
X_3487_ clknet_leaf_24_hz100 _0347_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem1\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2438_ net440 net174 _1187_ _1189_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__a22o_1
X_2369_ _1154_ net554 _1152_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__mux2_1
XFILLER_56_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap51 _1226_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1740_ net268 net261 matmult_inst.mem_inst.matrixB3\[12\] VGND VGND VPWR VPWR _0623_
+ sky130_fd_sc_hd__and3_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold308 matmult_inst.alu_inst.out\[17\] VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__dlygate4sd3_1
X_1671_ matmult_inst.fsm_inst.rx_data\[3\] net592 matmult_inst.spi_inst.rx_done_sys
+ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__mux2_1
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3410_ clknet_leaf_31_hz100 _0271_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r3.fa2.a
+ sky130_fd_sc_hd__dfxtp_1
Xhold319 matmult_inst.alu_inst.row1\[2\] VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__dlygate4sd3_1
X_3341_ clknet_leaf_1_hz100 _0206_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r0.fa0.b
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3272_ net291 _0014_ _0053_ VGND VGND VPWR VPWR matmult_inst.spi_inst.miso_shifter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2223_ net158 _0979_ _0980_ _0987_ _0988_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__a32o_1
X_2154_ _0950_ _0952_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__nand2_1
XFILLER_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2085_ _0883_ _0884_ _0885_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_36_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2987_ net561 net77 net35 VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__mux2_1
X_1938_ matmult_inst.spi_inst.tx_reg_sys\[4\] matmult_inst.spi_inst.miso_shifter\[3\]
+ net276 VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__mux2_1
X_1869_ matmult_inst.mem_inst.matrixA0\[1\] net168 _0739_ _0740_ VGND VGND VPWR VPWR
+ _0741_ sky130_fd_sc_hd__a211o_1
X_3608_ clknet_leaf_19_hz100 _0468_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA3\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_3539_ clknet_leaf_13_hz100 _0399_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem3\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2910_ net452 net78 net44 VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__mux2_1
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2841_ _1547_ _1548_ VGND VGND VPWR VPWR _1549_ sky130_fd_sc_hd__and2b_1
XFILLER_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2772_ _1488_ _1490_ VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__xnor2_1
X_1723_ matmult_inst.mem_inst.matrixA2\[14\] net188 net180 matmult_inst.mem_inst.matrixA1\[14\]
+ _0607_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__a221o_1
Xhold116 matmult_inst.mem_inst.matrixA2\[1\] VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold105 matmult_inst.alu_inst.col1\[6\] VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 matmult_inst.mem_inst.mem0\[10\] VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 matmult_inst.mem_inst.mem0\[6\] VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 matmult_inst.mem_inst.mem1\[8\] VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__dlygate4sd3_1
X_1654_ matmult_inst.spi_inst.mosi_shifter\[1\] matmult_inst.spi_inst.mosi_data_spi\[2\]
+ _0562_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__mux2_1
X_3324_ _0095_ _0193_ _0094_ VGND VGND VPWR VPWR matmult_inst.spi_inst.rx_done_spi
+ sky130_fd_sc_hd__dfrtp_1
X_3255_ clknet_leaf_26_hz100 _0144_ _0036_ VGND VGND VPWR VPWR matmult_inst.spi_inst.tx_reg_sys\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2206_ net253 net231 net232 net251 VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__a22o_1
X_3186_ net127 net117 VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__and2_1
XFILLER_81_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2137_ _0896_ _0935_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__nand2_1
XFILLER_81_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2068_ net239 net254 net252 net240 VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_14_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3040_ net326 net81 net30 VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__mux2_1
XFILLER_75_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2824_ _1527_ _1530_ _1528_ VGND VGND VPWR VPWR _1535_ sky130_fd_sc_hd__o21ai_1
X_2755_ net237 net400 net96 VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__mux2_1
X_2686_ _1426_ _1429_ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__xnor2_1
X_1706_ matmult_inst.mem_inst.matrixA0\[15\] net168 _0591_ net194 net115 VGND VGND
+ VPWR VPWR _0592_ sky130_fd_sc_hd__a221o_1
X_1637_ net131 net120 VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__and2_1
X_3307_ clknet_leaf_21_hz100 _0177_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB3\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3238_ clknet_leaf_26_hz100 net487 VGND VGND VPWR VPWR matmult_inst.fsm_inst.alu_result\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_3169_ net136 net117 VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__and2_1
XFILLER_73_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout22 _0800_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
XFILLER_54_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout33 _1588_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_4
Xfanout55 _0803_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_4
Xfanout44 _1583_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout88 _0802_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout77 _0814_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload14 clknet_leaf_19_hz100 VGND VGND VPWR VPWR clkload14/Y sky130_fd_sc_hd__clkinv_8
Xclkload25 clknet_leaf_12_hz100 VGND VGND VPWR VPWR clkload25/Y sky130_fd_sc_hd__bufinv_16
X_2540_ _1281_ _1285_ _1286_ VGND VGND VPWR VPWR _1288_ sky130_fd_sc_hd__nand3_1
XFILLER_5_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2471_ net221 net220 net213 net215 VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__nand4_1
X_3023_ net463 net79 net32 VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__mux2_1
XFILLER_48_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload8 clknet_leaf_0_hz100 VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__inv_12
X_2807_ net612 _1520_ net163 VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__mux2_1
X_2738_ _1475_ _1476_ _1477_ _1478_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__o31ai_1
X_2669_ net205 net207 net217 net216 VGND VGND VPWR VPWR _1413_ sky130_fd_sc_hd__and4_1
Xfanout201 matmult_inst.alu_inst.b0_reg\[7\] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__buf_2
Xfanout223 matmult_inst.alu_inst.a0_reg\[3\] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__buf_2
Xfanout212 matmult_inst.alu_inst.b0_reg\[2\] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout245 matmult_inst.alu_inst.a1_reg\[7\] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__buf_2
Xfanout256 matmult_inst.alu_inst.a1_reg\[1\] VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__clkbuf_2
Xfanout234 matmult_inst.alu_inst.b1_reg\[5\] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__buf_2
Xfanout289 net290 VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__buf_4
Xfanout267 net270 VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__buf_2
Xfanout278 net279 VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__clkbuf_4
XFILLER_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1971_ net486 net58 net21 matmult_inst.fsm_inst.alu_result\[13\] VGND VGND VPWR VPWR
+ _0136_ sky130_fd_sc_hd__a22o_1
X_3641_ clknet_leaf_23_hz100 _0501_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB1\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3572_ clknet_leaf_19_hz100 _0432_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA1\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2523_ _1268_ _1269_ _1246_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__a21o_1
X_2454_ _1179_ _1184_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__nor2_1
X_2385_ _1155_ net613 _1161_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__mux2_1
Xinput1 cs VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
X_3006_ net428 net77 net33 VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__mux2_1
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2170_ _0946_ _0953_ _0954_ _0967_ net147 VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__a311o_1
XFILLER_38_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1954_ matmult_inst.fsm_inst.count\[1\] _0783_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__nand2_1
X_1885_ net200 _0551_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__nor2_1
X_3624_ clknet_leaf_21_hz100 _0484_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB0\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_3555_ clknet_leaf_21_hz100 _0415_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA0\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2506_ _1253_ _1254_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__nor2_1
X_3486_ clknet_leaf_17_hz100 _0346_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem1\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2437_ net174 _1188_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__nor2_1
X_2368_ _0741_ net167 VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__and2_1
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2299_ net506 _1093_ net159 VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap63 net64 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_2
Xmax_cap52 _1058_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
XFILLER_55_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1670_ matmult_inst.fsm_inst.rx_data\[4\] net522 matmult_inst.spi_inst.rx_done_sys
+ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__mux2_1
Xhold309 _0140_ VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__dlygate4sd3_1
X_3340_ clknet_leaf_24_hz100 matmult_inst.fsm_inst.tx_ready VGND VGND VPWR VPWR matmult_inst.fsm_inst.tx_ready_delay
+ sky130_fd_sc_hd__dfxtp_1
X_3271_ net291 _0007_ _0052_ VGND VGND VPWR VPWR matmult_inst.spi_inst.miso_shifter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2222_ _0985_ _0986_ _0984_ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__a21bo_1
X_2153_ matmult_inst.alu_inst.b1_reg\[0\] matmult_inst.alu_inst.a1_reg\[7\] VGND VGND
+ VPWR VPWR _0952_ sky130_fd_sc_hd__nand2_1
XFILLER_19_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2084_ _0844_ _0863_ _0864_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__a21bo_1
XFILLER_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2986_ net366 net78 net36 VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__mux2_1
X_1937_ matmult_inst.spi_inst.tx_reg_sys\[3\] matmult_inst.spi_inst.miso_shifter\[2\]
+ net276 VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__mux2_1
X_1868_ net287 _0733_ _0738_ net277 VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__a22o_1
X_3607_ clknet_leaf_18_hz100 _0467_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA3\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_3538_ clknet_leaf_15_hz100 _0398_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem3\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_1799_ matmult_inst.mem_inst.matrixA2\[7\] net189 net181 matmult_inst.mem_inst.matrixA1\[7\]
+ _0676_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__a221o_1
X_3469_ clknet_leaf_26_hz100 _0329_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem0\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2840_ matmult_inst.alu_inst.adder_inst.r3.fa1.b matmult_inst.alu_inst.adder_inst.r3.fa1.a
+ VGND VGND VPWR VPWR _1548_ sky130_fd_sc_hd__nand2_1
XFILLER_43_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2771_ _1482_ _1489_ VGND VGND VPWR VPWR _1490_ sky130_fd_sc_hd__or2_1
X_1722_ net269 net262 matmult_inst.mem_inst.matrixA3\[14\] VGND VGND VPWR VPWR _0607_
+ sky130_fd_sc_hd__and3_1
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold106 matmult_inst.alu_inst.col1\[4\] VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 matmult_inst.mem_inst.matrixA1\[9\] VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__dlygate4sd3_1
X_1653_ matmult_inst.spi_inst.mosi_shifter\[2\] matmult_inst.spi_inst.mosi_data_spi\[3\]
+ _0562_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__mux2_1
Xhold139 matmult_inst.mem_inst.mem2\[15\] VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold128 matmult_inst.mem_inst.matrixB0\[6\] VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__dlygate4sd3_1
X_3323_ clknet_leaf_8_hz100 _0192_ _0093_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.rx_valid
+ sky130_fd_sc_hd__dfrtp_1
X_3254_ clknet_leaf_26_hz100 _0143_ _0035_ VGND VGND VPWR VPWR matmult_inst.spi_inst.tx_reg_sys\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2205_ net253 net230 net232 net251 VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__a22oi_1
X_3185_ net128 net117 VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__and2_1
X_2136_ _0868_ _0897_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__nand2_1
XFILLER_81_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2067_ net239 net241 net254 net252 VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__nand4_2
XFILLER_81_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2969_ net350 net76 net37 VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__mux2_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2823_ _1532_ _1533_ VGND VGND VPWR VPWR _1534_ sky130_fd_sc_hd__nand2_1
X_2754_ net239 net579 net96 VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__mux2_1
X_1705_ net278 matmult_inst.mem_inst.mem0\[15\] matmult_inst.mem_inst.matrixB0\[15\]
+ net283 VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__a22o_1
X_2685_ _1427_ _1428_ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__or2_1
X_1636_ _0554_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__inv_2
X_3306_ clknet_leaf_12_hz100 _0176_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB3\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_3237_ clknet_leaf_26_hz100 net343 VGND VGND VPWR VPWR matmult_inst.fsm_inst.alu_result\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_3168_ net128 net117 VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__and2_1
XFILLER_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2119_ _0917_ _0918_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__nand2b_1
XFILLER_81_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3099_ net355 _0812_ net24 VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout23 _1593_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_4
Xfanout34 _1588_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_4
Xfanout56 _0803_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_4
Xfanout78 _0813_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload15 clknet_leaf_20_hz100 VGND VGND VPWR VPWR clkload15/Y sky130_fd_sc_hd__inv_8
Xclkload26 clknet_leaf_13_hz100 VGND VGND VPWR VPWR clkload26/Y sky130_fd_sc_hd__clkinv_4
XFILLER_5_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2470_ net221 net214 net215 net220 VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__a22o_1
XFILLER_48_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3022_ net531 net80 net32 VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload9 clknet_leaf_3_hz100 VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__inv_8
X_2806_ _1518_ _1519_ VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__xnor2_1
X_2737_ net607 net174 VGND VGND VPWR VPWR _1478_ sky130_fd_sc_hd__nand2_1
X_2668_ net205 net216 VGND VGND VPWR VPWR _1412_ sky130_fd_sc_hd__and2_1
X_1619_ matmult_inst.fsm_inst.state\[4\] _0536_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__nand2_1
X_2599_ _1309_ _1310_ _1308_ VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__a21bo_1
Xfanout202 matmult_inst.alu_inst.b0_reg\[7\] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_2
Xfanout213 matmult_inst.alu_inst.b0_reg\[1\] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout224 matmult_inst.alu_inst.a0_reg\[2\] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__buf_2
Xfanout246 matmult_inst.alu_inst.a1_reg\[6\] VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout235 matmult_inst.alu_inst.b1_reg\[5\] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_2
Xfanout268 net270 VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkbuf_2
Xfanout279 matmult_inst.fsm_inst.sel\[2\] VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__buf_2
Xfanout257 net259 VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_57_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1970_ net342 net58 net21 matmult_inst.fsm_inst.alu_result\[12\] VGND VGND VPWR VPWR
+ _0135_ sky130_fd_sc_hd__a22o_1
X_3640_ clknet_leaf_21_hz100 _0500_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB1\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3571_ clknet_leaf_18_hz100 _0431_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA1\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_2522_ _1246_ _1268_ _1269_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__nand3_2
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2453_ _1195_ _1196_ net143 VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__or3b_1
X_2384_ _1154_ net456 _1161_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__mux2_1
Xinput2 mosi VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
X_3005_ net411 net78 net34 VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__mux2_1
XFILLER_51_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1953_ net655 net297 VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__nor2_1
X_1884_ matmult_inst.fsm_inst.state\[0\] _0550_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__nor2_1
X_3623_ clknet_leaf_25_hz100 _0483_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB0\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_3554_ clknet_leaf_18_hz100 _0414_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA0\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_2505_ _1251_ _1252_ _1221_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__a21oi_1
X_3485_ clknet_leaf_15_hz100 _0345_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem0\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_2436_ _1172_ _1175_ _1186_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__o21a_1
X_2367_ _1153_ net576 _1152_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__mux2_1
X_2298_ _1090_ _1092_ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_67_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap20 _1334_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
Xmax_cap64 _1165_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_2
XFILLER_62_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3270_ net292 net294 _0051_ VGND VGND VPWR VPWR matmult_inst.spi_inst.first_bit_sent
+ sky130_fd_sc_hd__dfrtp_1
X_2221_ _0926_ _0968_ _0969_ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__a21bo_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2152_ matmult_inst.alu_inst.b1_reg\[0\] matmult_inst.alu_inst.a1_reg\[7\] VGND VGND
+ VPWR VPWR _0951_ sky130_fd_sc_hd__and2_1
X_2083_ _0867_ net54 VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__or2_1
XFILLER_19_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2985_ net490 net79 net36 VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__mux2_1
X_1936_ matmult_inst.spi_inst.tx_reg_sys\[2\] matmult_inst.spi_inst.miso_shifter\[1\]
+ net276 VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__mux2_1
X_1867_ net194 _0734_ _0736_ net284 VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__a22o_1
X_3606_ clknet_leaf_22_hz100 _0466_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA3\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_1798_ net274 net263 matmult_inst.mem_inst.matrixA3\[7\] VGND VGND VPWR VPWR _0676_
+ sky130_fd_sc_hd__and3_1
X_3537_ clknet_leaf_22_hz100 _0397_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem3\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_3468_ clknet_leaf_17_hz100 _0328_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem0\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2419_ _1170_ _1171_ net228 net211 VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__and4bb_1
X_3399_ clknet_leaf_1_hz100 _0260_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r0.fa3.a
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_69_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_26_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2770_ matmult_inst.alu_inst.adder_inst.r0.fa1.b matmult_inst.alu_inst.adder_inst.r0.fa1.a
+ matmult_inst.alu_inst.adder_inst.r0.fa0.b matmult_inst.alu_inst.adder_inst.r0.fa0.a
+ VGND VGND VPWR VPWR _1489_ sky130_fd_sc_hd__a22oi_1
X_1721_ matmult_inst.mem_inst.matrixB2\[14\] net193 net185 matmult_inst.mem_inst.matrixB1\[14\]
+ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_44_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold107 matmult_inst.mem_inst.matrixB1\[17\] VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__dlygate4sd3_1
X_1652_ matmult_inst.spi_inst.mosi_shifter\[3\] matmult_inst.spi_inst.mosi_data_spi\[4\]
+ _0562_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__mux2_1
Xhold129 matmult_inst.mem_inst.matrixA3\[15\] VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 matmult_inst.alu_inst.adder_inst.r3.fa0.b VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__dlygate4sd3_1
X_3322_ _0092_ _0191_ _0091_ VGND VGND VPWR VPWR matmult_inst.spi_inst.mosi_shifter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_3253_ clknet_leaf_26_hz100 _0142_ _0034_ VGND VGND VPWR VPWR matmult_inst.spi_inst.tx_reg_sys\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2204_ _0977_ _0978_ _0976_ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__a21bo_1
X_3184_ net135 net125 VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_53_Left_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2135_ _0931_ _0932_ _0894_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_49_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2066_ _0851_ _0858_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_31_hz100 clknet_2_0__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_31_hz100
+ sky130_fd_sc_hd__clkbuf_8
X_2968_ net321 net77 net37 VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1919_ net282 _0785_ _0786_ _0775_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_62_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2899_ net652 _1578_ _1582_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__o21a_1
XFILLER_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Left_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_80_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2822_ matmult_inst.alu_inst.adder_inst.r2.fa2.b matmult_inst.alu_inst.adder_inst.r2.fa2.a
+ VGND VGND VPWR VPWR _1533_ sky130_fd_sc_hd__nand2_1
X_2753_ net241 net386 net96 VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__mux2_1
X_1704_ net628 net91 _0582_ _0590_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__o22a_1
X_2684_ net219 net201 _1388_ VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__and3_1
X_1635_ _0540_ _0542_ net197 VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__nand3_2
X_3305_ clknet_leaf_10_hz100 _0175_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB3\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3236_ clknet_leaf_26_hz100 net477 VGND VGND VPWR VPWR matmult_inst.fsm_inst.alu_result\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_3167_ net128 net117 VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__and2_1
XFILLER_39_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3098_ net609 _0811_ net24 VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__mux2_1
X_2118_ _0889_ _0915_ _0916_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__nand3_1
XFILLER_81_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2049_ _0849_ _0850_ _0838_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__a21oi_1
XFILLER_81_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout35 _1587_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_4
Xfanout24 _1593_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout57 net58 VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_2
Xfanout79 _0812_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_51 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload16 clknet_leaf_21_hz100 VGND VGND VPWR VPWR clkload16/Y sky130_fd_sc_hd__clkinv_4
Xclkload27 clknet_leaf_14_hz100 VGND VGND VPWR VPWR clkload27/Y sky130_fd_sc_hd__inv_6
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3021_ net538 net81 net32 VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__mux2_1
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2805_ _1509_ _1513_ _1510_ VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_14_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2736_ _1468_ _1473_ _1474_ VGND VGND VPWR VPWR _1477_ sky130_fd_sc_hd__a21oi_1
X_2667_ net551 _1411_ net160 VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__mux2_1
X_1618_ net199 net200 VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__or2_2
Xfanout203 matmult_inst.alu_inst.b0_reg\[6\] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__buf_2
Xfanout214 matmult_inst.alu_inst.b0_reg\[1\] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__dlymetal6s2s_1
X_2598_ net159 _1342_ _1343_ _1344_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__a31o_1
Xfanout225 matmult_inst.alu_inst.a0_reg\[2\] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout236 net237 VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__buf_2
Xfanout247 matmult_inst.alu_inst.a1_reg\[6\] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_2
Xfanout269 net270 VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__buf_1
Xfanout258 net259 VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__buf_1
XFILLER_74_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3219_ net292 VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__inv_2
XFILLER_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold290 matmult_inst.mem_inst.mem3\[13\] VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3570_ clknet_leaf_22_hz100 _0430_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA1\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2521_ net229 net227 net202 net204 VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__nand4_1
XFILLER_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2452_ _1195_ _1196_ net143 VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__o21bai_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2383_ _1153_ net389 _1161_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__mux2_1
XFILLER_56_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput3 spi_clk VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
X_3004_ net505 net79 net34 VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2719_ net217 net216 net201 net203 VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__nand4_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1952_ net653 net296 VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__and2b_1
X_1883_ matmult_inst.fsm_inst.state\[1\] matmult_inst.fsm_inst.state\[0\] VGND VGND
+ VPWR VPWR _0752_ sky130_fd_sc_hd__nor2_1
X_3622_ clknet_leaf_20_hz100 _0482_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB0\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3553_ clknet_leaf_18_hz100 _0413_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA0\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_2504_ _1221_ _1251_ _1252_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__and3_1
X_3484_ clknet_leaf_15_hz100 _0344_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem0\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_2435_ _1172_ _1175_ _1186_ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__or3_1
X_2366_ _0751_ net167 VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2297_ _1066_ _1091_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap10 _1550_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
Xmax_cap54 _0882_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_1
Xmax_cap65 net66 VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_2
XFILLER_43_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2220_ _1011_ net144 VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__xor2_1
X_2151_ net247 _0906_ _0948_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__a21bo_1
X_2082_ _0867_ _0882_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__nand2_1
XFILLER_19_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2984_ net419 net80 net36 VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1935_ matmult_inst.spi_inst.tx_reg_sys\[1\] matmult_inst.spi_inst.miso_shifter\[0\]
+ net276 VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__mux2_1
X_1866_ matmult_inst.mem_inst.mem2\[1\] net186 net178 matmult_inst.mem_inst.mem1\[1\]
+ _0737_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__a221o_1
X_3605_ clknet_leaf_23_hz100 _0465_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA3\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_1797_ matmult_inst.mem_inst.matrixB2\[7\] net189 net181 matmult_inst.mem_inst.matrixB1\[7\]
+ _0674_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__a221o_1
X_3536_ clknet_leaf_18_hz100 _0396_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem3\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_3467_ clknet_leaf_28_hz100 _0327_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.count\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2418_ net227 net225 net214 net215 VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__and4_1
X_3398_ clknet_leaf_1_hz100 _0259_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r0.fa2.a
+ sky130_fd_sc_hd__dfxtp_1
X_2349_ matmult_inst.alu_inst.complete _0551_ _0763_ _1137_ VGND VGND VPWR VPWR _1138_
+ sky130_fd_sc_hd__o31a_1
XFILLER_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1720_ net269 net262 matmult_inst.mem_inst.matrixB3\[14\] VGND VGND VPWR VPWR _0605_
+ sky130_fd_sc_hd__and3_1
Xhold108 matmult_inst.mem_inst.matrixA0\[12\] VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__dlygate4sd3_1
X_1651_ matmult_inst.spi_inst.mosi_shifter\[4\] matmult_inst.spi_inst.mosi_data_spi\[5\]
+ _0562_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__mux2_1
Xhold119 matmult_inst.mem_inst.matrixA0\[0\] VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__dlygate4sd3_1
X_3321_ _0090_ _0190_ _0089_ VGND VGND VPWR VPWR matmult_inst.spi_inst.mosi_shifter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3252_ clknet_leaf_17_hz100 _0141_ _0033_ VGND VGND VPWR VPWR matmult_inst.spi_inst.tx_reg_sys\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2203_ net624 _1000_ net161 VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__mux2_1
XFILLER_66_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3183_ net135 net124 VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__and2_1
X_2134_ _0894_ _0931_ _0932_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__nand3_1
XFILLER_26_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2065_ net605 _0866_ net162 VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__mux2_1
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2967_ net329 net78 net38 VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__mux2_1
X_1918_ matmult_inst.fsm_inst.count\[1\] matmult_inst.fsm_inst.count\[0\] VGND VGND
+ VPWR VPWR _0787_ sky130_fd_sc_hd__xor2_1
X_2898_ matmult_inst.fsm_inst.count\[3\] _1578_ _1581_ _1571_ VGND VGND VPWR VPWR
+ _1582_ sky130_fd_sc_hd__o2bb2a_1
X_1849_ net267 net260 matmult_inst.mem_inst.mem3\[2\] VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__and3_1
XFILLER_78_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3519_ clknet_leaf_22_hz100 _0379_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem2\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2821_ matmult_inst.alu_inst.adder_inst.r2.fa2.b matmult_inst.alu_inst.adder_inst.r2.fa2.a
+ VGND VGND VPWR VPWR _1532_ sky130_fd_sc_hd__or2_1
X_2752_ net243 net547 net96 VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__mux2_1
XFILLER_76_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1703_ net288 _0584_ _0589_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__a21o_1
X_2683_ net221 net201 net203 net219 VGND VGND VPWR VPWR _1427_ sky130_fd_sc_hd__a22oi_1
X_1634_ matmult_inst.fsm_inst.rx_ready_edge_delay net154 net155 VGND VGND VPWR VPWR
+ _0553_ sky130_fd_sc_hd__a21oi_2
X_3304_ clknet_leaf_10_hz100 _0174_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB3\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_3235_ clknet_leaf_26_hz100 net467 VGND VGND VPWR VPWR matmult_inst.fsm_inst.alu_result\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3166_ net128 net117 VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__and2_1
XFILLER_66_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3097_ net586 net81 net24 VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__mux2_1
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2117_ _0915_ _0916_ _0889_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__a21oi_1
XFILLER_81_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2048_ _0847_ _0848_ _0835_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_80_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout25 _1592_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_4
Xfanout36 _1587_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_4
Xfanout58 _0794_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_2
XFILLER_22_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload17 clknet_leaf_22_hz100 VGND VGND VPWR VPWR clkload17/Y sky130_fd_sc_hd__inv_6
XFILLER_70_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload28 clknet_leaf_15_hz100 VGND VGND VPWR VPWR clkload28/Y sky130_fd_sc_hd__inv_6
XFILLER_62_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_30_hz100 clknet_2_0__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_30_hz100
+ sky130_fd_sc_hd__clkbuf_8
X_3020_ net556 net82 net32 VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2804_ _1515_ _1517_ VGND VGND VPWR VPWR _1518_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_14_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2735_ _1439_ _1463_ _1446_ matmult_inst.alu_inst.a0_reg\[7\] net201 VGND VGND VPWR
+ VPWR _1476_ sky130_fd_sc_hd__o2111a_1
X_2666_ _1409_ _1410_ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__xnor2_1
X_1617_ net199 net200 VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__nor2_1
Xfanout204 matmult_inst.alu_inst.b0_reg\[6\] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__buf_2
X_2597_ matmult_inst.alu_inst.adder_inst.r2.fa0.a net174 VGND VGND VPWR VPWR _1344_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_6_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout215 matmult_inst.alu_inst.b0_reg\[0\] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__buf_2
Xfanout226 net227 VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__buf_2
Xfanout237 matmult_inst.alu_inst.b1_reg\[4\] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__buf_2
Xfanout259 matmult_inst.alu_inst.a1_reg\[0\] VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__clkbuf_2
Xfanout248 matmult_inst.alu_inst.a1_reg\[5\] VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__buf_2
X_3218_ net290 VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__inv_2
XFILLER_39_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3149_ net130 net122 VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__and2_1
XFILLER_54_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold280 matmult_inst.mem_inst.matrixB1\[1\] VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold291 matmult_inst.mem_inst.matrixB1\[14\] VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2520_ net229 net202 net204 net227 VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__a22o_1
XFILLER_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2451_ _1196_ net143 VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__nor2_1
X_2382_ _0537_ _0759_ _0766_ _0564_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__o22a_4
X_3003_ net471 net80 net34 VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2718_ net217 net201 net203 net216 VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__a22o_1
X_2649_ _1390_ _1391_ _1392_ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__or3b_1
XFILLER_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270__294 VGND VGND VPWR VPWR net294 _3270__294/LO sky130_fd_sc_hd__conb_1
XFILLER_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1951_ matmult_inst.spi_inst.current_state matmult_inst.spi_inst.cs_sync_prev _0797_
+ VGND VGND VPWR VPWR matmult_inst.spi_inst.next_state sky130_fd_sc_hd__o21a_1
X_1882_ net298 _0533_ matmult_inst.spi_inst.rx_done_sys VGND VGND VPWR VPWR _0122_
+ sky130_fd_sc_hd__a21o_1
X_3621_ clknet_leaf_13_hz100 _0481_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB0\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_3552_ clknet_leaf_21_hz100 _0412_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA0\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_2503_ _1249_ _1250_ _1248_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__a21o_1
X_3483_ clknet_leaf_21_hz100 _0343_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem0\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_2434_ _1179_ _1185_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__xnor2_1
X_2365_ _0791_ net150 VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__nor2_1
X_2296_ _0996_ _0997_ _1033_ _1034_ _1065_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_67_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_6_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap66 _1163_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_2
XFILLER_62_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2150_ net240 net242 net249 net247 VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__and4_1
XFILLER_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2081_ _0875_ net112 VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2983_ net429 _0810_ net36 VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1934_ net276 matmult_inst.spi_inst.tx_reg_sys\[0\] VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__and2b_1
X_1865_ net267 net260 matmult_inst.mem_inst.mem3\[1\] VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__and3_1
X_3604_ clknet_leaf_20_hz100 _0464_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA3\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_1796_ net273 net265 matmult_inst.mem_inst.matrixB3\[7\] VGND VGND VPWR VPWR _0674_
+ sky130_fd_sc_hd__and3_1
X_3535_ clknet_leaf_18_hz100 _0395_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem3\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_3466_ clknet_leaf_28_hz100 _0326_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.count\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2417_ net226 net214 net215 net225 VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__a22oi_1
X_3397_ clknet_leaf_1_hz100 _0258_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r0.fa1.a
+ sky130_fd_sc_hd__dfxtp_1
X_2348_ net156 _0545_ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__nand2_1
X_2279_ _1072_ _1073_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_27_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1650_ matmult_inst.spi_inst.mosi_shifter\[5\] matmult_inst.spi_inst.mosi_data_spi\[6\]
+ _0562_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__mux2_1
XFILLER_11_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold109 matmult_inst.mem_inst.matrixA1\[2\] VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__dlygate4sd3_1
X_3320_ _0088_ _0189_ _0087_ VGND VGND VPWR VPWR matmult_inst.spi_inst.mosi_shifter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3251_ net293 _0006_ _0032_ VGND VGND VPWR VPWR matmult_inst.spi_inst.miso_bit sky130_fd_sc_hd__dfrtp_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2202_ _0964_ _0999_ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__xnor2_1
X_3182_ net135 net124 VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__and2_1
XFILLER_66_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2133_ _0912_ _0930_ _0929_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__a21o_1
XFILLER_81_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2064_ _0844_ _0865_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__xnor2_1
X_2966_ net311 net79 net38 VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__mux2_1
X_2897_ _0771_ net166 net152 VGND VGND VPWR VPWR _1581_ sky130_fd_sc_hd__mux2_1
X_1917_ matmult_inst.fsm_inst.rx_ready_edge_delay matmult_inst.fsm_inst.rx_ready_edge
+ net154 _0771_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__and4b_4
X_1848_ net632 _0721_ net92 VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__mux2_1
X_1779_ net286 _0656_ _0658_ net280 VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__a22o_1
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3518_ clknet_leaf_19_hz100 _0378_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem2\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_3449_ clknet_leaf_27_hz100 _0309_ VGND VGND VPWR VPWR matmult_inst.alu_inst.a0_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2820_ net391 net46 net163 VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__mux2_1
X_2751_ net244 net448 net95 VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__mux2_1
X_2682_ _1424_ _1425_ VGND VGND VPWR VPWR _1426_ sky130_fd_sc_hd__nand2b_1
X_1702_ net286 _0586_ _0588_ net280 VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__a22o_1
X_1633_ _0537_ _0551_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__nor2_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3303_ clknet_leaf_16_hz100 _0173_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB3\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3234_ clknet_leaf_7_hz100 net392 VGND VGND VPWR VPWR matmult_inst.fsm_inst.alu_result\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_3165_ net135 net124 VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__and2_1
X_3096_ net553 _0809_ net24 VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__mux2_1
X_2116_ _0900_ _0901_ net69 VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__or3_1
X_2047_ _0835_ _0847_ _0848_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_80_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout37 _1586_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_4
Xfanout26 _1592_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2949_ net370 net77 net39 VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__mux2_1
Xmax_cap170 _1282_ VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload18 clknet_leaf_23_hz100 VGND VGND VPWR VPWR clkload18/Y sky130_fd_sc_hd__inv_6
Xclkload29 clknet_leaf_16_hz100 VGND VGND VPWR VPWR clkload29/Y sky130_fd_sc_hd__bufinv_16
XFILLER_70_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2803_ matmult_inst.alu_inst.adder_inst.r1.fa3.b matmult_inst.alu_inst.adder_inst.r1.fa3.a
+ VGND VGND VPWR VPWR _1517_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_14_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2734_ _1468_ _1473_ _1474_ net174 VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__a31o_1
X_2665_ _1339_ _1376_ _1380_ net14 VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__a31o_1
X_1616_ net268 net261 VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__and2_1
X_2596_ net17 _1340_ _1341_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__o21ai_1
XFILLER_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout205 matmult_inst.alu_inst.b0_reg\[5\] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__buf_2
Xfanout216 matmult_inst.alu_inst.a0_reg\[7\] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout227 matmult_inst.alu_inst.a0_reg\[1\] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_2
Xfanout238 matmult_inst.alu_inst.b1_reg\[3\] VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__buf_2
Xfanout249 matmult_inst.alu_inst.a1_reg\[5\] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__clkbuf_2
X_3217_ net292 VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__inv_2
X_3148_ net130 net122 VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__and2_1
X_3079_ net597 _0811_ net26 VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_59_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_68_Left_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold270 matmult_inst.mem_inst.mem2\[3\] VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold281 matmult_inst.mem_inst.matrixB2\[13\] VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 matmult_inst.mem_inst.matrixB2\[6\] VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2450_ _1197_ _1200_ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__xnor2_1
X_2381_ _1160_ net527 net108 VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__mux2_1
X_3002_ net542 net81 net34 VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__mux2_1
XFILLER_51_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2717_ net615 _1459_ net160 VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__mux2_1
XFILLER_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2648_ _1390_ _1391_ _1392_ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__o21bai_1
X_2579_ _1288_ _1295_ _1325_ _1287_ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__a211o_1
XFILLER_42_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1950_ matmult_inst.spi_inst.current_state matmult_inst.spi_inst.cs_sync_prev matmult_inst.spi_inst.cs_sync
+ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__a21bo_1
X_1881_ net633 _0751_ net92 VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__mux2_1
X_3620_ clknet_leaf_16_hz100 _0480_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB0\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3551_ clknet_leaf_23_hz100 _0411_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA0\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_2502_ _1248_ _1249_ _1250_ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__nand3_1
X_3482_ clknet_leaf_18_hz100 _0342_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem0\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2433_ _1183_ _1184_ VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__or2_1
X_2364_ _1141_ _1149_ _1151_ _1139_ net260 VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__o32a_1
X_2295_ _1088_ _1089_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_67_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap12 _1454_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_1
Xmax_cap67 _0990_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_1
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap89 net90 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_1
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2080_ _0846_ _0880_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__xnor2_1
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2982_ net375 net82 net36 VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__mux2_1
X_1933_ matmult_inst.spi_inst.tx_reg_sys\[16\] matmult_inst.spi_inst.miso_shifter\[15\]
+ net275 VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__mux2_1
X_1864_ matmult_inst.mem_inst.matrixB2\[1\] net187 net179 matmult_inst.mem_inst.matrixB1\[1\]
+ _0735_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__a221o_1
X_3603_ clknet_leaf_12_hz100 _0463_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA3\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_1795_ net281 matmult_inst.mem_inst.mem0\[7\] matmult_inst.mem_inst.matrixB0\[7\]
+ net285 VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__a22o_1
X_3534_ clknet_leaf_22_hz100 _0394_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem3\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_3465_ clknet_leaf_24_hz100 _0325_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.count\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2416_ net651 net175 _1167_ _1169_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__a22o_1
X_3396_ clknet_leaf_1_hz100 _0257_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r0.fa0.a
+ sky130_fd_sc_hd__dfxtp_1
X_2347_ matmult_inst.fsm_inst.tx_start_send _0554_ _0773_ VGND VGND VPWR VPWR _1136_
+ sky130_fd_sc_hd__o21bai_1
X_2278_ _1047_ _1048_ net172 VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_27_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3250_ clknet_leaf_9_hz100 matmult_inst.spi_inst.mosi_data_spi\[7\] _0031_ VGND VGND
+ VPWR VPWR matmult_inst.spi_inst.mosi_data_sync\[7\] sky130_fd_sc_hd__dfrtp_1
X_2201_ _0995_ _0996_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__nand2b_1
X_3181_ net135 net124 VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_77_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2132_ _0912_ _0929_ _0930_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__nand3_1
XFILLER_19_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2063_ _0863_ _0864_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_22_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2965_ net315 net80 net38 VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__mux2_1
X_2896_ _1580_ matmult_inst.fsm_inst.count\[2\] _1571_ VGND VGND VPWR VPWR _0326_
+ sky130_fd_sc_hd__mux2_1
X_1916_ net156 _0784_ _0782_ _0776_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__a211o_1
X_1847_ matmult_inst.mem_inst.matrixA0\[3\] net168 _0719_ _0720_ VGND VGND VPWR VPWR
+ _0721_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_31_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3517_ clknet_leaf_18_hz100 _0377_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem2\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_1778_ matmult_inst.mem_inst.mem2\[9\] net191 net183 matmult_inst.mem_inst.mem1\[9\]
+ _0657_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__a221o_1
X_3448_ clknet_leaf_27_hz100 _0308_ VGND VGND VPWR VPWR matmult_inst.alu_inst.a0_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3379_ clknet_leaf_29_hz100 _0241_ VGND VGND VPWR VPWR matmult_inst.alu_inst.col0\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_40_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2750_ net245 net544 net95 VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__mux2_1
X_2681_ _1400_ _1423_ VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__or2_1
X_1701_ matmult_inst.mem_inst.mem2\[16\] net191 net183 matmult_inst.mem_inst.mem1\[16\]
+ _0587_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__a221o_1
XFILLER_8_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1632_ matmult_inst.fsm_inst.state\[4\] _0549_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__or2_2
X_3302_ clknet_leaf_17_hz100 _0172_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB3\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3233_ clknet_leaf_7_hz100 net581 VGND VGND VPWR VPWR matmult_inst.fsm_inst.alu_result\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3164_ net134 net123 VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__and2_1
XFILLER_66_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3095_ net495 net83 net24 VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__mux2_1
X_2115_ _0900_ _0901_ net69 VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__o21ai_1
XFILLER_66_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2046_ net239 net256 net237 net258 VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_80_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout27 _1591_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_4
Xfanout38 _1586_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2948_ net444 net78 net40 VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__mux2_1
X_2879_ net202 net533 net93 VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap171 _1221_ VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__buf_1
XFILLER_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload19 clknet_leaf_24_hz100 VGND VGND VPWR VPWR clkload19/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2802_ _1515_ VGND VGND VPWR VPWR _1516_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2733_ matmult_inst.alu_inst.a0_reg\[7\] net201 _1446_ _1463_ _1439_ VGND VGND VPWR
+ VPWR _1474_ sky130_fd_sc_hd__a311o_1
X_2664_ _1407_ _1408_ VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__nor2_1
X_1615_ net289 VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__inv_2
X_2595_ net17 _1340_ _1341_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__or3_1
Xfanout217 matmult_inst.alu_inst.a0_reg\[6\] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__buf_2
Xfanout206 matmult_inst.alu_inst.b0_reg\[5\] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout228 net229 VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_2
Xfanout239 matmult_inst.alu_inst.b1_reg\[3\] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__clkbuf_2
X_3216_ net131 net120 VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__and2_1
XFILLER_39_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3147_ net130 net118 VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__and2_1
X_3078_ net368 net81 net26 VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__mux2_1
X_2029_ _0825_ _0831_ net162 VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__o21ai_1
XFILLER_24_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold260 matmult_inst.alu_inst.row0\[1\] VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 matmult_inst.spi_inst.mosi_data_sync\[1\] VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold282 matmult_inst.alu_inst.row0\[0\] VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 matmult_inst.mem_inst.matrixB2\[10\] VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2380_ _0680_ net167 VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__and2_2
XFILLER_36_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3001_ net491 net82 net34 VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__mux2_1
XFILLER_24_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2716_ _1456_ _1458_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__xor2_1
X_2647_ net209 net216 VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__nand2_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2578_ _1323_ _1324_ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__xnor2_1
XFILLER_27_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1880_ matmult_inst.mem_inst.matrixA0\[0\] net169 _0749_ _0750_ VGND VGND VPWR VPWR
+ _0751_ sky130_fd_sc_hd__a211o_1
X_3550_ clknet_leaf_20_hz100 _0410_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA0\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_2501_ net211 net221 net220 net213 VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__nand4_1
X_3481_ clknet_leaf_18_hz100 _0341_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem0\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_2432_ _1171_ _1181_ _1182_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2363_ net89 net176 net109 _0764_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__a211o_1
X_2294_ _1086_ _1087_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__nand2_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2981_ net427 net83 net36 VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__mux2_1
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1932_ matmult_inst.spi_inst.tx_reg_sys\[17\] matmult_inst.spi_inst.miso_bit net275
+ VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__mux2_1
X_1863_ net270 net260 matmult_inst.mem_inst.matrixB3\[1\] VGND VGND VPWR VPWR _0735_
+ sky130_fd_sc_hd__and3_1
X_3602_ clknet_leaf_12_hz100 _0462_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA3\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_1794_ matmult_inst.mem_inst.mem2\[7\] net189 net181 matmult_inst.mem_inst.mem1\[7\]
+ _0671_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__a221o_1
X_3533_ clknet_leaf_23_hz100 _0393_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem3\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_3464_ clknet_leaf_28_hz100 _0324_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.count\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2415_ net174 _1168_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__nor2_1
X_3395_ clknet_leaf_25_hz100 net299 VGND VGND VPWR VPWR matmult_inst.fsm_inst.rx_ready_edge_delay
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2346_ net623 net175 VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__and2_1
X_2277_ _1070_ _1071_ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_27_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2200_ _0996_ _0997_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__and2_1
X_3180_ net136 net125 VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_77_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2131_ _0877_ _0909_ _0910_ _0904_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__a31o_1
XFILLER_81_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2062_ _0859_ _0860_ _0862_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__nand3_1
XFILLER_81_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2964_ net383 net81 net37 VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__mux2_1
X_1915_ _0543_ net177 VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2895_ _1572_ _1577_ _1579_ VGND VGND VPWR VPWR _1580_ sky130_fd_sc_hd__and3_1
X_1846_ net287 _0713_ _0718_ net284 VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__a22o_1
X_1777_ net273 net265 matmult_inst.mem_inst.mem3\[9\] VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__and3_1
X_3516_ clknet_leaf_22_hz100 _0376_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem2\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3447_ clknet_leaf_1_hz100 _0307_ VGND VGND VPWR VPWR matmult_inst.alu_inst.out\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_3378_ clknet_leaf_24_hz100 _0005_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.tx_start_send
+ sky130_fd_sc_hd__dfxtp_1
X_2329_ _1099_ net111 VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__or2_1
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2680_ _1400_ _1423_ VGND VGND VPWR VPWR _1424_ sky130_fd_sc_hd__and2_1
X_1700_ net272 net264 matmult_inst.mem_inst.mem3\[16\] VGND VGND VPWR VPWR _0587_
+ sky130_fd_sc_hd__and3_1
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1631_ matmult_inst.fsm_inst.state\[4\] matmult_inst.fsm_inst.state\[1\] _0537_ VGND
+ VGND VPWR VPWR _0550_ sky130_fd_sc_hd__or3_1
X_3301_ clknet_leaf_8_hz100 _0171_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB3\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3232_ clknet_leaf_7_hz100 net537 VGND VGND VPWR VPWR matmult_inst.fsm_inst.alu_result\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_3163_ net135 net124 VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__and2_1
X_2114_ _0904_ _0913_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3094_ net502 net84 net23 VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__mux2_1
X_2045_ net239 net257 net256 net237 VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_80_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout28 _1591_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_4
XFILLER_62_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout39 _1585_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_4
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2947_ net438 net79 net40 VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__mux2_1
X_2878_ net204 net508 net93 VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__mux2_1
X_1829_ net281 matmult_inst.mem_inst.mem0\[4\] matmult_inst.mem_inst.matrixB0\[4\]
+ net285 VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__a22o_1
Xmax_cap150 _0799_ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_1
Xmax_cap172 _1046_ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2801_ matmult_inst.alu_inst.adder_inst.r1.fa3.b matmult_inst.alu_inst.adder_inst.r1.fa3.a
+ VGND VGND VPWR VPWR _1515_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_14_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2732_ _1433_ _1453_ _1457_ _1469_ _1454_ VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__a311o_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2663_ _1375_ _1406_ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__nor2_1
X_1614_ net2 VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__inv_2
X_2594_ _1302_ _1303_ net18 VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__a21o_1
Xfanout218 matmult_inst.alu_inst.a0_reg\[6\] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__clkbuf_2
Xfanout207 matmult_inst.alu_inst.b0_reg\[4\] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__buf_2
Xfanout229 matmult_inst.alu_inst.a0_reg\[0\] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__buf_2
X_3215_ net290 VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__inv_2
X_3146_ net130 net118 VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__and2_1
XFILLER_27_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3077_ net430 _0809_ net26 VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__mux2_1
XFILLER_54_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2028_ _0825_ _0831_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__and2_1
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold261 matmult_inst.mem_inst.mem1\[14\] VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold250 matmult_inst.alu_inst.row1\[7\] VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 matmult_inst.alu_inst.row0\[2\] VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 matmult_inst.alu_inst.col1\[7\] VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 _0160_ VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3000_ net431 _0808_ net33 VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__mux2_1
XFILLER_36_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2715_ _1433_ _1457_ VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__nand2_1
X_2646_ net205 net207 net219 net217 VGND VGND VPWR VPWR _1391_ sky130_fd_sc_hd__and4_1
X_2577_ _1291_ _1292_ _1290_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__a21bo_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3129_ net130 net118 VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_53_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2500_ net212 net221 net220 net213 VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__a22o_1
X_3480_ clknet_leaf_21_hz100 _0340_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem0\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_2431_ _1181_ _1182_ _1171_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__a21oi_1
X_2362_ net198 _0541_ net194 _0756_ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__o31ai_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2293_ _1086_ _1087_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__nor2_1
XFILLER_37_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_466 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2629_ net50 _1371_ _1372_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__a21bo_1
XFILLER_47_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap47 net48 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2980_ net407 net84 net35 VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__mux2_1
X_1931_ _0796_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_72_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1862_ net279 matmult_inst.mem_inst.mem0\[1\] matmult_inst.mem_inst.matrixB0\[1\]
+ net282 VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__a22o_1
X_3601_ clknet_leaf_10_hz100 _0461_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA3\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_1793_ net271 net263 matmult_inst.mem_inst.mem3\[7\] VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__and3_1
X_3532_ clknet_leaf_20_hz100 _0392_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem3\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_3463_ clknet_leaf_29_hz100 _0323_ VGND VGND VPWR VPWR matmult_inst.alu_inst.b0_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2414_ net228 net226 net214 net215 VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__and4_1
X_3394_ clknet_leaf_4_hz100 _0256_ VGND VGND VPWR VPWR matmult_inst.alu_inst.col1\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2345_ _1131_ _1132_ _1134_ _1135_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__a31oi_1
X_2276_ net246 net234 net245 net236 VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__a22o_1
XFILLER_25_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2130_ _0927_ _0928_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__nand2_1
X_2061_ _0859_ _0860_ _0862_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_49_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2963_ net359 net82 net38 VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__mux2_1
X_1914_ matmult_inst.fsm_inst.count\[0\] _0544_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_32_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2894_ matmult_inst.fsm_inst.count\[2\] _0542_ VGND VGND VPWR VPWR _1579_ sky130_fd_sc_hd__or2_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1845_ net194 _0714_ _0716_ net279 VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__a22o_1
X_1776_ matmult_inst.mem_inst.matrixB2\[9\] net191 net183 matmult_inst.mem_inst.matrixB1\[9\]
+ _0655_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__a221o_1
X_3515_ clknet_leaf_23_hz100 _0375_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem2\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_3446_ clknet_leaf_1_hz100 _0306_ VGND VGND VPWR VPWR matmult_inst.alu_inst.out\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_3377_ clknet_leaf_2_hz100 _0240_ VGND VGND VPWR VPWR matmult_inst.alu_inst.row1\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2328_ _1096_ _1120_ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__xnor2_1
X_2259_ _1044_ _1051_ _1052_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__or3_1
XFILLER_72_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1630_ matmult_inst.fsm_inst.state\[1\] matmult_inst.fsm_inst.state\[0\] VGND VGND
+ VPWR VPWR _0549_ sky130_fd_sc_hd__nand2b_1
X_3300_ clknet_leaf_25_hz100 _0170_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB3\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3231_ clknet_leaf_7_hz100 net347 VGND VGND VPWR VPWR matmult_inst.fsm_inst.alu_result\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3162_ net135 net124 VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__and2_1
XFILLER_39_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2113_ _0911_ _0912_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__and2b_1
X_3093_ net462 _0806_ net23 VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__mux2_1
XFILLER_81_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2044_ net255 net237 VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__and2_1
XFILLER_81_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout29 _1590_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_4
X_2946_ net394 net80 net40 VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__mux2_1
X_2877_ net206 net437 net93 VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__mux2_1
X_1828_ matmult_inst.mem_inst.mem2\[4\] net190 net182 matmult_inst.mem_inst.mem1\[4\]
+ _0702_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__a221o_1
Xmax_cap151 _0790_ VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_1
X_1759_ net629 net91 _0640_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__o21a_1
Xmax_cap173 _0877_ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__buf_1
XFILLER_77_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3429_ clknet_leaf_4_hz100 _0289_ VGND VGND VPWR VPWR matmult_inst.alu_inst.b1_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2800_ net346 _1514_ net163 VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2731_ net634 _1472_ net160 VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__mux2_1
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2662_ _1375_ _1406_ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__and2_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1613_ net625 VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__inv_2
X_2593_ _1334_ _1335_ _1337_ _1279_ VGND VGND VPWR VPWR _1340_ sky130_fd_sc_hd__o211a_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout208 matmult_inst.alu_inst.b0_reg\[4\] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_2
Xfanout219 net220 VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__buf_2
X_3214_ net290 VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_19_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3145_ net131 net121 VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__and2_1
X_3076_ net501 net83 net26 VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__mux2_1
X_2027_ _0829_ _0830_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__nor2_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2929_ net559 net78 net42 VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__mux2_1
Xhold240 matmult_inst.mem_inst.mem2\[2\] VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 matmult_inst.mem_inst.mem2\[13\] VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 matmult_inst.mem_inst.matrixA2\[5\] VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 matmult_inst.mem_inst.matrixA1\[12\] VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 matmult_inst.mem_inst.matrixA2\[10\] VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 matmult_inst.mem_inst.matrixB0\[4\] VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2714_ _1407_ _1432_ _1435_ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__or3b_1
X_2645_ net205 net219 net217 net207 VGND VGND VPWR VPWR _1390_ sky130_fd_sc_hd__a22oi_2
XFILLER_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2576_ net227 net202 _1233_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__and3_1
XFILLER_55_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3128_ net129 net119 VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__and2_1
XFILLER_27_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3059_ net422 net81 net28 VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__mux2_1
XFILLER_42_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2430_ net229 net210 net211 net226 VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__a22o_1
X_2361_ _0564_ net166 _1148_ VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__and3_1
X_2292_ _1042_ _1062_ _1061_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__o21a_1
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2628_ _1371_ _1372_ net49 VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__a21o_1
X_2559_ net161 _1305_ _1306_ _1267_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__a31o_1
Xmax_cap59 net60 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_38_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1930_ matmult_inst.alu_inst.state\[0\] matmult_inst.alu_inst.state\[1\] VGND VGND
+ VPWR VPWR _0796_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_72_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1861_ matmult_inst.mem_inst.matrixA2\[1\] net186 net178 matmult_inst.mem_inst.matrixA1\[1\]
+ _0732_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__a221o_1
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3600_ clknet_leaf_16_hz100 _0460_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA3\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3531_ clknet_leaf_12_hz100 _0391_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem3\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_1792_ net617 net91 _0670_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__o21a_1
X_3462_ clknet_leaf_29_hz100 _0322_ VGND VGND VPWR VPWR matmult_inst.alu_inst.b0_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_2413_ net228 net214 net215 net226 VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__a22o_1
X_3393_ clknet_leaf_2_hz100 _0255_ VGND VGND VPWR VPWR matmult_inst.alu_inst.col1\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_2344_ net627 net159 VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__nor2_1
X_2275_ net246 net236 net234 net245 VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__and4_1
XFILLER_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2060_ _0840_ _0861_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__nor2_1
XFILLER_19_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2962_ net382 net83 net38 VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__mux2_1
X_1913_ _0781_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_32_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2893_ _1571_ _1577_ VGND VGND VPWR VPWR _1578_ sky130_fd_sc_hd__nor2_1
X_1844_ matmult_inst.mem_inst.matrixB2\[3\] net187 net179 matmult_inst.mem_inst.matrixB1\[3\]
+ _0717_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__a221o_1
X_1775_ net273 net265 matmult_inst.mem_inst.matrixB3\[9\] VGND VGND VPWR VPWR _0655_
+ sky130_fd_sc_hd__and3_1
X_3514_ clknet_leaf_20_hz100 _0374_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem2\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_3445_ clknet_leaf_26_hz100 _0305_ VGND VGND VPWR VPWR matmult_inst.alu_inst.out\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_3376_ clknet_leaf_4_hz100 _0239_ VGND VGND VPWR VPWR matmult_inst.alu_inst.row1\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_2327_ _1117_ _1118_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__xnor2_1
X_2258_ _1051_ _1052_ _1044_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__o21ai_1
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2189_ _0984_ _0985_ _0986_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__a21o_1
XFILLER_80_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3230_ clknet_leaf_6_hz100 _0128_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.alu_result\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3161_ net136 net125 VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__and2_1
XFILLER_39_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2112_ _0909_ _0910_ _0877_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__a21o_1
X_3092_ net519 net86 net23 VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__mux2_1
XFILLER_81_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2043_ _0844_ _0845_ net649 net175 VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_45_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2945_ net405 net81 net39 VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__mux2_1
X_2876_ net208 net590 net94 VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__mux2_1
X_1827_ net271 net263 matmult_inst.mem_inst.mem3\[4\] VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__and3_1
Xmax_cap152 net153 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__buf_1
Xmax_cap141 _1254_ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_1
X_1758_ net283 _0634_ _0639_ _0632_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__a211o_1
X_1689_ net272 net264 matmult_inst.mem_inst.mem3\[17\] VGND VGND VPWR VPWR _0577_
+ sky130_fd_sc_hd__and3_1
X_3428_ clknet_leaf_2_hz100 _0288_ VGND VGND VPWR VPWR matmult_inst.alu_inst.b1_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3359_ clknet_leaf_24_hz100 _0223_ VGND VGND VPWR VPWR matmult_inst.addr\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_13_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2730_ _1470_ _1471_ VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__xnor2_1
X_2661_ _1386_ _1405_ VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__xnor2_1
X_1612_ net277 VGND VGND VPWR VPWR _1606_ sky130_fd_sc_hd__inv_2
X_2592_ _1338_ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__inv_2
Xfanout209 matmult_inst.alu_inst.b0_reg\[3\] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_4
XFILLER_67_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3213_ net290 VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__inv_2
X_3144_ net132 net121 VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__and2_1
XFILLER_39_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3075_ net459 net84 net25 VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__mux2_1
X_2026_ net258 net241 _0827_ _0828_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2928_ net432 net79 net42 VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__mux2_1
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2859_ _1562_ _1563_ VGND VGND VPWR VPWR _1564_ sky130_fd_sc_hd__xnor2_1
Xhold241 matmult_inst.mem_inst.matrixA2\[11\] VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 matmult_inst.mem_inst.matrixA2\[3\] VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 matmult_inst.mem_inst.matrixB1\[13\] VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 matmult_inst.alu_inst.col0\[4\] VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 matmult_inst.mem_inst.matrixB0\[0\] VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 matmult_inst.alu_inst.col1\[3\] VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 matmult_inst.mem_inst.matrixB0\[8\] VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2713_ _1453_ _1455_ VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__nand2_1
X_2644_ net212 net216 _1357_ _1358_ net219 VGND VGND VPWR VPWR _1389_ sky130_fd_sc_hd__a32oi_2
X_2575_ _1315_ _1321_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__xnor2_1
X_3127_ net130 net118 VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__and2_1
XFILLER_35_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3058_ net464 net82 net28 VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__mux2_1
X_2009_ matmult_inst.fsm_inst.alu_result\[15\] net114 VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_53_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0__f_hz100 clknet_0_hz100 VGND VGND VPWR VPWR clknet_2_0__leaf_hz100 sky130_fd_sc_hd__clkbuf_16
XFILLER_23_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_47_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2360_ net260 _0783_ _0784_ net200 VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__o22a_1
X_2291_ _1082_ _1085_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_56_Left_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_65_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2627_ net49 _1371_ _1372_ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__nand3_1
X_2558_ _1301_ net18 _1303_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__o21ai_1
X_2489_ _1222_ _1234_ _1235_ _1236_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__nand4_1
XPHY_EDGE_ROW_74_Left_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap49 net50 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_38_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1860_ net267 net260 matmult_inst.mem_inst.matrixA3\[1\] VGND VGND VPWR VPWR _0732_
+ sky130_fd_sc_hd__and3_1
X_1791_ net285 _0664_ _0669_ _0662_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__a211o_1
X_3530_ clknet_leaf_13_hz100 _0390_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem3\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3461_ clknet_leaf_29_hz100 _0321_ VGND VGND VPWR VPWR matmult_inst.alu_inst.b0_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_2412_ net646 net175 _1166_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__a21o_1
XFILLER_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3392_ clknet_leaf_2_hz100 _0254_ VGND VGND VPWR VPWR matmult_inst.alu_inst.col1\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_2343_ net159 _1116_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__and2_1
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2274_ net234 net245 VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__and2_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1989_ matmult_inst.fsm_inst.rx_data\[5\] _0786_ net113 matmult_inst.fsm_inst.alu_result\[5\]
+ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__a22o_1
XFILLER_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3659_ clknet_leaf_23_hz100 _0519_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB2\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2961_ net323 _0807_ net37 VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__mux2_1
X_1912_ matmult_inst.alu_inst.complete _0779_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_32_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2892_ matmult_inst.fsm_inst.count\[2\] _0542_ VGND VGND VPWR VPWR _1577_ sky130_fd_sc_hd__nand2_1
XFILLER_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1843_ net267 net260 matmult_inst.mem_inst.matrixB3\[3\] VGND VGND VPWR VPWR _0717_
+ sky130_fd_sc_hd__and3_1
X_1774_ matmult_inst.mem_inst.matrixA2\[9\] net191 net183 matmult_inst.mem_inst.matrixA1\[9\]
+ _0653_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__a221o_1
X_3513_ clknet_leaf_12_hz100 _0373_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem2\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_3444_ clknet_leaf_1_hz100 _0304_ VGND VGND VPWR VPWR matmult_inst.alu_inst.out\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_3375_ clknet_leaf_4_hz100 _0238_ VGND VGND VPWR VPWR matmult_inst.alu_inst.row1\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_2326_ _1117_ _1118_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__nor2_1
XFILLER_69_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2257_ _1045_ _1049_ _1050_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_48_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2188_ net242 net245 VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__nand2_1
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3160_ net134 net123 VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__and2_1
X_3091_ net540 _0804_ net23 VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__mux2_1
X_2111_ _0877_ _0909_ _0910_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__and3_1
Xhold1 matmult_inst.spi_inst.cs_sync VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__dlygate4sd3_1
X_2042_ _0829_ _0832_ _0843_ net162 VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__o31ai_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2944_ net515 net82 net40 VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__mux2_1
X_2875_ net210 net489 net93 VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__mux2_1
X_1826_ net621 _0701_ net91 VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__mux2_1
X_1757_ net287 _0636_ _0638_ net278 VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__a22o_1
Xmax_cap142 _1216_ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_1
X_1688_ matmult_inst.mem_inst.matrixA2\[17\] net192 net184 matmult_inst.mem_inst.matrixA1\[17\]
+ _0575_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__a221o_1
Xmax_cap197 _0543_ VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3427_ clknet_leaf_2_hz100 _0287_ VGND VGND VPWR VPWR matmult_inst.alu_inst.b1_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3358_ clknet_leaf_8_hz100 net296 VGND VGND VPWR VPWR matmult_inst.fsm_inst.rx_valid_delay
+ sky130_fd_sc_hd__dfxtp_1
X_2309_ net248 net230 net233 net246 VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__a22o_1
X_3289_ clknet_leaf_9_hz100 net469 _0070_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.rx_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2660_ _1402_ _1403_ VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__xor2_1
X_1611_ matmult_inst.fsm_inst.count\[3\] VGND VGND VPWR VPWR _1605_ sky130_fd_sc_hd__inv_2
XFILLER_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2591_ _1279_ _1337_ _1335_ net20 VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__a211oi_1
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3212_ net289 VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__inv_2
X_3143_ net134 net123 VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__and2_1
X_3074_ net496 _0806_ net25 VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__mux2_1
X_2025_ _0827_ _0828_ net258 net241 VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__and4bb_1
XFILLER_50_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2927_ net397 net80 net42 VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__mux2_1
X_2858_ _1557_ net7 _1558_ VGND VGND VPWR VPWR _1563_ sky130_fd_sc_hd__o21ai_2
Xhold220 matmult_inst.mem_inst.matrixA2\[15\] VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__dlygate4sd3_1
X_1809_ net272 net264 matmult_inst.mem_inst.matrixB3\[6\] VGND VGND VPWR VPWR _0686_
+ sky130_fd_sc_hd__and3_1
X_2789_ matmult_inst.alu_inst.adder_inst.r1.fa1.b matmult_inst.alu_inst.adder_inst.r1.fa1.a
+ VGND VGND VPWR VPWR _1505_ sky130_fd_sc_hd__or2_1
Xhold231 matmult_inst.alu_inst.adder_inst.r2.fa1.b VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 matmult_inst.alu_inst.col1\[1\] VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 matmult_inst.fsm_inst.alu_result\[7\] VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 matmult_inst.mem_inst.mem0\[14\] VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 matmult_inst.alu_inst.out\[0\] VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold286 matmult_inst.alu_inst.out\[8\] VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 matmult_inst.mem_inst.mem1\[11\] VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_56_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2712_ net12 VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__inv_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2643_ net221 net203 VGND VGND VPWR VPWR _1388_ sky130_fd_sc_hd__and2_1
X_2574_ _1319_ _1320_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__or2_1
X_3126_ net134 net123 VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__and2_1
XFILLER_55_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3057_ net578 net83 net28 VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__mux2_1
X_2008_ net310 net73 net55 VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__mux2_1
XFILLER_35_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2290_ _1083_ _1084_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__or2_1
XFILLER_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2626_ _1326_ _1362_ _1370_ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__nand3_1
X_2557_ _1301_ _1303_ net18 VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__or3_1
X_2488_ _1234_ _1235_ _1236_ _1222_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__a22o_1
XFILLER_28_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap17 _1338_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3109_ matmult_inst.fsm_inst.tx_start_send _0554_ _0781_ _1569_ VGND VGND VPWR VPWR
+ _1594_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_66_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1790_ matmult_inst.fsm_inst.sel\[0\] _0666_ _0668_ net280 VGND VGND VPWR VPWR _0669_
+ sky130_fd_sc_hd__a22o_1
X_3460_ clknet_leaf_29_hz100 _0320_ VGND VGND VPWR VPWR matmult_inst.alu_inst.b0_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_2411_ net228 net215 net161 VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__and3_1
X_3391_ clknet_leaf_2_hz100 _0253_ VGND VGND VPWR VPWR matmult_inst.alu_inst.col1\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2342_ _1131_ _1132_ _1133_ net174 net614 VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__a32o_1
X_2273_ net619 _1068_ net159 VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__mux2_1
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1988_ net340 net83 net56 VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__mux2_1
X_3658_ clknet_leaf_21_hz100 _0518_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB2\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_2609_ _1353_ _1354_ VGND VGND VPWR VPWR _1355_ sky130_fd_sc_hd__nor2_1
X_3589_ clknet_leaf_18_hz100 _0449_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA2\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout190 net192 VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2960_ net344 net85 net37 VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__mux2_1
X_2891_ _1576_ matmult_inst.fsm_inst.count\[1\] _1571_ VGND VGND VPWR VPWR _0325_
+ sky130_fd_sc_hd__mux2_1
X_1911_ _0779_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_32_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1842_ matmult_inst.mem_inst.mem2\[3\] net187 net179 matmult_inst.mem_inst.mem1\[3\]
+ _0715_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__a221o_1
XFILLER_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1773_ net273 net265 matmult_inst.mem_inst.matrixA3\[9\] VGND VGND VPWR VPWR _0653_
+ sky130_fd_sc_hd__and3_1
X_3512_ clknet_leaf_13_hz100 _0372_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem2\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3443_ clknet_leaf_26_hz100 _0303_ VGND VGND VPWR VPWR matmult_inst.alu_inst.out\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_3374_ clknet_leaf_2_hz100 _0237_ VGND VGND VPWR VPWR matmult_inst.alu_inst.row1\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_2325_ _1069_ _1105_ _1103_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__o21ai_1
X_2256_ _1045_ _1049_ _1050_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__and3_1
XFILLER_69_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2187_ net238 net240 net249 net247 VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__nand4_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2110_ _0905_ _0907_ _0908_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__or3b_1
X_3090_ net282 net186 _0802_ VGND VGND VPWR VPWR _1593_ sky130_fd_sc_hd__and3_1
Xhold2 matmult_inst.fsm_inst.rx_valid VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2041_ _0829_ _0832_ _0843_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_45_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2943_ net465 net83 net40 VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__mux2_1
X_2874_ net211 net595 net94 VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__mux2_1
X_1825_ _0695_ _0698_ _0700_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__or3_1
X_1756_ matmult_inst.mem_inst.mem2\[11\] net186 net178 matmult_inst.mem_inst.mem1\[11\]
+ _0637_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__a221o_1
Xmax_cap165 _0774_ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__buf_1
Xmax_cap154 _0552_ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dlymetal6s2s_1
X_1687_ net272 net264 matmult_inst.mem_inst.matrixA3\[17\] VGND VGND VPWR VPWR _0575_
+ sky130_fd_sc_hd__and3_1
X_3426_ clknet_leaf_2_hz100 _0286_ VGND VGND VPWR VPWR matmult_inst.alu_inst.b1_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3357_ clknet_leaf_1_hz100 _0222_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.fa.b
+ sky130_fd_sc_hd__dfxtp_1
X_2308_ net246 net233 VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__nand2_1
X_3288_ clknet_leaf_11_hz100 net298 _0069_ VGND VGND VPWR VPWR matmult_inst.spi_inst.rx_done2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2239_ _0998_ _1034_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__nand2_1
XFILLER_38_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1610_ matmult_inst.fsm_inst.count\[0\] VGND VGND VPWR VPWR _1604_ sky130_fd_sc_hd__inv_2
XFILLER_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2590_ _1280_ _1296_ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__nand2_1
X_3211_ net289 VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__inv_2
X_3142_ net129 net118 VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__and2_1
XFILLER_79_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3073_ net574 net86 net25 VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__mux2_1
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2024_ net256 net243 net254 net244 VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__and4_1
XFILLER_62_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2926_ net610 net81 net41 VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__mux2_1
X_2857_ matmult_inst.alu_inst.adder_inst.fa.b matmult_inst.alu_inst.adder_inst.fa.a
+ VGND VGND VPWR VPWR _1562_ sky130_fd_sc_hd__xnor2_1
X_1808_ matmult_inst.mem_inst.matrixA2\[6\] net189 net181 matmult_inst.mem_inst.matrixA1\[6\]
+ _0684_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__a221o_1
Xhold210 matmult_inst.mem_inst.mem1\[10\] VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__dlygate4sd3_1
X_2788_ matmult_inst.alu_inst.adder_inst.r1.fa1.b matmult_inst.alu_inst.adder_inst.r1.fa1.a
+ VGND VGND VPWR VPWR _1504_ sky130_fd_sc_hd__nor2_1
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1739_ matmult_inst.mem_inst.matrixA0\[12\] net168 _0621_ net195 net115 VGND VGND
+ VPWR VPWR _0622_ sky130_fd_sc_hd__a221o_1
Xhold232 matmult_inst.mem_inst.matrixA0\[16\] VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 matmult_inst.mem_inst.mem2\[5\] VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 _0130_ VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 matmult_inst.mem_inst.matrixB0\[13\] VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 matmult_inst.alu_inst.out\[4\] VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 _0131_ VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 matmult_inst.mem_inst.mem1\[9\] VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__dlygate4sd3_1
X_3409_ clknet_leaf_31_hz100 _0270_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r3.fa1.a
+ sky130_fd_sc_hd__dfxtp_1
Xhold298 matmult_inst.spi_inst.mosi_data_sync\[3\] VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2711_ net16 _1452_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__nor2_1
X_2642_ _1352_ _1360_ _1354_ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__a21o_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2573_ _1316_ _1317_ _1318_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__a21oi_1
X_3125_ net131 net120 VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__and2_1
X_3056_ net517 net84 net27 VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__mux2_1
X_2007_ matmult_inst.fsm_inst.alu_result\[14\] net114 VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_53_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2909_ net494 net79 net44 VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__mux2_1
XFILLER_76_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2625_ _1326_ _1362_ _1370_ VGND VGND VPWR VPWR _1371_ sky130_fd_sc_hd__a21o_1
X_2556_ _1297_ _1298_ _1300_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__a21oi_1
X_2487_ net205 net229 _1220_ net171 _1190_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__a41o_1
Xmax_cap18 _1304_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_1
X_3108_ net458 net70 net24 VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3039_ net328 net82 net30 VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2410_ _1160_ net577 net63 VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__mux2_1
X_3390_ clknet_leaf_2_hz100 _0252_ VGND VGND VPWR VPWR matmult_inst.alu_inst.col1\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2341_ _1123_ _1127_ _1130_ net159 VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__o31a_1
X_2272_ _1035_ _1067_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__xnor2_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1987_ matmult_inst.fsm_inst.rx_data\[4\] _0786_ net113 matmult_inst.fsm_inst.alu_result\[4\]
+ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__a22o_1
X_3657_ clknet_leaf_12_hz100 _0517_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB2\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_3588_ clknet_leaf_22_hz100 _0448_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA2\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_2608_ _1345_ _1350_ _1351_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__and3_1
X_2539_ _1285_ _1286_ _1281_ VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__a21oi_1
XFILLER_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire60 _1322_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
XFILLER_24_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout180 net185 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_4
Xfanout191 net192 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_4
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2890_ net166 _1575_ _0787_ VGND VGND VPWR VPWR _1576_ sky130_fd_sc_hd__o21a_1
X_1910_ _0549_ _0778_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__or2_1
XFILLER_30_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1841_ net270 net260 matmult_inst.mem_inst.mem3\[3\] VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__and3_1
XFILLER_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1772_ matmult_inst.mem_inst.matrixA0\[9\] net169 _0651_ net196 net115 VGND VGND
+ VPWR VPWR _0652_ sky130_fd_sc_hd__a221o_1
X_3511_ clknet_leaf_13_hz100 _0371_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem2\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_3442_ clknet_leaf_26_hz100 _0302_ VGND VGND VPWR VPWR matmult_inst.alu_inst.out\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_3373_ clknet_leaf_4_hz100 _0236_ VGND VGND VPWR VPWR matmult_inst.alu_inst.row1\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2324_ _1115_ _1116_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__nand2_1
X_2255_ _1049_ _1050_ _1045_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__a21oi_1
X_2186_ net238 net249 net247 net240 VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__a22o_1
XFILLER_25_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3 matmult_inst.fsm_inst.tx_ready_delay VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__dlygate4sd3_1
X_2040_ _0836_ _0842_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__xnor2_1
X_2942_ net564 _0807_ net39 VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__mux2_1
X_2873_ net214 net367 net94 VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__mux2_1
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1824_ matmult_inst.mem_inst.matrixA0\[5\] net169 _0699_ net195 VGND VGND VPWR VPWR
+ _0700_ sky130_fd_sc_hd__a22o_1
X_1755_ net268 net261 matmult_inst.mem_inst.mem3\[11\] VGND VGND VPWR VPWR _0637_
+ sky130_fd_sc_hd__and3_1
Xmax_cap144 _1016_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_1
Xmax_cap177 _0770_ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__buf_1
Xmax_cap155 _0548_ VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__buf_1
X_1686_ matmult_inst.mem_inst.matrixB2\[17\] net191 net183 matmult_inst.mem_inst.matrixB1\[17\]
+ _0573_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__a221o_1
X_3425_ clknet_leaf_6_hz100 _0285_ VGND VGND VPWR VPWR matmult_inst.alu_inst.b1_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3356_ clknet_leaf_3_hz100 _0221_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r3.fa3.b
+ sky130_fd_sc_hd__dfxtp_1
X_2307_ _1099_ _1100_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__nand2b_1
X_3287_ clknet_leaf_10_hz100 matmult_inst.spi_inst.next_state _0068_ VGND VGND VPWR
+ VPWR matmult_inst.spi_inst.current_state sky130_fd_sc_hd__dfrtp_4
X_2238_ _0996_ _0997_ _1033_ _1034_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__a31o_1
XFILLER_72_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2169_ _0965_ _0966_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_0_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3210_ net289 VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__inv_2
XFILLER_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3141_ net129 net119 VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__and2_1
XFILLER_67_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3072_ net455 _0804_ net25 VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__mux2_1
X_2023_ net256 net242 net254 net244 VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__a22oi_1
X_2925_ net573 net82 net42 VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_17_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2856_ net450 net6 net164 VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1807_ net271 net263 matmult_inst.mem_inst.matrixA3\[6\] VGND VGND VPWR VPWR _0684_
+ sky130_fd_sc_hd__and3_1
X_2787_ matmult_inst.alu_inst.adder_inst.r1.fa1.b matmult_inst.alu_inst.adder_inst.r1.fa1.a
+ VGND VGND VPWR VPWR _1503_ sky130_fd_sc_hd__nand2_1
Xhold200 matmult_inst.mem_inst.mem0\[8\] VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 matmult_inst.mem_inst.matrixA1\[8\] VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 matmult_inst.alu_inst.row0\[7\] VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 matmult_inst.mem_inst.matrixB1\[11\] VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__dlygate4sd3_1
X_1738_ net278 matmult_inst.mem_inst.mem0\[12\] matmult_inst.mem_inst.matrixB0\[12\]
+ net283 VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__a22o_1
Xhold244 matmult_inst.mem_inst.matrixA2\[6\] VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 matmult_inst.mem_inst.mem2\[12\] VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 matmult_inst.mem_inst.mem0\[0\] VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__dlygate4sd3_1
X_1669_ matmult_inst.fsm_inst.rx_data\[5\] net571 matmult_inst.spi_inst.rx_done_sys
+ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__mux2_1
Xhold277 matmult_inst.spi_inst.mosi_data_sync\[5\] VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__dlygate4sd3_1
X_3408_ clknet_leaf_31_hz100 _0269_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r3.fa0.a
+ sky130_fd_sc_hd__dfxtp_1
Xhold299 _0162_ VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 matmult_inst.spi_inst.mosi_data_sync\[7\] VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__dlygate4sd3_1
X_3339_ clknet_leaf_24_hz100 net92 VGND VGND VPWR VPWR matmult_inst.fsm_inst.load_delay
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2710_ net16 _1452_ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__nand2_1
XFILLER_71_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2641_ _1383_ _1385_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_10_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2572_ _1316_ _1317_ _1318_ VGND VGND VPWR VPWR _1319_ sky130_fd_sc_hd__and3_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3124_ net134 net123 VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__and2_1
X_3055_ net518 net85 net27 VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__mux2_1
X_2006_ net348 net74 net55 VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2908_ net483 net80 net44 VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2839_ matmult_inst.alu_inst.adder_inst.r3.fa1.b matmult_inst.alu_inst.adder_inst.r3.fa1.a
+ VGND VGND VPWR VPWR _1547_ sky130_fd_sc_hd__nor2_1
XFILLER_76_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_25_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2624_ _1367_ _1369_ VGND VGND VPWR VPWR _1370_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_34_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2555_ _1227_ _1261_ _1263_ _1260_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__o31a_1
X_2486_ net205 net227 net204 net229 VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__a22o_1
X_3107_ net373 net71 net24 VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__mux2_1
XFILLER_43_419 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3038_ net317 net83 net29 VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__mux2_1
XFILLER_70_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_52_Left_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_70_Left_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2340_ _1123_ _1127_ _1130_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__o21ai_1
X_2271_ _1065_ _1066_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__nand2b_1
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1986_ net352 net84 net55 VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__mux2_1
X_3656_ clknet_leaf_10_hz100 _0516_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB2\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3587_ clknet_leaf_22_hz100 _0447_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA2\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_2607_ _1352_ VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__inv_2
X_2538_ net170 _1283_ _1284_ VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__o21ai_1
X_2469_ _1193_ _1217_ _1218_ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__a21o_1
XFILLER_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire50 _1361_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_5_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout181 net184 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_4
Xfanout192 net193 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1840_ net279 matmult_inst.mem_inst.mem0\[3\] matmult_inst.mem_inst.matrixB0\[3\]
+ net282 VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__a22o_1
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3510_ clknet_leaf_15_hz100 _0370_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem2\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_1771_ net280 matmult_inst.mem_inst.mem0\[9\] matmult_inst.mem_inst.matrixB0\[9\]
+ net286 VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__a22o_1
X_3441_ clknet_leaf_26_hz100 _0301_ VGND VGND VPWR VPWR matmult_inst.alu_inst.out\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3372_ clknet_leaf_6_hz100 _0235_ VGND VGND VPWR VPWR matmult_inst.alu_inst.row1\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2323_ net246 net230 net233 net245 VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__nand4_1
XFILLER_69_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2254_ net172 _1047_ _1048_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__o21ai_1
X_2185_ _0981_ _0982_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__nand2_1
XFILLER_25_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1969_ net476 net58 net21 matmult_inst.fsm_inst.alu_result\[11\] VGND VGND VPWR VPWR
+ _0134_ sky130_fd_sc_hd__a22o_1
XFILLER_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3639_ clknet_leaf_12_hz100 _0499_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB1\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold4 matmult_inst.spi_inst.rx_done1 VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2941_ net534 net85 net39 VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__mux2_1
X_2872_ net604 net600 net94 VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__mux2_1
X_1823_ net281 matmult_inst.mem_inst.mem0\[5\] matmult_inst.mem_inst.matrixB0\[5\]
+ net285 VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__a22o_1
X_1754_ matmult_inst.mem_inst.matrixA2\[11\] net186 net178 matmult_inst.mem_inst.matrixA1\[11\]
+ _0635_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__a221o_1
Xmax_cap101 net102 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
Xmax_cap112 _0881_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_1
Xmax_cap145 _0967_ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_1
X_1685_ net272 net264 matmult_inst.mem_inst.matrixB3\[17\] VGND VGND VPWR VPWR _0573_
+ sky130_fd_sc_hd__and3_1
X_3424_ clknet_leaf_5_hz100 _0284_ VGND VGND VPWR VPWR matmult_inst.alu_inst.b1_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3355_ clknet_leaf_3_hz100 _0220_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r3.fa2.b
+ sky130_fd_sc_hd__dfxtp_1
X_3286_ net293 _0013_ _0067_ VGND VGND VPWR VPWR matmult_inst.spi_inst.miso_shifter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_2306_ _1076_ _1098_ _1097_ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__a21o_1
X_2237_ _0974_ _1031_ _1032_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__and3_1
XFILLER_53_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2168_ _0949_ _0951_ _0948_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__o21ai_1
XFILLER_80_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2099_ _0896_ _0897_ _0868_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__a21o_1
XFILLER_80_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_3__f_hz100 clknet_0_hz100 VGND VGND VPWR VPWR clknet_2_3__leaf_hz100 sky130_fd_sc_hd__clkbuf_16
XFILLER_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3140_ net129 net119 VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_8_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3071_ net282 net178 _0802_ VGND VGND VPWR VPWR _1592_ sky130_fd_sc_hd__and3_1
XFILLER_67_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2022_ net650 net175 _0824_ _0826_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2924_ net398 net83 net42 VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__mux2_1
X_2855_ _1559_ _1560_ VGND VGND VPWR VPWR _1561_ sky130_fd_sc_hd__xnor2_1
X_1806_ net281 matmult_inst.mem_inst.mem0\[6\] matmult_inst.mem_inst.matrixB0\[6\]
+ net286 VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__a22o_1
X_2786_ net570 _1502_ net163 VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__mux2_1
Xhold201 matmult_inst.mem_inst.matrixB2\[4\] VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 matmult_inst.mem_inst.matrixB0\[3\] VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__dlygate4sd3_1
X_1737_ net642 net92 _0612_ _0620_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__o22a_1
Xhold234 matmult_inst.mem_inst.matrixA1\[13\] VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 matmult_inst.alu_inst.adder_inst.r2.fa3.b VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 matmult_inst.mem_inst.matrixA0\[10\] VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 matmult_inst.mem_inst.mem0\[5\] VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 matmult_inst.fsm_inst.alu_result\[5\] VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold278 _0164_ VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__dlygate4sd3_1
X_1668_ matmult_inst.fsm_inst.rx_data\[6\] net335 matmult_inst.spi_inst.rx_done_sys
+ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__mux2_1
X_3407_ clknet_leaf_31_hz100 _0268_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r2.fa3.a
+ sky130_fd_sc_hd__dfxtp_1
Xhold289 _0166_ VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__dlygate4sd3_1
X_3338_ _0121_ _0205_ _0120_ VGND VGND VPWR VPWR matmult_inst.spi_inst.rx_bit_count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3269_ clknet_leaf_12_hz100 _0158_ _0050_ VGND VGND VPWR VPWR matmult_inst.spi_inst.tx_reg_sys\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2640_ net222 net202 _1384_ VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_10_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2571_ net213 matmult_inst.alu_inst.a0_reg\[7\] VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__nand2_1
X_3123_ matmult_inst.fsm_inst.state\[0\] _0778_ _1137_ _1595_ _0550_ VGND VGND VPWR
+ VPWR _0532_ sky130_fd_sc_hd__o2111ai_1
X_3054_ net511 net86 net27 VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__mux2_1
X_2005_ matmult_inst.fsm_inst.alu_result\[13\] net114 VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_53_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2907_ net443 _0810_ net44 VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2838_ net342 net11 net164 VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__mux2_1
X_2769_ _1486_ _1487_ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__and2b_1
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3672_ clknet_leaf_27_hz100 _0532_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.state\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2623_ net227 net201 _1368_ VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__and3_1
X_2554_ _1297_ _1298_ _1300_ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__nand3_1
X_2485_ net206 net229 net227 net204 VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__nand4_2
X_3106_ net562 _0819_ net23 VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__mux2_1
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3037_ net338 net84 net29 VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__mux2_1
XFILLER_70_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2270_ _1029_ _1064_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__or2_1
XFILLER_77_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1985_ matmult_inst.fsm_inst.rx_data\[3\] _0786_ net113 matmult_inst.fsm_inst.alu_result\[3\]
+ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__a22o_1
XFILLER_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3655_ clknet_leaf_10_hz100 _0515_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB2\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2606_ _1350_ _1351_ _1345_ VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__a21o_1
X_3586_ clknet_leaf_21_hz100 _0446_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA2\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_2537_ _1282_ _1283_ _1284_ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__or3_1
X_2468_ _1193_ _1216_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__nor2_1
XFILLER_57_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2399_ _1159_ net508 net65 VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__mux2_1
XFILLER_28_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire62 _1256_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_24_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout160 net161 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_2
Xfanout182 net184 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout193 _0571_ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1770_ net638 net92 _0650_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__o21a_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3440_ clknet_leaf_26_hz100 _0300_ VGND VGND VPWR VPWR matmult_inst.alu_inst.out\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_3371_ clknet_leaf_2_hz100 _0234_ VGND VGND VPWR VPWR matmult_inst.alu_inst.row1\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2322_ net246 net230 net233 net245 VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__a22o_1
XFILLER_69_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2253_ _1046_ _1047_ _1048_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__or3_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2184_ net158 _0979_ _0980_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_48_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1968_ net466 net58 net21 matmult_inst.fsm_inst.alu_result\[10\] VGND VGND VPWR VPWR
+ _0133_ sky130_fd_sc_hd__a22o_1
X_1899_ _0755_ _0758_ _0764_ net153 VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__nor4_1
X_3638_ clknet_leaf_10_hz100 _0498_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB1\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3569_ clknet_leaf_23_hz100 _0429_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA1\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold5 matmult_inst.fsm_inst.rx_ready_edge VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_81_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2940_ net478 net86 net39 VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__mux2_1
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2871_ net216 net527 net93 VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__mux2_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1822_ net195 _0697_ net288 VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__and3b_1
X_1753_ net268 net261 matmult_inst.mem_inst.matrixA3\[11\] VGND VGND VPWR VPWR _0635_
+ sky130_fd_sc_hd__and3_1
X_1684_ net261 net268 VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__and2b_1
Xmax_cap102 _0527_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__buf_1
Xmax_cap146 _0955_ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_1
Xmax_cap157 _1312_ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_1
X_3423_ clknet_leaf_6_hz100 _0283_ VGND VGND VPWR VPWR matmult_inst.alu_inst.b1_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3354_ clknet_leaf_31_hz100 _0219_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r3.fa1.b
+ sky130_fd_sc_hd__dfxtp_1
X_3285_ net293 _0012_ _0066_ VGND VGND VPWR VPWR matmult_inst.spi_inst.miso_shifter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_2305_ _1076_ _1097_ _1098_ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__and3_1
X_2236_ _0974_ _1032_ _1031_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__a21o_1
X_2167_ net255 net231 _0892_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_0_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2098_ _0868_ _0896_ _0897_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__nand3_1
XFILLER_80_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3070_ net357 net70 net28 VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__mux2_1
X_2021_ net175 _0825_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__nor2_1
XFILLER_35_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2923_ net599 net84 net41 VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__mux2_1
X_2854_ _1552_ _1555_ _1553_ VGND VGND VPWR VPWR _1560_ sky130_fd_sc_hd__a21boi_1
X_1805_ matmult_inst.mem_inst.mem2\[6\] net189 net181 matmult_inst.mem_inst.mem1\[6\]
+ _0681_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__a221o_1
X_2785_ _1499_ _1501_ VGND VGND VPWR VPWR _1502_ sky130_fd_sc_hd__xnor2_1
Xhold202 matmult_inst.mem_inst.matrixB1\[2\] VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__dlygate4sd3_1
X_1736_ net278 _0617_ _0619_ net283 _0615_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__a221o_1
Xhold235 matmult_inst.mem_inst.matrixB1\[15\] VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 matmult_inst.mem_inst.matrixB0\[2\] VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 matmult_inst.mem_inst.mem2\[16\] VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 matmult_inst.mem_inst.matrixB2\[15\] VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 matmult_inst.alu_inst.adder_inst.r2.fa2.a VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 matmult_inst.mem_inst.matrixB2\[0\] VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__dlygate4sd3_1
X_1667_ matmult_inst.fsm_inst.rx_data\[7\] net582 matmult_inst.spi_inst.rx_done_sys
+ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__mux2_1
X_3406_ clknet_leaf_0_hz100 _0267_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r2.fa2.a
+ sky130_fd_sc_hd__dfxtp_1
Xhold279 matmult_inst.mem_inst.mem1\[5\] VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3337_ _0119_ _0204_ _0118_ VGND VGND VPWR VPWR matmult_inst.spi_inst.rx_bit_count\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_3268_ clknet_leaf_14_hz100 _0157_ _0049_ VGND VGND VPWR VPWR matmult_inst.spi_inst.tx_reg_sys\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3199_ net289 VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__inv_2
X_2219_ _1012_ _1015_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2570_ net209 net212 net219 net218 VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__nand4_1
X_3122_ _0548_ _1596_ _1603_ _0781_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__o31a_1
XFILLER_67_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3053_ net568 net87 net27 VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__mux2_1
X_2004_ net318 _0816_ net55 VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__mux2_1
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2906_ net539 net82 net44 VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2837_ _1544_ _1545_ VGND VGND VPWR VPWR _1546_ sky130_fd_sc_hd__xnor2_1
X_2768_ matmult_inst.alu_inst.adder_inst.r0.fa2.b matmult_inst.alu_inst.adder_inst.r0.fa2.a
+ VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__nand2_1
X_2699_ _1420_ _1422_ _1419_ VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__a21o_1
X_1719_ matmult_inst.mem_inst.mem2\[14\] net193 net185 matmult_inst.mem_inst.mem1\[14\]
+ _0603_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_69_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3671_ clknet_leaf_27_hz100 _0531_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.state\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2622_ _1233_ _1324_ VGND VGND VPWR VPWR _1368_ sky130_fd_sc_hd__nand2_1
XFILLER_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2553_ _1297_ _1298_ _1300_ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__and3_1
X_2484_ net229 net204 VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__nand2_1
XFILLER_28_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3105_ net472 _0818_ net23 VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__mux2_1
X_3036_ net390 net85 net29 VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1984_ net314 net85 net55 VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3654_ clknet_leaf_18_hz100 _0514_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB2\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_2605_ _1346_ _1348_ _1349_ VGND VGND VPWR VPWR _1351_ sky130_fd_sc_hd__or3_1
X_3585_ clknet_leaf_12_hz100 _0445_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA2\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_2536_ net209 matmult_inst.alu_inst.a0_reg\[4\] VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__and2_1
X_2467_ _1191_ net142 VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__xnor2_1
X_2398_ _1158_ net437 net65 VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__mux2_1
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3019_ net372 _0808_ net31 VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__mux2_1
XFILLER_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout161 net162 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_4
Xfanout183 net184 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_4
Xfanout194 net195 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__buf_2
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3370_ clknet_leaf_2_hz100 _0233_ VGND VGND VPWR VPWR matmult_inst.alu_inst.row1\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2321_ net412 _1114_ net159 VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__mux2_1
X_2252_ net238 net245 VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__and2_1
XFILLER_69_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2183_ _0979_ _0980_ _0975_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_48_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1967_ net391 net57 net21 matmult_inst.fsm_inst.alu_result\[9\] VGND VGND VPWR VPWR
+ _0132_ sky130_fd_sc_hd__a22o_1
X_1898_ _0537_ _0539_ _0759_ net200 _0766_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__o221ai_1
X_3637_ clknet_leaf_10_hz100 _0497_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB1\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_3568_ clknet_leaf_20_hz100 _0428_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA1\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_2519_ matmult_inst.alu_inst.adder_inst.r1.fa3.a net174 VGND VGND VPWR VPWR _1267_
+ sky130_fd_sc_hd__and2_1
X_3499_ clknet_leaf_18_hz100 _0359_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem1\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Left_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_58_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold6 matmult_inst.alu_inst.out\[14\] VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_47_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2870_ net217 net354 net93 VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__mux2_1
XFILLER_30_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1821_ matmult_inst.mem_inst.matrixA2\[5\] net190 net182 matmult_inst.mem_inst.matrixA1\[5\]
+ _0696_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__a221o_1
X_1752_ matmult_inst.mem_inst.matrixB3\[11\] net198 _0633_ VGND VGND VPWR VPWR _0634_
+ sky130_fd_sc_hd__a21o_1
X_1683_ net268 net261 VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__and2b_1
XFILLER_7_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap103 _1450_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
Xmax_cap147 _0945_ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_1
X_3422_ clknet_leaf_2_hz100 _0282_ VGND VGND VPWR VPWR matmult_inst.alu_inst.b1_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xmax_cap158 _0975_ VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_1
X_3353_ clknet_leaf_3_hz100 _0218_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r3.fa0.b
+ sky130_fd_sc_hd__dfxtp_1
X_3284_ net293 _0011_ _0065_ VGND VGND VPWR VPWR matmult_inst.spi_inst.miso_shifter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_2304_ _1075_ _1078_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__or2_1
XFILLER_57_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2235_ _0990_ _0973_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__nand2b_1
X_2166_ _0960_ _0962_ _0959_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__a21o_1
XFILLER_65_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2097_ _0878_ _0893_ _0894_ _0895_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__nand4_1
XFILLER_80_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2999_ net436 net84 net33 VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__mux2_1
XFILLER_79_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2020_ net259 net256 net242 net244 VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__and4_1
XFILLER_75_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2922_ net598 net85 net41 VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__mux2_1
X_2853_ _1557_ _1558_ VGND VGND VPWR VPWR _1559_ sky130_fd_sc_hd__and2b_1
X_1804_ net272 net264 matmult_inst.mem_inst.mem3\[6\] VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__and3_1
X_2784_ _1492_ _1500_ VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__or2_1
X_1735_ matmult_inst.mem_inst.matrixB2\[13\] net187 net179 matmult_inst.mem_inst.matrixB1\[13\]
+ _0618_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__a221o_1
Xhold203 matmult_inst.mem_inst.matrixA2\[2\] VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 matmult_inst.alu_inst.col0\[6\] VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 matmult_inst.mem_inst.matrixB2\[1\] VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__dlygate4sd3_1
X_1666_ _0534_ matmult_inst.spi_inst.mosi_shifter\[0\] _0563_ VGND VGND VPWR VPWR
+ _0185_ sky130_fd_sc_hd__mux2_1
Xhold269 matmult_inst.mem_inst.mem3\[12\] VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 matmult_inst.mem_inst.matrixA1\[14\] VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 matmult_inst.alu_inst.adder_inst.fa.a VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 matmult_inst.fsm_inst.alu_result\[0\] VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__dlygate4sd3_1
X_3405_ clknet_leaf_3_hz100 _0266_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r2.fa1.a
+ sky130_fd_sc_hd__dfxtp_1
X_3336_ _0117_ _0203_ _0116_ VGND VGND VPWR VPWR matmult_inst.spi_inst.rx_bit_count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ clknet_leaf_21_hz100 _0156_ _0048_ VGND VGND VPWR VPWR matmult_inst.spi_inst.tx_reg_sys\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_3198_ net135 net124 VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__and2_1
X_2218_ _1013_ _1014_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__nand2_1
X_2149_ net240 net249 net247 net242 VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__a22o_1
XFILLER_53_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3121_ _0761_ _1601_ _1602_ _1137_ VGND VGND VPWR VPWR _1603_ sky130_fd_sc_hd__or4b_1
X_3052_ net282 net194 net88 VGND VGND VPWR VPWR _1591_ sky130_fd_sc_hd__and3_1
X_2003_ matmult_inst.fsm_inst.alu_result\[12\] net114 VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_18_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2905_ net484 net83 net44 VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__mux2_1
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2836_ _1537_ _1540_ _1538_ VGND VGND VPWR VPWR _1545_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_61_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2767_ matmult_inst.alu_inst.adder_inst.r0.fa2.b matmult_inst.alu_inst.adder_inst.r0.fa2.a
+ VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__nor2_1
X_2698_ _1438_ _1440_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__and2_1
XFILLER_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1718_ net269 net262 matmult_inst.mem_inst.mem3\[14\] VGND VGND VPWR VPWR _0603_
+ sky130_fd_sc_hd__and3_1
X_1649_ matmult_inst.spi_inst.mosi_shifter\[6\] matmult_inst.spi_inst.mosi_data_spi\[7\]
+ _0562_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__mux2_1
X_3319_ _0086_ _0188_ _0085_ VGND VGND VPWR VPWR matmult_inst.spi_inst.mosi_shifter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3670_ clknet_leaf_28_hz100 _0530_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.state\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2621_ _1365_ _1366_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__nand2b_1
X_2552_ _1244_ _1299_ VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__nor2_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2483_ _1218_ _1225_ _1193_ _1217_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3104_ net575 net74 net23 VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__mux2_1
X_3035_ net337 net86 net29 VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2819_ _1529_ _1530_ VGND VGND VPWR VPWR _1531_ sky130_fd_sc_hd__xor2_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_21_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1983_ matmult_inst.fsm_inst.rx_data\[2\] _0786_ net114 matmult_inst.fsm_inst.alu_result\[2\]
+ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__a22o_1
XFILLER_60_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3653_ clknet_leaf_16_hz100 _0513_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB2\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_2604_ _1346_ _1348_ _1349_ VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__o21ai_1
X_3584_ clknet_leaf_12_hz100 _0444_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA2\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_2535_ net206 net208 net224 net222 VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__and4_1
X_2466_ _1214_ _1215_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__xnor2_1
X_2397_ _1157_ net590 net66 VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_19_hz100 clknet_2_2__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_19_hz100
+ sky130_fd_sc_hd__clkbuf_8
X_3018_ net524 net84 net31 VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__mux2_1
Xwire53 _1017_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_34_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire97 net98 VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout162 _0526_ VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_4
Xfanout195 _0566_ VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_4
Xfanout184 net185 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_2
XFILLER_63_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2320_ _1112_ _1113_ VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2251_ net248 net246 net236 net234 VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__and4_1
XFILLER_69_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2182_ _0976_ _0977_ _0978_ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__a21o_1
XFILLER_80_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1966_ net580 net57 net21 matmult_inst.fsm_inst.alu_result\[8\] VGND VGND VPWR VPWR
+ _0131_ sky130_fd_sc_hd__a22o_1
X_1897_ matmult_inst.fsm_inst.state\[4\] _0539_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__or2_2
X_3636_ clknet_leaf_15_hz100 _0496_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB1\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3567_ clknet_leaf_12_hz100 _0427_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA1\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_2518_ net161 _1265_ _1266_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__a21oi_1
X_3498_ clknet_leaf_22_hz100 _0358_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem1\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_2449_ _1198_ _1199_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__nand2b_1
XFILLER_71_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold7 _0137_ VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1820_ net271 net266 matmult_inst.mem_inst.matrixA3\[5\] VGND VGND VPWR VPWR _0696_
+ sky130_fd_sc_hd__and3_1
X_1751_ matmult_inst.mem_inst.matrixB2\[11\] net186 net178 matmult_inst.mem_inst.matrixB1\[11\]
+ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__a22o_1
XFILLER_7_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap126 _0553_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
Xmax_cap104 net105 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
X_1682_ matmult_inst.mem_inst.matrixA0\[17\] net169 _0569_ net196 net115 VGND VGND
+ VPWR VPWR _0570_ sky130_fd_sc_hd__a221o_1
Xmax_cap137 _1360_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_1
X_3421_ clknet_leaf_3_hz100 _0281_ VGND VGND VPWR VPWR matmult_inst.alu_inst.a1_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xmax_cap148 _0872_ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_1
X_3352_ clknet_leaf_3_hz100 _0217_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r2.fa3.b
+ sky130_fd_sc_hd__dfxtp_1
X_2303_ _1084_ _1095_ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__xnor2_1
X_3283_ net293 _0010_ _0064_ VGND VGND VPWR VPWR matmult_inst.spi_inst.miso_shifter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_2234_ net53 _1027_ _1029_ _1030_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__a22oi_1
X_2165_ net616 _0963_ net162 VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__mux2_1
XFILLER_65_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2096_ _0893_ _0894_ _0895_ _0878_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2998_ net403 net85 net33 VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__mux2_1
XFILLER_21_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1949_ matmult_inst.spi_inst.tx_reg_sys\[15\] matmult_inst.spi_inst.miso_shifter\[14\]
+ net275 VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__mux2_1
X_3619_ clknet_leaf_16_hz100 _0479_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB0\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_8_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2921_ net446 net86 net41 VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__mux2_1
X_2852_ matmult_inst.alu_inst.adder_inst.r3.fa3.b matmult_inst.alu_inst.adder_inst.r3.fa3.a
+ VGND VGND VPWR VPWR _1558_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_13_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2783_ _1482_ _1486_ _1489_ _1493_ _1487_ VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__o311a_1
X_1803_ net618 _0680_ net91 VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__mux2_1
X_1734_ net272 net264 matmult_inst.mem_inst.matrixB3\[13\] VGND VGND VPWR VPWR _0618_
+ sky130_fd_sc_hd__and3_1
XFILLER_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold226 matmult_inst.alu_inst.out\[5\] VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 matmult_inst.fsm_inst.alu_result\[4\] VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 matmult_inst.spi_inst.mosi_data_sync\[2\] VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__dlygate4sd3_1
X_1665_ matmult_inst.spi_inst.mosi_shifter\[0\] matmult_inst.spi_inst.mosi_shifter\[1\]
+ _0563_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__mux2_1
X_3404_ clknet_leaf_0_hz100 _0265_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r2.fa0.a
+ sky130_fd_sc_hd__dfxtp_1
Xhold259 matmult_inst.mem_inst.matrixB2\[5\] VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 matmult_inst.mem_inst.matrixA1\[6\] VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 matmult_inst.mem_inst.matrixA2\[7\] VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__dlygate4sd3_1
X_3335_ _0115_ _0202_ _0114_ VGND VGND VPWR VPWR matmult_inst.spi_inst.rx_bit_count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3266_ clknet_leaf_19_hz100 _0155_ _0047_ VGND VGND VPWR VPWR matmult_inst.spi_inst.tx_reg_sys\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2217_ net238 net248 net247 net237 VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__nand4_1
X_3197_ net131 net120 VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__and2_1
X_2148_ _0945_ _0946_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_77_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2079_ net257 _0879_ _0878_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__a21bo_1
XFILLER_53_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3120_ net200 _0752_ matmult_inst.fsm_inst.state\[4\] net199 VGND VGND VPWR VPWR
+ _1602_ sky130_fd_sc_hd__and4b_1
X_3051_ net307 _0821_ net30 VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__mux2_1
X_2002_ net351 _0815_ net55 VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__mux2_1
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2904_ net485 net84 net43 VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__mux2_1
X_2835_ _1542_ _1543_ VGND VGND VPWR VPWR _1544_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_61_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2766_ net305 _1485_ net163 VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__mux2_1
X_2697_ _1413_ _1417_ _1428_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__or3_1
X_1717_ matmult_inst.mem_inst.matrixA0\[14\] net168 _0601_ net195 net115 VGND VGND
+ VPWR VPWR _0602_ sky130_fd_sc_hd__a221o_1
X_1648_ matmult_inst.spi_inst.rx_bit_count\[2\] net1 _0558_ VGND VGND VPWR VPWR _0562_
+ sky130_fd_sc_hd__nand3_4
X_3318_ _0084_ _0187_ _0083_ VGND VGND VPWR VPWR matmult_inst.spi_inst.mosi_shifter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3249_ clknet_leaf_5_hz100 matmult_inst.spi_inst.mosi_data_spi\[6\] _0030_ VGND VGND
+ VPWR VPWR matmult_inst.spi_inst.mosi_data_sync\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2620_ _1313_ _1363_ _1364_ VGND VGND VPWR VPWR _1366_ sky130_fd_sc_hd__or3_1
X_2551_ _1243_ net62 VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__nor2_1
X_2482_ net648 _1231_ net161 VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__mux2_1
XFILLER_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3103_ net416 net75 net23 VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__mux2_1
X_3034_ net339 net87 net30 VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2818_ _1516_ _1521_ _1524_ _1522_ VGND VGND VPWR VPWR _1530_ sky130_fd_sc_hd__o31a_1
X_2749_ net246 net388 net95 VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1982_ net415 net86 net55 VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3652_ clknet_leaf_8_hz100 _0512_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB2\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_2603_ net205 net221 VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__and2_1
X_3583_ clknet_leaf_10_hz100 _0443_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA2\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2534_ net206 net224 net222 net208 VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__a22oi_1
X_2465_ _1197_ _1198_ _1199_ VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__o21ai_2
X_2396_ _1156_ net489 net66 VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__mux2_1
XFILLER_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3017_ net497 net85 net31 VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__mux2_1
Xwire98 net99 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_34_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout130 net132 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
Xfanout174 net175 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__buf_2
Xfanout163 net164 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_4
Xfanout185 _0572_ VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
Xfanout196 _0566_ VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2250_ net246 net236 net234 net248 VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__a22oi_1
XFILLER_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2181_ _0976_ _0977_ _0978_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_48_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1965_ matmult_inst.alu_inst.out\[7\] _0794_ net22 net536 VGND VGND VPWR VPWR _0130_
+ sky130_fd_sc_hd__a22o_1
X_1896_ matmult_inst.fsm_inst.state\[4\] _0539_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__nor2_1
X_3635_ clknet_leaf_16_hz100 _0495_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB1\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3566_ clknet_leaf_12_hz100 _0426_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA1\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3497_ clknet_leaf_23_hz100 _0357_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem1\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_2517_ net641 net161 VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__nor2_1
X_2448_ net225 net211 net213 net223 VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__a22o_1
X_2379_ _1159_ net354 net108 VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold8 matmult_inst.alu_inst.row0\[5\] VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1750_ matmult_inst.mem_inst.matrixA0\[11\] net168 _0631_ net195 net115 VGND VGND
+ VPWR VPWR _0632_ sky130_fd_sc_hd__a221o_1
XFILLER_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap105 _1327_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_18_hz100 clknet_2_2__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_18_hz100
+ sky130_fd_sc_hd__clkbuf_8
X_1681_ net280 matmult_inst.mem_inst.mem0\[17\] matmult_inst.mem_inst.matrixB0\[17\]
+ net286 VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__a22o_1
Xmax_cap138 _1325_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_1
X_3420_ clknet_leaf_4_hz100 _0280_ VGND VGND VPWR VPWR matmult_inst.alu_inst.a1_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3351_ clknet_leaf_3_hz100 _0216_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r2.fa2.b
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2302_ _1095_ _1084_ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__and2b_1
X_3282_ net293 _0009_ _0063_ VGND VGND VPWR VPWR matmult_inst.spi_inst.miso_shifter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_2233_ net53 _1028_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__or2_1
X_2164_ _0961_ _0962_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2095_ net257 net235 _0876_ net173 _0846_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__a41o_1
XFILLER_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2997_ net442 net86 net33 VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__mux2_1
X_1948_ matmult_inst.spi_inst.tx_reg_sys\[14\] matmult_inst.spi_inst.miso_shifter\[13\]
+ net275 VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__mux2_1
X_1879_ net281 _0743_ _0746_ net285 VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__a22o_1
X_3618_ clknet_leaf_15_hz100 _0478_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB0\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3549_ clknet_leaf_13_hz100 _0409_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA0\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_48_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2920_ net543 net87 net42 VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__mux2_1
X_2851_ matmult_inst.alu_inst.adder_inst.r3.fa3.b matmult_inst.alu_inst.adder_inst.r3.fa3.a
+ VGND VGND VPWR VPWR _1557_ sky130_fd_sc_hd__nor2_1
XFILLER_79_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2782_ _1497_ _1498_ VGND VGND VPWR VPWR _1499_ sky130_fd_sc_hd__and2b_1
X_1802_ matmult_inst.mem_inst.matrixA0\[7\] net168 _0678_ _0679_ VGND VGND VPWR VPWR
+ _0680_ sky130_fd_sc_hd__a211o_1
X_1733_ matmult_inst.mem_inst.mem3\[13\] net198 _0616_ VGND VGND VPWR VPWR _0617_
+ sky130_fd_sc_hd__a21o_1
XFILLER_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold216 matmult_inst.alu_inst.adder_inst.r0.fa2.b VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 _0161_ VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__dlygate4sd3_1
X_1664_ matmult_inst.spi_inst.mosi_shifter\[1\] matmult_inst.spi_inst.mosi_shifter\[2\]
+ _0563_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__mux2_1
Xhold238 matmult_inst.mem_inst.matrixA0\[2\] VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__dlygate4sd3_1
X_3403_ clknet_leaf_0_hz100 _0264_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r1.fa3.a
+ sky130_fd_sc_hd__dfxtp_1
Xhold249 matmult_inst.mem_inst.mem1\[0\] VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 matmult_inst.mem_inst.matrixB3\[9\] VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ clknet_leaf_9_hz100 matmult_inst.cs _0113_ VGND VGND VPWR VPWR matmult_inst.spi_inst.cs_sync
+ sky130_fd_sc_hd__dfstp_1
X_3265_ clknet_leaf_18_hz100 _0154_ _0046_ VGND VGND VPWR VPWR matmult_inst.spi_inst.tx_reg_sys\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2216_ net238 net247 net236 net248 VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__a22o_1
XFILLER_38_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3196_ net132 net119 VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__and2_1
XFILLER_81_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2147_ _0939_ _0943_ _0944_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__nand3_1
X_2078_ net235 _0876_ net173 VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__and3_1
XFILLER_30_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3050_ net327 net71 net30 VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__mux2_1
X_2001_ matmult_inst.fsm_inst.alu_result\[11\] net114 VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_18_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2903_ net461 net85 net43 VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__mux2_1
X_2834_ matmult_inst.alu_inst.adder_inst.r3.fa0.b matmult_inst.alu_inst.adder_inst.r3.fa0.a
+ VGND VGND VPWR VPWR _1543_ sky130_fd_sc_hd__nand2_1
X_2765_ _1480_ _1484_ VGND VGND VPWR VPWR _1485_ sky130_fd_sc_hd__xnor2_1
X_2696_ _1438_ VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__inv_2
X_1716_ net278 matmult_inst.mem_inst.mem0\[14\] matmult_inst.mem_inst.matrixB0\[14\]
+ net283 VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__a22o_1
X_1647_ _0557_ _0561_ net1 VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__and3b_1
Xwire6 _1561_ VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_3317_ _0082_ _0186_ _0081_ VGND VGND VPWR VPWR matmult_inst.spi_inst.mosi_shifter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3248_ clknet_leaf_5_hz100 matmult_inst.spi_inst.mosi_data_spi\[5\] _0029_ VGND VGND
+ VPWR VPWR matmult_inst.spi_inst.mosi_data_sync\[5\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3179_ net135 net123 VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__and2_1
XFILLER_26_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2550_ _1279_ _1280_ net61 VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__a21o_1
X_2481_ _1229_ _1230_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__xnor2_1
X_3102_ net361 net76 net23 VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__mux2_1
X_3033_ net198 _0567_ net88 VGND VGND VPWR VPWR _1590_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_66_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2817_ _1527_ _1528_ VGND VGND VPWR VPWR _1529_ sky130_fd_sc_hd__nand2b_1
X_2748_ net248 net379 net95 VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__mux2_1
X_2679_ _1421_ _1422_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1981_ matmult_inst.fsm_inst.rx_data\[1\] _0786_ net113 matmult_inst.fsm_inst.alu_result\[1\]
+ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_71_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3651_ clknet_leaf_25_hz100 _0511_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB2\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2602_ net224 net222 net202 net204 VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__and4_1
X_3582_ clknet_leaf_16_hz100 _0442_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA2\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2533_ _1248_ _1250_ _1249_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__a21bo_1
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2464_ _1212_ _1213_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__nand2_1
X_2395_ _1155_ net595 _1163_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire11 _1546_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
X_3016_ net410 net86 net31 VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__mux2_1
Xwire99 net101 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_34_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout131 net132 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
Xfanout120 net121 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_2
Xfanout164 _0003_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_4
Xfanout186 net187 VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__buf_2
Xfanout175 _0822_ VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__buf_2
XFILLER_47_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2180_ net250 net236 VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_76_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1964_ net346 net57 net22 matmult_inst.fsm_inst.alu_result\[6\] VGND VGND VPWR VPWR
+ _0129_ sky130_fd_sc_hd__a22o_1
X_1895_ net199 net200 _0762_ _0761_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__a31o_1
X_3634_ clknet_leaf_10_hz100 _0494_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB1\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3565_ clknet_leaf_10_hz100 _0425_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA1\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3496_ clknet_leaf_20_hz100 _0356_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem1\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_2516_ _1262_ _1264_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__xnor2_1
X_2447_ net225 net223 net211 net213 VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__and4_1
X_2378_ _0690_ net167 VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_39_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_18_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold9 matmult_inst.mem_inst.matrixB3\[16\] VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_74_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1680_ _0567_ net194 net287 VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__mux2_1
Xmax_cap106 _1274_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__buf_1
Xmax_cap139 _1287_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__buf_1
X_3350_ clknet_leaf_3_hz100 _0215_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r2.fa1.b
+ sky130_fd_sc_hd__dfxtp_1
X_2301_ _1070_ _1073_ _1071_ VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__o21ai_1
X_3281_ net292 _0008_ _0062_ VGND VGND VPWR VPWR matmult_inst.spi_inst.miso_shifter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2232_ net53 _1028_ _1027_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__a21oi_1
X_2163_ _0883_ _0918_ _0920_ _0917_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__a31o_1
XFILLER_65_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2094_ net257 net255 net233 net235 VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__nand4_2
XFILLER_61_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2996_ net475 net87 net34 VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__mux2_1
X_1947_ matmult_inst.spi_inst.tx_reg_sys\[13\] matmult_inst.spi_inst.miso_shifter\[12\]
+ net275 VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__mux2_1
X_1878_ net195 _0744_ _0748_ net288 VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__a22o_1
X_3617_ clknet_leaf_7_hz100 _0477_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB0\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3548_ clknet_leaf_16_hz100 _0408_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA0\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3479_ clknet_leaf_18_hz100 _0339_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem0\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2850_ net300 net8 net164 VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__mux2_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1801_ net195 _0673_ _0677_ net288 VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__a22o_1
X_2781_ matmult_inst.alu_inst.adder_inst.r1.fa0.b matmult_inst.alu_inst.adder_inst.r1.fa0.a
+ VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_13_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1732_ matmult_inst.mem_inst.mem2\[13\] net187 net179 matmult_inst.mem_inst.mem1\[13\]
+ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__a22o_1
XFILLER_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold217 matmult_inst.mem_inst.matrixB0\[1\] VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold206 matmult_inst.alu_inst.adder_inst.r0.fa0.b VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__dlygate4sd3_1
X_1663_ matmult_inst.spi_inst.mosi_shifter\[2\] matmult_inst.spi_inst.mosi_shifter\[3\]
+ _0563_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__mux2_1
Xhold239 matmult_inst.alu_inst.col0\[7\] VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__dlygate4sd3_1
X_3402_ clknet_leaf_1_hz100 _0263_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r1.fa2.a
+ sky130_fd_sc_hd__dfxtp_1
Xhold228 matmult_inst.spi_inst.mosi_data_sync\[4\] VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__dlygate4sd3_1
X_3333_ _0112_ _0201_ _0111_ VGND VGND VPWR VPWR matmult_inst.spi_inst.mosi_data_spi\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3264_ clknet_leaf_11_hz100 _0153_ _0045_ VGND VGND VPWR VPWR matmult_inst.spi_inst.tx_reg_sys\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_2215_ net240 matmult_inst.alu_inst.a1_reg\[7\] VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__nand2_1
X_3195_ net133 net122 VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__and2_1
X_2146_ _0943_ _0944_ _0939_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__a21oi_1
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2077_ net257 net235 _0876_ net173 VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__a22o_1
XFILLER_81_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2979_ net532 net85 net35 VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__mux2_1
XFILLER_30_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_17_hz100 clknet_2_2__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_17_hz100
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_55_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2000_ net316 net77 net55 VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__mux2_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2902_ net596 _0805_ net43 VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__mux2_1
XFILLER_31_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2833_ matmult_inst.alu_inst.adder_inst.r3.fa0.b matmult_inst.alu_inst.adder_inst.r3.fa0.a
+ VGND VGND VPWR VPWR _1542_ sky130_fd_sc_hd__or2_1
X_2764_ _1482_ _1483_ VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__nor2_1
X_1715_ net647 net92 _0592_ _0600_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__o22a_1
X_2695_ _1413_ _1417_ _1428_ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__o21ai_2
X_1646_ matmult_inst.spi_inst.rx_bit_count\[0\] matmult_inst.spi_inst.rx_bit_count\[3\]
+ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__nand2b_1
X_3316_ _0080_ _0185_ _0079_ VGND VGND VPWR VPWR matmult_inst.spi_inst.mosi_shifter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3247_ clknet_leaf_5_hz100 matmult_inst.spi_inst.mosi_data_spi\[4\] _0028_ VGND VGND
+ VPWR VPWR matmult_inst.spi_inst.mosi_data_sync\[4\] sky130_fd_sc_hd__dfrtp_1
X_3178_ net134 net123 VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__and2_1
X_2129_ _0924_ _0925_ _0903_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__a21o_1
XFILLER_25_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2480_ _1188_ _1207_ _1208_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__a21bo_1
X_3101_ net587 _0814_ net23 VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__mux2_1
X_3032_ net364 _0821_ net32 VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2816_ matmult_inst.alu_inst.adder_inst.r2.fa1.b matmult_inst.alu_inst.adder_inst.r2.fa1.a
+ VGND VGND VPWR VPWR _1528_ sky130_fd_sc_hd__nand2_1
XFILLER_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2747_ net250 net493 net95 VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__mux2_1
X_2678_ _1388_ _1395_ _1397_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__o21a_1
X_1629_ _0538_ _0547_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__nor2_1
XFILLER_27_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1980_ net325 net87 net55 VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__mux2_1
XFILLER_60_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3650_ clknet_leaf_23_hz100 _0510_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB2\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2601_ net224 net202 net203 net222 VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__a22o_1
X_3581_ clknet_leaf_8_hz100 _0441_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA2\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_2532_ _1275_ _1276_ _1278_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__nand3_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2463_ net225 net210 net223 net211 VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__a22o_1
X_2394_ _1154_ net367 net66 VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3015_ net441 net87 net32 VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__mux2_1
Xwire45 _1535_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_1
XFILLER_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout121 net122 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout132 net133 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
Xfanout198 _0535_ VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__buf_2
Xfanout187 net193 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_4
XFILLER_74_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1963_ net520 net57 net22 net550 VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__a22o_1
X_1894_ net199 matmult_inst.fsm_inst.state\[3\] VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__nand2_1
X_3633_ clknet_leaf_25_hz100 _0493_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB1\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3564_ clknet_leaf_16_hz100 _0424_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA1\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_2515_ _1227_ _1263_ VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__nor2_1
X_3495_ clknet_leaf_13_hz100 _0355_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem1\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_2446_ net221 matmult_inst.alu_inst.b0_reg\[0\] VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__and2_1
X_2377_ _1158_ net302 net108 VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__mux2_1
XFILLER_56_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap107 _1225_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_1
X_2300_ _1081_ _1085_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__nand2_1
X_3280_ net292 _0022_ _0061_ VGND VGND VPWR VPWR matmult_inst.spi_inst.miso_shifter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2231_ _1018_ _1025_ _1026_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__nand3_1
XFILLER_78_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2162_ _0959_ _0960_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__nand2b_1
X_2093_ net257 net232 net235 net255 VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__a22o_1
X_2995_ _0567_ net178 net88 VGND VGND VPWR VPWR _1588_ sky130_fd_sc_hd__and3_1
XFILLER_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1946_ matmult_inst.spi_inst.tx_reg_sys\[12\] matmult_inst.spi_inst.miso_shifter\[11\]
+ net275 VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__mux2_1
X_1877_ matmult_inst.mem_inst.matrixA2\[0\] net189 net181 matmult_inst.mem_inst.matrixA1\[0\]
+ _0747_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__a221o_1
X_3616_ clknet_leaf_8_hz100 _0476_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB0\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3547_ clknet_leaf_8_hz100 _0407_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA0\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_3478_ clknet_leaf_20_hz100 _0338_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem0\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_2429_ net228 net226 net210 net211 VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_42_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1800_ net280 _0672_ _0675_ net285 VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__a22o_1
X_2780_ matmult_inst.alu_inst.adder_inst.r1.fa0.b matmult_inst.alu_inst.adder_inst.r1.fa0.a
+ VGND VGND VPWR VPWR _1497_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_13_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1731_ net288 _0614_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__and2_1
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold207 matmult_inst.mem_inst.matrixB1\[4\] VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__dlygate4sd3_1
X_1662_ matmult_inst.spi_inst.mosi_shifter\[3\] matmult_inst.spi_inst.mosi_shifter\[4\]
+ _0563_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__mux2_1
Xhold218 matmult_inst.mem_inst.matrixB0\[15\] VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__dlygate4sd3_1
X_3401_ clknet_leaf_1_hz100 _0262_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r1.fa1.a
+ sky130_fd_sc_hd__dfxtp_1
Xhold229 _0163_ VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__dlygate4sd3_1
X_3332_ _0110_ _0200_ _0109_ VGND VGND VPWR VPWR matmult_inst.spi_inst.mosi_data_spi\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_37_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3263_ clknet_leaf_10_hz100 _0152_ _0044_ VGND VGND VPWR VPWR matmult_inst.spi_inst.tx_reg_sys\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_3194_ net133 net122 VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__and2_1
X_2214_ _1009_ _1010_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__nor2_1
X_2145_ _0940_ _0941_ _0942_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__o21ai_1
XFILLER_38_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2076_ net242 matmult_inst.alu_inst.b1_reg\[0\] net250 net249 VGND VGND VPWR VPWR
+ _0877_ sky130_fd_sc_hd__nand4_1
XFILLER_34_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2978_ net454 _0805_ net35 VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__mux2_1
X_1929_ net155 _0793_ net58 _0795_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__or4_1
XFILLER_30_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_hz100 hz100 VGND VGND VPWR VPWR clknet_0_hz100 sky130_fd_sc_hd__clkbuf_16
XFILLER_30_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Left_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_64_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Left_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold90 matmult_inst.alu_inst.col1\[5\] VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2901_ net560 net87 net43 VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__mux2_1
X_2832_ net476 net15 net164 VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__mux2_1
X_2763_ matmult_inst.alu_inst.adder_inst.r0.fa1.b matmult_inst.alu_inst.adder_inst.r0.fa1.a
+ VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__and2_1
X_1714_ net287 _0596_ _0599_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__a21o_1
X_2694_ net611 _1437_ net159 VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__mux2_1
X_1645_ _0558_ _0560_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__nor2_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire8 _1556_ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
X_3315_ clknet_leaf_10_hz100 matmult_inst.spi_inst.rx_done_spi _0078_ VGND VGND VPWR
+ VPWR matmult_inst.spi_inst.rx_done1 sky130_fd_sc_hd__dfrtp_1
X_3246_ clknet_leaf_5_hz100 matmult_inst.spi_inst.mosi_data_spi\[3\] _0027_ VGND VGND
+ VPWR VPWR matmult_inst.spi_inst.mosi_data_sync\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_39_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3177_ net134 net123 VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__and2_1
X_2128_ _0903_ _0924_ _0925_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__nand3_1
XFILLER_81_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2059_ _0836_ _0841_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__nor2_1
XFILLER_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3100_ net365 _0813_ net24 VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__mux2_1
X_3031_ net387 _0820_ net32 VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2815_ matmult_inst.alu_inst.adder_inst.r2.fa1.b matmult_inst.alu_inst.adder_inst.r2.fa1.a
+ VGND VGND VPWR VPWR _1527_ sky130_fd_sc_hd__nor2_1
XFILLER_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2746_ net252 net377 net95 VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__mux2_1
X_2677_ _1419_ _1420_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_16_hz100 clknet_2_3__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_16_hz100
+ sky130_fd_sc_hd__clkbuf_8
X_1628_ matmult_inst.fsm_inst.state\[0\] matmult_inst.fsm_inst.state\[1\] VGND VGND
+ VPWR VPWR _0547_ sky130_fd_sc_hd__nand2b_1
X_3229_ clknet_leaf_6_hz100 _0127_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.alu_result\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2600_ net224 net202 net204 net222 VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__a22oi_1
X_3580_ clknet_leaf_8_hz100 _0440_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA2\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_2531_ _1275_ _1276_ _1278_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__a21o_1
XFILLER_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2462_ net225 net209 net223 net212 VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__nand4_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2393_ _1153_ net600 net66 VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__mux2_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3014_ _0567_ net186 net88 VGND VGND VPWR VPWR _1589_ sky130_fd_sc_hd__and3_1
Xwire13 _1430_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire46 _1531_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
Xwire68 _0956_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2729_ _1433_ _1453_ _1457_ net12 VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__a31o_1
Xfanout122 net126 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
Xfanout133 _0546_ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout166 net167 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__buf_2
Xfanout199 matmult_inst.fsm_inst.state\[2\] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_2
Xfanout188 net193 VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1962_ net570 net57 net22 net509 VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__a22o_1
X_1893_ _0551_ _0759_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__nand2_1
X_3632_ clknet_leaf_25_hz100 _0492_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB1\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3563_ clknet_leaf_8_hz100 _0423_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA1\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_2514_ _1211_ net51 _1230_ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__a21oi_1
X_3494_ clknet_leaf_12_hz100 _0354_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem1\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_2445_ _1180_ _1193_ _1194_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2376_ _0701_ net167 VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__and2_2
XFILLER_56_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap108 _1152_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_2
XFILLER_23_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2230_ _1025_ _1026_ _1018_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__a21oi_1
XFILLER_38_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2161_ _0957_ _0958_ _0923_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__a21o_1
X_2092_ net257 net232 VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2994_ net360 net70 net36 VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__mux2_1
X_1945_ matmult_inst.spi_inst.tx_reg_sys\[11\] matmult_inst.spi_inst.miso_shifter\[10\]
+ net276 VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__mux2_1
X_1876_ net271 net263 matmult_inst.mem_inst.matrixA3\[0\] VGND VGND VPWR VPWR _0747_
+ sky130_fd_sc_hd__and3_1
X_3615_ clknet_leaf_25_hz100 _0475_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB0\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3546_ clknet_leaf_16_hz100 _0406_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA0\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3477_ clknet_leaf_13_hz100 _0337_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem0\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_2428_ net228 net226 net210 net211 VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__and4_1
X_2359_ net267 _1139_ _1141_ _1147_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__o22a_1
XFILLER_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1730_ matmult_inst.mem_inst.matrixA2\[13\] net187 net179 matmult_inst.mem_inst.matrixA1\[13\]
+ _0613_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__a221o_1
Xhold208 matmult_inst.mem_inst.matrixB2\[3\] VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__dlygate4sd3_1
X_1661_ matmult_inst.spi_inst.mosi_shifter\[4\] matmult_inst.spi_inst.mosi_shifter\[5\]
+ _0563_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__mux2_1
Xhold219 matmult_inst.alu_inst.row0\[4\] VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__dlygate4sd3_1
X_3400_ clknet_leaf_1_hz100 _0261_ VGND VGND VPWR VPWR matmult_inst.alu_inst.adder_inst.r1.fa0.a
+ sky130_fd_sc_hd__dfxtp_1
X_3331_ _0108_ _0199_ _0107_ VGND VGND VPWR VPWR matmult_inst.spi_inst.mosi_data_spi\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3262_ clknet_leaf_12_hz100 _0151_ _0043_ VGND VGND VPWR VPWR matmult_inst.spi_inst.tx_reg_sys\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2213_ _1001_ _1006_ _1007_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__and3_1
X_3193_ net130 net118 VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__and2_1
X_2144_ _0940_ _0941_ _0942_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__or3_1
XFILLER_38_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2075_ net242 net250 net248 net244 VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__a22o_1
XFILLER_34_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2977_ net413 net87 net35 VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__mux2_1
X_1928_ _1606_ _0784_ _0541_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__a21oi_1
X_1859_ net643 _0731_ net92 VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__mux2_1
XFILLER_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3529_ clknet_leaf_8_hz100 _0389_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem3\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold91 matmult_inst.mem_inst.matrixA0\[11\] VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 matmult_inst.mem_inst.mem2\[17\] VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2900_ net277 net194 net88 VGND VGND VPWR VPWR _1583_ sky130_fd_sc_hd__and3_1
X_2831_ _1539_ _1540_ VGND VGND VPWR VPWR _1541_ sky130_fd_sc_hd__xnor2_1
XFILLER_77_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2762_ matmult_inst.alu_inst.adder_inst.r0.fa1.b matmult_inst.alu_inst.adder_inst.r0.fa1.a
+ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__nor2_1
X_1713_ net283 _0594_ _0598_ net278 VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__a22o_1
X_2693_ _1434_ _1436_ VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__xor2_1
X_1644_ matmult_inst.spi_inst.rx_bit_count\[1\] _0557_ net1 VGND VGND VPWR VPWR _0560_
+ sky130_fd_sc_hd__o21ai_1
Xwire9 _1551_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
X_3314_ clknet_leaf_13_hz100 _0184_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB3\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_3245_ clknet_leaf_5_hz100 matmult_inst.spi_inst.mosi_data_spi\[2\] _0026_ VGND VGND
+ VPWR VPWR matmult_inst.spi_inst.mosi_data_sync\[2\] sky130_fd_sc_hd__dfrtp_1
X_3176_ net133 net116 VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_16_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2127_ _0903_ _0924_ _0925_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__and3_1
XFILLER_81_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2058_ _0851_ _0852_ net149 VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_52_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3030_ net514 net72 net31 VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2814_ net580 _1526_ net163 VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__mux2_1
X_2745_ net254 net613 net96 VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__mux2_1
X_2676_ _1385_ _1418_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__or2_1
X_1627_ net198 _0541_ _0545_ matmult_inst.fsm_inst.tx_start_send VGND VGND VPWR VPWR
+ _0546_ sky130_fd_sc_hd__or4b_4
X_3228_ clknet_leaf_1_hz100 net381 VGND VGND VPWR VPWR matmult_inst.fsm_inst.alu_result\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_29_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3159_ net134 net123 VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__and2_1
XFILLER_14_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2530_ _1237_ _1277_ VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__nand2_1
XFILLER_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2461_ _1195_ _1202_ VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__nor2_1
X_2392_ _0766_ _0774_ _1162_ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__o21ai_1
X_3013_ net408 net70 net34 VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__mux2_1
Xwire14 _1377_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
Xwire69 _0914_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_34_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2728_ net48 _1467_ VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__xnor2_1
X_2659_ _1402_ _1403_ VGND VGND VPWR VPWR _1404_ sky130_fd_sc_hd__nand2_1
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout134 net135 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_2
Xfanout123 net124 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
Xfanout167 _0765_ VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_2
Xfanout178 net179 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__buf_2
Xfanout189 net192 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_hz100 clknet_2_3__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_15_hz100
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1961_ net380 net57 net22 matmult_inst.fsm_inst.alu_result\[3\] VGND VGND VPWR VPWR
+ _0126_ sky130_fd_sc_hd__a22o_1
XFILLER_53_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1892_ _0757_ _0759_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_31_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3631_ clknet_leaf_17_hz100 _0491_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB1\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3562_ clknet_leaf_8_hz100 _0422_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA1\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_2513_ _1259_ _1261_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__nor2_1
X_3493_ clknet_leaf_8_hz100 _0353_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem1\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2444_ _1193_ _1194_ _1180_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__a21oi_1
X_2375_ _1157_ net513 net108 VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__mux2_1
XFILLER_59_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2160_ _0923_ _0957_ _0958_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__and3_1
X_2091_ _0870_ _0871_ _0890_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2993_ net526 net71 net36 VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__mux2_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1944_ matmult_inst.spi_inst.tx_reg_sys\[10\] matmult_inst.spi_inst.miso_shifter\[9\]
+ net275 VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__mux2_1
X_3614_ clknet_leaf_25_hz100 _0474_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB0\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1875_ matmult_inst.mem_inst.matrixB2\[0\] net189 net181 matmult_inst.mem_inst.matrixB1\[0\]
+ _0745_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__a221o_1
X_3545_ clknet_leaf_7_hz100 _0405_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA0\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3476_ clknet_leaf_16_hz100 _0336_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem0\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_2427_ _1177_ _1178_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__nor2_1
X_2358_ _1604_ net90 _0771_ _1146_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__a31o_1
X_2289_ net248 net230 _1044_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__and3_1
XFILLER_52_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire140 _1272_ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_1
X_1660_ matmult_inst.spi_inst.mosi_shifter\[5\] matmult_inst.spi_inst.mosi_shifter\[6\]
+ _0563_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__mux2_1
Xhold209 matmult_inst.mem_inst.matrixA1\[11\] VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__dlygate4sd3_1
X_3330_ _0106_ _0198_ _0105_ VGND VGND VPWR VPWR matmult_inst.spi_inst.mosi_data_spi\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3261_ clknet_leaf_12_hz100 _0150_ _0042_ VGND VGND VPWR VPWR matmult_inst.spi_inst.tx_reg_sys\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2212_ _1008_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__inv_2
X_3192_ net130 net118 VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__and2_1
X_2143_ net238 net250 VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__and2_1
X_2074_ _0849_ _0873_ _0874_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__a21oi_1
XFILLER_46_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2976_ net194 _0567_ net88 VGND VGND VPWR VPWR _1587_ sky130_fd_sc_hd__and3_1
X_1927_ matmult_inst.alu_inst.complete _0780_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__and2_1
X_1858_ matmult_inst.mem_inst.matrixA0\[2\] net168 _0729_ _0730_ VGND VGND VPWR VPWR
+ _0731_ sky130_fd_sc_hd__a211o_1
X_1789_ matmult_inst.mem_inst.mem2\[8\] net191 net183 matmult_inst.mem_inst.mem1\[8\]
+ _0667_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__a221o_1
XFILLER_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3528_ clknet_leaf_16_hz100 _0388_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem3\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_3459_ clknet_leaf_28_hz100 _0319_ VGND VGND VPWR VPWR matmult_inst.alu_inst.b0_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold70 matmult_inst.mem_inst.matrixA2\[17\] VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 matmult_inst.mem_inst.matrixA0\[5\] VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 matmult_inst.alu_inst.col1\[2\] VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_18_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2830_ _1532_ net45 _1533_ VGND VGND VPWR VPWR _1540_ sky130_fd_sc_hd__a21bo_1
X_2761_ net569 _0796_ _1480_ _1481_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__a22o_1
X_1712_ matmult_inst.mem_inst.mem2\[15\] net188 net180 matmult_inst.mem_inst.mem1\[15\]
+ _0597_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__a221o_1
X_2692_ _1407_ _1435_ VGND VGND VPWR VPWR _1436_ sky130_fd_sc_hd__and2b_1
X_1643_ matmult_inst.spi_inst.rx_bit_count\[2\] _0558_ _0559_ VGND VGND VPWR VPWR
+ _0204_ sky130_fd_sc_hd__o21a_1
XFILLER_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_1 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3313_ clknet_leaf_14_hz100 _0183_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB3\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_3244_ clknet_leaf_9_hz100 matmult_inst.spi_inst.mosi_data_spi\[1\] _0025_ VGND VGND
+ VPWR VPWR matmult_inst.spi_inst.mosi_data_sync\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3175_ net127 net116 VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__and2_1
XFILLER_66_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2126_ net257 net255 net231 net232 VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__nand4_1
XFILLER_81_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2057_ _0851_ _0852_ net149 VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_52_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2959_ net371 net86 net37 VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__mux2_1
XFILLER_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2813_ _1523_ _1525_ VGND VGND VPWR VPWR _1526_ sky130_fd_sc_hd__xnor2_1
X_2744_ net256 net456 net96 VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__mux2_1
X_2675_ _1385_ _1418_ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__and2_1
X_1626_ _0542_ net197 VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__nand2_1
X_3227_ clknet_leaf_26_hz100 net425 VGND VGND VPWR VPWR matmult_inst.fsm_inst.alu_result\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3158_ net133 net122 VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__and2_1
X_2109_ _0905_ _0907_ _0908_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__o21bai_1
XFILLER_14_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3089_ net401 net70 net26 VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__mux2_1
XFILLER_22_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2460_ net640 _1210_ net161 VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__mux2_1
X_2391_ _0564_ net166 _0784_ net150 VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_79_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3012_ net435 _0820_ net34 VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__mux2_1
Xwire15 _1541_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
Xwire48 _1466_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_1
XFILLER_36_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2727_ net47 _1467_ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__nor2_1
X_2658_ _1366_ _1369_ _1365_ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__a21o_1
X_1609_ net1 VGND VGND VPWR VPWR matmult_inst.cs sky130_fd_sc_hd__inv_2
X_2589_ net60 _1333_ _1331_ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__a21oi_1
Xfanout113 net114 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_4
Xfanout124 net125 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
Xfanout135 net136 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
Xfanout179 net185 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__buf_2
Xfanout168 _0568_ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_4
XFILLER_74_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1960_ net424 net58 net21 matmult_inst.fsm_inst.alu_result\[2\] VGND VGND VPWR VPWR
+ _0125_ sky130_fd_sc_hd__a22o_1
X_1891_ _0759_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3630_ clknet_leaf_17_hz100 _0490_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB1\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3561_ clknet_leaf_25_hz100 _0421_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA1\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2512_ _1232_ _1257_ _1258_ VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__and3_1
XFILLER_52_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3492_ clknet_leaf_15_hz100 _0352_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem1\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_2443_ _1191_ _1192_ _1178_ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__a21o_1
X_2374_ _0711_ net167 VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__and2_2
XFILLER_68_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2090_ _0870_ _0871_ _0847_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__a21o_1
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2992_ net414 net72 net35 VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1943_ matmult_inst.spi_inst.tx_reg_sys\[9\] matmult_inst.spi_inst.miso_shifter\[8\]
+ net275 VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__mux2_1
X_3613_ clknet_leaf_26_hz100 _0473_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB0\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1874_ net271 net263 matmult_inst.mem_inst.matrixB3\[0\] VGND VGND VPWR VPWR _0745_
+ sky130_fd_sc_hd__and3_1
X_3544_ clknet_leaf_8_hz100 _0404_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA0\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3475_ clknet_leaf_16_hz100 _0335_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem0\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2426_ net225 net223 net213 matmult_inst.alu_inst.b0_reg\[0\] VGND VGND VPWR VPWR
+ _1178_ sky130_fd_sc_hd__and4_1
XFILLER_69_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2357_ _0758_ _1143_ _1144_ _1145_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__or4_1
X_2288_ net250 net230 net233 net248 VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__a22oi_1
XFILLER_52_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_hz100 clknet_2_3__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_14_hz100
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_hz100 clknet_2_0__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_29_hz100
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_47_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ clknet_leaf_11_hz100 _0149_ _0041_ VGND VGND VPWR VPWR matmult_inst.spi_inst.tx_reg_sys\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2211_ _1006_ _1007_ _1001_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__a21o_1
X_3191_ net131 net120 VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__and2_1
XFILLER_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2142_ net253 net251 net236 net234 VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__and4_1
X_2073_ _0849_ _0872_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__nor2_1
XFILLER_61_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2975_ net304 net70 net38 VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__mux2_1
X_1926_ _0776_ _0780_ net277 VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__o21a_1
X_1857_ net194 _0724_ _0728_ net287 VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__a22o_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3527_ clknet_leaf_8_hz100 _0387_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem3\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_1788_ net273 net265 matmult_inst.mem_inst.mem3\[8\] VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__and3_1
X_3458_ clknet_leaf_28_hz100 _0318_ VGND VGND VPWR VPWR matmult_inst.alu_inst.b0_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2409_ _1159_ net399 net63 VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__mux2_1
X_3389_ clknet_leaf_6_hz100 _0251_ VGND VGND VPWR VPWR matmult_inst.alu_inst.col1\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_69_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_24_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_33_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold82 matmult_inst.mem_inst.matrixA3\[12\] VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 matmult_inst.alu_inst.row0\[6\] VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 matmult_inst.mem_inst.matrixB2\[9\] VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 matmult_inst.mem_inst.matrixA2\[16\] VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2760_ matmult_inst.alu_inst.adder_inst.r0.fa0.b matmult_inst.alu_inst.adder_inst.r0.fa0.a
+ net163 VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__o21a_1
X_1711_ net268 net261 matmult_inst.mem_inst.mem3\[15\] VGND VGND VPWR VPWR _0597_
+ sky130_fd_sc_hd__and3_1
X_2691_ _1339_ _1376_ _1380_ _1408_ _1377_ VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__a311o_1
XANTENNA_2 matmult_inst.fsm_inst.alu_result\[17\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1642_ matmult_inst.spi_inst.rx_bit_count\[2\] _0558_ matmult_inst.cs VGND VGND VPWR
+ VPWR _0559_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3312_ clknet_leaf_21_hz100 _0182_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB3\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_60_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3243_ clknet_leaf_9_hz100 matmult_inst.spi_inst.mosi_data_spi\[0\] _0024_ VGND VGND
+ VPWR VPWR matmult_inst.spi_inst.mosi_data_sync\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_39_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3174_ net127 net116 VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__and2_1
XFILLER_54_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2125_ net257 net231 net232 net255 VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__a22o_1
X_2056_ _0852_ net149 VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_52_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2958_ net334 net87 net38 VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1909_ _0538_ _0777_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__and2_1
X_2889_ _0541_ _0544_ net153 VGND VGND VPWR VPWR _1575_ sky130_fd_sc_hd__o21ai_1
XFILLER_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput4 net4 VGND VGND VPWR VPWR miso sky130_fd_sc_hd__buf_2
XFILLER_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2812_ _1516_ _1524_ VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__nor2_1
X_2743_ net259 net389 net95 VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__mux2_1
X_2674_ _1415_ _1416_ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__xnor2_1
X_1625_ matmult_inst.fsm_inst.count\[2\] matmult_inst.fsm_inst.count\[3\] VGND VGND
+ VPWR VPWR _0544_ sky130_fd_sc_hd__or2_1
XFILLER_39_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3226_ clknet_leaf_7_hz100 net306 VGND VGND VPWR VPWR matmult_inst.fsm_inst.alu_result\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3157_ net133 net122 VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_65_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2108_ matmult_inst.alu_inst.b1_reg\[0\] net247 VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__nand2_1
X_3088_ net363 net71 net26 VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__mux2_1
XFILLER_35_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2039_ _0840_ _0841_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__or2_1
XFILLER_52_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold360 matmult_inst.spi_inst.current_state VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2390_ _1160_ net544 _1161_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3011_ net492 net72 net33 VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__mux2_1
Xwire16 _1451_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_62_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2726_ net47 _1467_ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__nand2_1
X_2657_ _1400_ _1401_ VGND VGND VPWR VPWR _1402_ sky130_fd_sc_hd__and2_1
X_1608_ net654 VGND VGND VPWR VPWR matmult_inst.fsm_inst.tx_ready sky130_fd_sc_hd__inv_2
X_2588_ _1331_ _1332_ net59 VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__o21a_1
Xfanout114 _0801_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_4
Xfanout136 _0546_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout125 net126 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout169 _0568_ VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__buf_2
X_3209_ net290 VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__inv_2
XFILLER_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold190 matmult_inst.mem_inst.mem0\[4\] VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1890_ matmult_inst.fsm_inst.state\[4\] _0547_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_31_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3560_ clknet_leaf_23_hz100 _0420_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA1\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2511_ _1257_ _1258_ _1232_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__a21o_1
X_3491_ clknet_leaf_8_hz100 _0351_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem1\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2442_ _1178_ _1191_ _1192_ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__nand3_1
XFILLER_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2373_ _1156_ net426 net108 VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__mux2_1
XFILLER_68_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2709_ _1424_ _1429_ _1425_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__o21a_1
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2991_ net453 net73 net35 VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1942_ matmult_inst.spi_inst.tx_reg_sys\[8\] matmult_inst.spi_inst.miso_shifter\[7\]
+ net275 VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__mux2_1
X_1873_ net281 matmult_inst.mem_inst.mem0\[0\] matmult_inst.mem_inst.matrixB0\[0\]
+ net285 VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__a22o_1
X_3612_ clknet_leaf_17_hz100 _0472_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB0\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3543_ clknet_leaf_25_hz100 _0403_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA0\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3474_ clknet_leaf_15_hz100 _0334_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem0\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_2425_ net225 net213 net215 net223 VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__a22oi_1
XFILLER_69_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2356_ net267 _0541_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__nor2_1
XFILLER_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2287_ _1080_ _1081_ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__nand2_1
XFILLER_37_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire153 _0767_ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__buf_1
XFILLER_50_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2210_ _1002_ _1004_ _1005_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__or3_1
XFILLER_78_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3190_ net131 net121 VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__and2_1
X_2141_ net251 net236 net234 net253 VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__a22oi_2
XFILLER_81_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2072_ _0847_ net148 VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2974_ net312 net71 net38 VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__mux2_1
X_1925_ net287 _0785_ _0789_ _0792_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__a211o_1
X_1856_ net277 _0723_ _0726_ net282 VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__a22o_1
X_1787_ matmult_inst.mem_inst.matrixA2\[8\] net191 net183 matmult_inst.mem_inst.matrixA1\[8\]
+ _0665_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__a221o_1
X_3526_ clknet_leaf_8_hz100 _0386_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem3\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3457_ clknet_leaf_29_hz100 _0317_ VGND VGND VPWR VPWR matmult_inst.alu_inst.b0_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3388_ clknet_leaf_6_hz100 _0250_ VGND VGND VPWR VPWR matmult_inst.alu_inst.col1\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2408_ _1158_ net384 net63 VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__mux2_1
X_2339_ _1096_ _1119_ _1102_ net230 net245 VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__o2111ai_2
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold50 matmult_inst.mem_inst.mem3\[2\] VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 matmult_inst.mem_inst.matrixA0\[9\] VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 matmult_inst.alu_inst.row1\[3\] VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 matmult_inst.mem_inst.matrixB2\[8\] VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 matmult_inst.alu_inst.row1\[6\] VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_18_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1710_ matmult_inst.mem_inst.matrixA3\[15\] net198 _0595_ VGND VGND VPWR VPWR _0596_
+ sky130_fd_sc_hd__a21o_1
X_2690_ _1432_ _1433_ VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__nand2b_1
X_1641_ matmult_inst.spi_inst.rx_bit_count\[1\] _0557_ VGND VGND VPWR VPWR _0558_
+ sky130_fd_sc_hd__and2_2
XFILLER_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3311_ clknet_leaf_19_hz100 _0181_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB3\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_3242_ clknet_leaf_7_hz100 net603 VGND VGND VPWR VPWR matmult_inst.fsm_inst.alu_result\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_3173_ net127 net116 VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__and2_1
X_2124_ _0900_ net69 _0901_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__o21ba_1
X_2055_ _0853_ _0856_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_13_hz100 clknet_2_3__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_13_hz100
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2957_ net277 net198 net88 VGND VGND VPWR VPWR _1586_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_60_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2888_ _1574_ matmult_inst.fsm_inst.count\[0\] _1571_ VGND VGND VPWR VPWR _0324_
+ sky130_fd_sc_hd__mux2_1
X_1908_ matmult_inst.fsm_inst.state\[4\] _0536_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_28_hz100 clknet_2_0__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_28_hz100
+ sky130_fd_sc_hd__clkbuf_8
X_1839_ matmult_inst.mem_inst.matrixA2\[3\] net187 net179 matmult_inst.mem_inst.matrixA1\[3\]
+ _0712_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__a221o_1
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3509_ clknet_leaf_16_hz100 _0369_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem2\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput5 net5 VGND VGND VPWR VPWR ready sky130_fd_sc_hd__buf_2
XFILLER_56_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2811_ _1504_ _1509_ _1512_ _1517_ _1510_ VGND VGND VPWR VPWR _1524_ sky130_fd_sc_hd__o311a_1
X_2742_ matmult_inst.alu_inst.state\[0\] matmult_inst.alu_inst.state\[1\] _0778_ _0752_
+ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__nor4b_1
XFILLER_31_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2673_ _1414_ _1416_ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__nor2_1
X_1624_ matmult_inst.fsm_inst.count\[2\] matmult_inst.fsm_inst.count\[3\] VGND VGND
+ VPWR VPWR _0543_ sky130_fd_sc_hd__nor2_1
X_3225_ clknet_leaf_7_hz100 _0123_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.alu_result\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3156_ net127 net116 VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__and2_1
X_3087_ net529 _0819_ net25 VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2107_ net240 net242 matmult_inst.alu_inst.a1_reg\[4\] net249 VGND VGND VPWR VPWR
+ _0907_ sky130_fd_sc_hd__and4_1
X_2038_ _0828_ _0837_ _0839_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_37_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold350 matmult_inst.alu_inst.adder_inst.r3.fa3.a VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 matmult_inst.spi_inst.current_state VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3010_ net552 net73 net33 VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__mux2_1
XFILLER_36_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2725_ _1443_ net103 _1444_ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__o21bai_2
X_2656_ _1387_ _1398_ _1399_ VGND VGND VPWR VPWR _1401_ sky130_fd_sc_hd__nand3_1
X_2587_ net59 _1331_ _1332_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__nor3_1
Xfanout115 _0565_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_4
Xfanout159 net160 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_4
X_3208_ net290 VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__inv_2
XFILLER_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3139_ net129 net119 VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__and2_1
XFILLER_27_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold180 matmult_inst.mem_inst.matrixA0\[13\] VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold191 matmult_inst.mem_inst.mem0\[3\] VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_2__f_hz100 clknet_0_hz100 VGND VGND VPWR VPWR clknet_2_2__leaf_hz100 sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_31_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2510_ _1257_ _1258_ _1232_ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__a21oi_1
X_3490_ clknet_leaf_8_hz100 _0350_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem1\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2441_ net228 net207 net210 net226 VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__a22o_1
X_2372_ _0721_ net166 VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__and2_2
XFILLER_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2708_ _1445_ _1450_ VGND VGND VPWR VPWR _1451_ sky130_fd_sc_hd__xnor2_1
X_2639_ net224 net204 _1347_ _1349_ VGND VGND VPWR VPWR _1384_ sky130_fd_sc_hd__a22o_1
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_74 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2990_ net474 _0817_ net35 VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1941_ matmult_inst.spi_inst.tx_reg_sys\[7\] matmult_inst.spi_inst.miso_shifter\[6\]
+ net275 VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__mux2_1
X_1872_ matmult_inst.mem_inst.mem2\[0\] net189 net181 matmult_inst.mem_inst.mem1\[0\]
+ _0742_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__a221o_1
X_3611_ clknet_leaf_14_hz100 _0471_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA3\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_3542_ clknet_leaf_25_hz100 _0402_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixA0\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3473_ clknet_leaf_7_hz100 _0333_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem0\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_2424_ _1175_ _1176_ net645 net174 VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__a2bb2o_1
X_2355_ net267 net165 net166 matmult_inst.fsm_inst.state\[2\] VGND VGND VPWR VPWR
+ _1144_ sky130_fd_sc_hd__o211a_1
X_2286_ _1057_ _1079_ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__or2_1
XFILLER_64_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire110 _1150_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_1
Xwire143 _1201_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
Xwire176 _0787_ VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__buf_1
XFILLER_3_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2140_ _0905_ _0908_ _0907_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__o21ba_1
XFILLER_66_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2071_ _0870_ _0871_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2973_ net345 net72 net37 VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__mux2_1
X_1924_ _0753_ _0760_ _0790_ _0791_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__or4_1
X_1855_ matmult_inst.mem_inst.matrixA2\[2\] net187 net179 matmult_inst.mem_inst.matrixA1\[2\]
+ _0727_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_12_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1786_ net273 net265 matmult_inst.mem_inst.matrixA3\[8\] VGND VGND VPWR VPWR _0665_
+ sky130_fd_sc_hd__and3_1
X_3525_ clknet_leaf_17_hz100 _0385_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem3\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3456_ clknet_leaf_29_hz100 _0316_ VGND VGND VPWR VPWR matmult_inst.alu_inst.b0_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3387_ clknet_leaf_2_hz100 _0249_ VGND VGND VPWR VPWR matmult_inst.alu_inst.col1\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2407_ _1157_ net400 net64 VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__mux2_1
XFILLER_69_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2338_ net230 net245 _1102_ _1119_ _1096_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__a311o_1
X_2269_ _1029_ _1064_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__and2_1
XFILLER_25_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold40 matmult_inst.mem_inst.mem3\[0\] VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 matmult_inst.mem_inst.mem3\[15\] VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 matmult_inst.alu_inst.col0\[1\] VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 matmult_inst.mem_inst.mem1\[16\] VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 matmult_inst.alu_inst.row1\[0\] VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 matmult_inst.mem_inst.matrixB1\[8\] VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1640_ matmult_inst.spi_inst.rx_bit_count\[3\] matmult_inst.spi_inst.rx_bit_count\[0\]
+ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_9_hz100 clknet_2_3__leaf_hz100 VGND VGND VPWR VPWR clknet_leaf_9_hz100
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3310_ clknet_leaf_17_hz100 _0180_ VGND VGND VPWR VPWR matmult_inst.mem_inst.matrixB3\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3241_ clknet_leaf_26_hz100 net309 VGND VGND VPWR VPWR matmult_inst.fsm_inst.alu_result\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3172_ net127 net116 VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__and2_1
X_2123_ net601 _0922_ net162 VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__mux2_1
XFILLER_26_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2054_ _0854_ _0855_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__nand2b_1
XFILLER_81_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2956_ net374 net70 net40 VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__mux2_1
X_2887_ net152 _0771_ _1572_ _1573_ _1604_ VGND VGND VPWR VPWR _1574_ sky130_fd_sc_hd__o221a_1
X_1907_ net166 _0775_ _0773_ _0769_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_60_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1838_ net270 net262 matmult_inst.mem_inst.matrixA3\[3\] VGND VGND VPWR VPWR _0712_
+ sky130_fd_sc_hd__and3_1
X_1769_ net284 _0644_ _0649_ _0642_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__a211o_1
X_3508_ clknet_leaf_8_hz100 _0368_ VGND VGND VPWR VPWR matmult_inst.mem_inst.mem2\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3439_ clknet_leaf_7_hz100 _0299_ VGND VGND VPWR VPWR matmult_inst.alu_inst.out\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2810_ _1521_ _1522_ VGND VGND VPWR VPWR _1523_ sky130_fd_sc_hd__nand2b_1
X_2741_ net541 net175 VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__and2_1
X_2672_ _1390_ _1392_ _1391_ VGND VGND VPWR VPWR _1416_ sky130_fd_sc_hd__o21ba_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1623_ matmult_inst.fsm_inst.count\[1\] matmult_inst.fsm_inst.count\[0\] VGND VGND
+ VPWR VPWR _0542_ sky130_fd_sc_hd__and2_1
X_3224_ clknet_leaf_25_hz100 _0002_ VGND VGND VPWR VPWR matmult_inst.fsm_inst.sel\[2\]
+ sky130_fd_sc_hd__dfxtp_1
.ends


* NGSPICE file created from pwm_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt pwm_wrapper CLK VGND VPWR addr[0] addr[10] addr[11] addr[12] addr[13] addr[14]
+ addr[15] addr[16] addr[17] addr[18] addr[19] addr[1] addr[20] addr[21] addr[22]
+ addr[23] addr[24] addr[25] addr[26] addr[27] addr[28] addr[29] addr[2] addr[30]
+ addr[31] addr[3] addr[4] addr[5] addr[6] addr[7] addr[8] addr[9] error nRST pwm_out[0]
+ pwm_out[1] rdata[0] rdata[10] rdata[11] rdata[12] rdata[13] rdata[14] rdata[15]
+ rdata[16] rdata[17] rdata[18] rdata[19] rdata[1] rdata[20] rdata[21] rdata[22] rdata[23]
+ rdata[24] rdata[25] rdata[26] rdata[27] rdata[28] rdata[29] rdata[2] rdata[30] rdata[31]
+ rdata[3] rdata[4] rdata[5] rdata[6] rdata[7] rdata[8] rdata[9] ren request_stall
+ strobe[0] strobe[1] strobe[2] strobe[3] wdata[0] wdata[10] wdata[11] wdata[12] wdata[13]
+ wdata[14] wdata[15] wdata[16] wdata[17] wdata[18] wdata[19] wdata[1] wdata[20] wdata[21]
+ wdata[22] wdata[23] wdata[24] wdata[25] wdata[26] wdata[27] wdata[28] wdata[29]
+ wdata[2] wdata[30] wdata[31] wdata[3] wdata[4] wdata[5] wdata[6] wdata[7] wdata[8]
+ wdata[9] wen
XFILLER_0_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3155_ _0759_ _0824_ _0929_ _0990_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__a31oi_4
X_3086_ net106 _0919_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__nand2_1
X_2106_ net340 net56 _1546_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2037_ net285 net60 net87 VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3988_ net183 VGND VGND VPWR VPWR rdata[11] sky130_fd_sc_hd__buf_2
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2939_ _0516_ _0538_ _0546_ _0513_ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__and4b_1
XFILLER_0_72_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2954__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout75_A _1540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3196__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3370__A1 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_6_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_6_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_47_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3911_ clknet_leaf_4_CLK _0237_ net151 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[60\]
+ sky130_fd_sc_hd__dfrtp_2
X_3842_ clknet_leaf_5_CLK _0168_ net152 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3773_ clknet_leaf_10_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[20\]
+ net158 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_14_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2722__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2724_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[43\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[11\]
+ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2655_ _0489_ _0490_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_74_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2586_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[10\]
+ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__xor2_1
Xfanout127 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[3\] VGND VGND VPWR VPWR net127
+ sky130_fd_sc_hd__buf_2
Xfanout116 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[6\] VGND VGND VPWR VPWR net116
+ sky130_fd_sc_hd__buf_2
Xfanout138 net33 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_2
Xfanout105 _1535_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__buf_2
Xfanout149 net33 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_4
X_3207_ _1027_ _1041_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3138_ _1610_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[41\] VGND VGND VPWR
+ VPWR _0974_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout165_X net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3069_ _0898_ _0901_ _0904_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2124__S net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout78_X net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2034__S net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1873__S net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2440_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\]
+ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2371_ _1769_ _1770_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[23\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3825_ clknet_leaf_18_CLK _0151_ net167 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_15_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3756_ clknet_leaf_23_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[3\] net161
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3987__182 VGND VGND VPWR VPWR _3987__182/HI net182 sky130_fd_sc_hd__conb_1
X_2707_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[38\]
+ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3687_ clknet_leaf_33_CLK _0047_ net139 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2638_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[53\] _0473_ VGND VGND VPWR
+ VPWR _0474_ sky130_fd_sc_hd__nor2_1
X_2569_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\] _0407_ net69 VGND VGND VPWR
+ VPWR _0410_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2119__S net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1958__S net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2362__B myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_80_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3325__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input55_A wdata[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1887__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2029__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1868__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1940_ net208 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[42\] net101 VGND
+ VGND VPWR VPWR _0089_ sky130_fd_sc_hd__mux2_1
XANTENNA__2064__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1871_ net214 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] net105 VGND
+ VGND VPWR VPWR _0023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3610_ _1387_ _1388_ _1444_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__and3b_1
XFILLER_0_71_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3541_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] _1372_ _1375_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\]
+ VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3472_ _1080_ _1083_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2423_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] _1768_ VGND VGND VPWR
+ VPWR _0293_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_71_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2354_ net121 _1756_ _1758_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[18\]
+ sky130_fd_sc_hd__o21a_1
X_2285_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[28\]
+ VGND VGND VPWR VPWR _1707_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2055__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3808_ clknet_leaf_6_CLK _0134_ net155 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3739_ clknet_leaf_0_CLK _0099_ net135 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1869__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2046__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input58_X net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2548__A _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2070_ net285 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[36\] net92 VGND
+ VGND VPWR VPWR _0213_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_11_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2037__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2972_ _0805_ _0806_ _0807_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1923_ net304 net52 net77 VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_26_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1854_ net257 net51 net81 VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3524_ _1135_ _1358_ VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3455_ _1080_ _1081_ VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2406_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] _1722_ _1728_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\]
+ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__a2bb2o_1
X_3386_ _1011_ _1220_ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__xnor2_1
X_2337_ _1712_ _1745_ _1746_ VGND VGND VPWR VPWR _1747_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2268_ _1554_ net125 _1562_ net123 _1689_ VGND VGND VPWR VPWR _1690_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_68_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4007_ net202 VGND VGND VPWR VPWR rdata[30] sky130_fd_sc_hd__buf_2
X_2199_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[24\] VGND VGND VPWR VPWR
+ _1621_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1971__S net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold41 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[0\] VGND VGND VPWR VPWR net245
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[26\] VGND VGND VPWR VPWR net234
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold74 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[5\] VGND VGND VPWR VPWR net278
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[49\] VGND VGND VPWR VPWR net267
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[2\] VGND VGND VPWR VPWR net256
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[21\] VGND VGND VPWR VPWR net300
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[39\] VGND VGND VPWR VPWR net289
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input18_A addr[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2267__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_85_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2019__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2042__S net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1881__S net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3240_ _1072_ _1074_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3171_ _1004_ _1005_ _0999_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__a21o_1
X_2122_ net206 net40 net81 VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2053_ net276 net46 net86 VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2955_ _0493_ _0497_ _0762_ _0789_ _0494_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__o221a_1
X_2886_ _0677_ _0720_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__nor2_1
X_1906_ net216 net65 net80 VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__mux2_1
X_1837_ net13 net16 net15 net18 VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_77_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3507_ _1331_ _1333_ _1340_ _1341_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_9_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3438_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[24\] _1268_ _1271_ _1272_ VGND VGND
+ VPWR VPWR _1273_ sky130_fd_sc_hd__o211a_1
X_3369_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[1\] _1200_ _1203_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\]
+ _1202_ VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__o221a_1
XFILLER_0_95_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1966__S net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2037__S net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1876__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2412__B2 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2740_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[17\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[49\]
+ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2671_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[42\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\]
+ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_41_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3223_ _1053_ _1057_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__nand2_1
X_3154_ _0935_ _0939_ _0989_ _0937_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__a31oi_2
X_2105_ net317 net45 _1546_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__mux2_1
X_3085_ net106 _0919_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__or2_1
X_2036_ net258 net59 net87 VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3671__RESET_B net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3567__A _1560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3987_ net182 VGND VGND VPWR VPWR rdata[10] sky130_fd_sc_hd__buf_2
XFILLER_0_43_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_2__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_2_2__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_2938_ _0524_ _0688_ _0771_ _0773_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2954__A2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2869_ _0552_ _0555_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2646__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2642__A1 _1621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input40_X net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2556__A myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3910_ clknet_leaf_4_CLK _0236_ net152 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[59\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_86_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3841_ clknet_leaf_6_CLK _0167_ net155 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_3772_ clknet_leaf_10_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[19\]
+ net158 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__2291__A myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_2723_ _0507_ _0558_ _0508_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__a21oi_1
X_2654_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\]
+ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__nand2b_1
X_2585_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[0\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[0\]
+ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_74_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout117 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[30\] VGND VGND VPWR VPWR net117
+ sky130_fd_sc_hd__clkbuf_4
Xfanout106 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[27\] VGND VGND VPWR VPWR net106
+ sky130_fd_sc_hd__buf_2
Xfanout128 net132 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_4
Xfanout139 net141 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_4
X_3206_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] _1667_ _1032_ _1039_
+ _1029_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__a221o_2
X_3137_ _1607_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[39\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[38\]
+ _1605_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3068_ _0847_ _0902_ _0903_ _0849_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__or4b_1
XANTENNA_fanout158_X net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2019_ net300 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] net95 VGND
+ VGND VPWR VPWR _0165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_470 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1832__X _1521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2312__B1 _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2615__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2050__S net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2370_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\] _1767_ _1713_ VGND VGND VPWR
+ VPWR _1770_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3824_ clknet_leaf_21_CLK _0150_ net162 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_82_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3755_ clknet_leaf_12_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[2\] net159
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_15_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3686_ clknet_leaf_40_CLK _0046_ net130 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_mod\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2706_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[38\]
+ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2637_ _0471_ _0472_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__and2b_2
XFILLER_0_42_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2568_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\] _0407_ VGND VGND VPWR VPWR
+ _0409_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2499_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\] _0358_ VGND VGND VPWR VPWR _0364_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2196__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1974__S net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout90_X net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3774__RESET_B net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input48_A wdata[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3703__RESET_B net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2045__S net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1870_ net236 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\] net105 VGND
+ VGND VPWR VPWR _0022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3013__A1 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__1884__S net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3540_ _1365_ _1374_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3471_ _1299_ _1301_ _1305_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__a21o_2
XFILLER_0_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2422_ _0277_ _0278_ _0290_ _0291_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_71_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2353_ net121 _1756_ net72 VGND VGND VPWR VPWR _1758_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2284_ _1565_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[15\] _1590_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\]
+ VGND VGND VPWR VPWR _1706_ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2827__A1 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3807_ clknet_leaf_6_CLK _0133_ net155 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1999_ net235 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] net96 VGND VGND
+ VPWR VPWR _0145_ sky130_fd_sc_hd__mux2_1
X_3738_ clknet_leaf_1_CLK _0098_ net135 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\]
+ sky130_fd_sc_hd__dfrtp_2
X_3669_ clknet_leaf_39_CLK _0029_ net131 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2818__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1969__S net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3482__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1879__S net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2971_ _0604_ _0608_ _0804_ _0606_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1922_ net310 net51 net77 VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1853_ net207 net50 net82 VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3523_ _1131_ _1347_ VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__nand2_1
X_3454_ _1069_ _1070_ _1288_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__or3_1
X_2405_ _1551_ _1719_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__xnor2_1
X_3385_ _1004_ _1115_ _1118_ _1006_ VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__a31o_1
X_2336_ net123 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\] _1742_ VGND VGND VPWR
+ VPWR _1746_ sky130_fd_sc_hd__and3_1
X_2267_ _1549_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[0\] _1570_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\]
+ VGND VGND VPWR VPWR _1689_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_68_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4006_ net201 VGND VGND VPWR VPWR rdata[29] sky130_fd_sc_hd__buf_2
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2198_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] VGND VGND VPWR VPWR
+ _1620_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout98_A _1538_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold31 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[1\] VGND VGND VPWR VPWR net235
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[34\] VGND VGND VPWR VPWR net224
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[14\] VGND VGND VPWR VPWR net246
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[25\] VGND VGND VPWR VPWR net257
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[37\] VGND VGND VPWR VPWR net268
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[8\] VGND VGND VPWR VPWR net301
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold86 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[53\] VGND VGND VPWR VPWR net290
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[30\] VGND VGND VPWR VPWR net279
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2384__A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2559__A myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_3170_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[53\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\]
+ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__and2b_1
X_2121_ net246 net39 net83 VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__mux2_1
X_2052_ net328 net44 net86 VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2294__A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2954_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\]
+ _0788_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1905_ net239 net64 net79 VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__mux2_1
X_2885_ net112 _0679_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1836_ net17 net20 net19 net22 VGND VGND VPWR VPWR _1524_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3506_ net117 _1330_ _1332_ _1671_ _1329_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__a311o_1
XANTENNA_fanout100_A _1538_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3437_ net119 _1266_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__xnor2_1
X_3368_ _1032_ _1039_ VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__xnor2_1
X_2319_ net125 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[7\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[8\]
+ _1727_ VGND VGND VPWR VPWR _1734_ sky130_fd_sc_hd__and4_1
XFILLER_0_57_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3299_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[58\]
+ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1982__S net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_10_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input30_A addr[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1999__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2053__S net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2670_ _0505_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1892__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1923__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3222_ _1027_ _1041_ _1056_ _1055_ _1048_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__a32oi_4
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3153_ _0983_ _0988_ _0960_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__o21ai_1
X_2104_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable net34 _1546_ VGND VGND
+ VPWR VPWR _0245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3084_ net106 _0919_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2035_ net255 net56 net87 VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__mux2_1
XANTENNA__2100__A1 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_99_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3986_ net181 VGND VGND VPWR VPWR rdata[9] sky130_fd_sc_hd__buf_2
XANTENNA__2752__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout148_A net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2937_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[3\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[35\]
+ _0688_ _0768_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__a31o_1
XFILLER_0_94_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3640__RESET_B net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2868_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\] _0702_ VGND VGND VPWR VPWR _0704_
+ sky130_fd_sc_hd__nand2_1
X_1819_ _1594_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[63\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[62\]
+ _1593_ VGND VGND VPWR VPWR _1508_ sky130_fd_sc_hd__a2bb2o_1
X_2799_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[62\]
+ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1914__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout103_X net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2199__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[24\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1977__S net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3799__RESET_B net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1905__A1 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input33_X net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2048__S net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1887__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3840_ clknet_leaf_6_CLK _0166_ net155 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\]
+ sky130_fd_sc_hd__dfrtp_4
X_3771_ clknet_leaf_10_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[18\]
+ net158 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2722_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[41\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\]
+ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_42_503 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2653_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\]
+ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__nand2b_2
X_2584_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[0\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[0\]
+ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_74_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout118 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[27\] VGND VGND VPWR VPWR net118
+ sky130_fd_sc_hd__buf_2
Xfanout129 net132 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_4
Xfanout107 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[21\] VGND VGND VPWR VPWR net107
+ sky130_fd_sc_hd__buf_2
X_3205_ _1032_ _1039_ _1029_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__a21oi_1
X_3136_ _1605_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[38\] _0965_ _0971_
+ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__a22o_1
X_3067_ net111 _0900_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__nor2_1
X_2018_ net270 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] net95 VGND
+ VGND VPWR VPWR _0164_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_555 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3969_ clknet_leaf_24_CLK _0261_ net145 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout80_A _1537_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3909__RESET_B net154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3398__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3823_ clknet_leaf_22_CLK _0149_ net162 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_62_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3754_ clknet_leaf_23_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[1\] net160
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_15_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3685_ clknet_leaf_40_CLK _0045_ net130 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\]
+ sky130_fd_sc_hd__dfrtp_2
X_2705_ _0519_ _0533_ _0537_ _0539_ _0540_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__a311o_1
XFILLER_0_42_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2636_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\]
+ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__nand2_1
X_2567_ _0407_ _0408_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[28\]
+ sky130_fd_sc_hd__nor2_1
X_2498_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\] _0358_ VGND VGND VPWR VPWR _0363_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout170_X net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3119_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] _1636_ _1637_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[22\]
+ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_591 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2533__A1 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__1990__S net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout83_X net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Left_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2061__S net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3470_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[40\]
+ _1303_ _1304_ VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2421_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[20\]
+ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_71_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2352_ _1756_ _1757_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[17\]
+ sky130_fd_sc_hd__nor2_1
X_2283_ _1553_ net126 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] _1563_
+ VGND VGND VPWR VPWR _1705_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_63_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_72_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3806_ clknet_leaf_7_CLK _0132_ net156 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2760__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_1998_ net245 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[0\] net96 VGND VGND
+ VPWR VPWR _0144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3737_ clknet_leaf_1_CLK _0097_ net138 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3668_ clknet_leaf_34_CLK _0028_ net139 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_30_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3599_ _1425_ _1426_ _1432_ _1433_ VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2619_ _1625_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[26\] VGND VGND VPWR
+ VPWR _0456_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_81_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2654__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_90_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1985__S net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2451__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input60_A wdata[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3467__C1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3977__172 VGND VGND VPWR VPWR _3977__172/HI net172 sky130_fd_sc_hd__conb_1
XFILLER_0_88_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2056__S net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2970_ _0595_ _0599_ _0596_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1921_ net315 net50 net78 VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1852_ net312 net49 net82 VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3522_ _1347_ _1356_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3453_ _1061_ _1065_ VGND VGND VPWR VPWR _1288_ sky130_fd_sc_hd__nand2_1
X_2404_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] _1716_ _1725_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\]
+ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__o2bb2a_1
X_3384_ _1216_ _1217_ _1218_ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__a21o_1
X_2335_ net123 _1742_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\] VGND VGND VPWR
+ VPWR _1745_ sky130_fd_sc_hd__a21oi_1
X_2266_ _1554_ net125 _1561_ net124 _1687_ VGND VGND VPWR VPWR _1688_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_68_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4005_ net200 VGND VGND VPWR VPWR rdata[28] sky130_fd_sc_hd__buf_2
X_2197_ net109 VGND VGND VPWR VPWR _1619_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_38_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_38_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold32 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[8\] VGND VGND VPWR VPWR net236
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[9\] VGND VGND VPWR VPWR net214
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[3\] VGND VGND VPWR VPWR net225
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[48\] VGND VGND VPWR VPWR net269
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[33\] VGND VGND VPWR VPWR net247
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[35\] VGND VGND VPWR VPWR net258
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold76 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[26\] VGND VGND VPWR VPWR net280
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[32\] VGND VGND VPWR VPWR net291
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold98 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[51\] VGND VGND VPWR VPWR net302
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_29_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_29_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input63_X net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2120_ net227 net38 net84 VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__mux2_1
X_2051_ net334 net43 net86 VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2953_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\]
+ _0788_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1904_ net289 net63 net80 VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2884_ _1613_ _0673_ _0676_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__and3_1
X_1835_ net21 net25 net24 VGND VGND VPWR VPWR _1523_ sky130_fd_sc_hd__or3_1
XFILLER_0_72_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3505_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] _1338_ _1339_ VGND VGND VPWR
+ VPWR _1340_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3436_ net120 _1269_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3367_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[1\] _1200_ _1201_ _1037_ VGND VGND
+ VPWR VPWR _1202_ sky130_fd_sc_hd__a211o_1
X_2318_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[8\] _1731_ VGND VGND VPWR VPWR _1733_
+ sky130_fd_sc_hd__nor2_1
X_3298_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[58\]
+ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__nor2_1
XANTENNA__2485__A _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2249_ myPWM.g_pwm_channel\[1\].CHANNEL.alignment VGND VGND VPWR VPWR _1671_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input23_A addr[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3221_ _1025_ _1045_ _1055_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_9_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_9_CLK sky130_fd_sc_hd__clkbuf_8
X_3152_ _0955_ _0959_ _0984_ _0987_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__or4b_1
X_2103_ net12 net1 net23 _1542_ VGND VGND VPWR VPWR _1546_ sky130_fd_sc_hd__and4bb_1
X_3083_ _0597_ _0918_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__xnor2_1
X_2034_ net247 net45 net87 VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3985_ net180 VGND VGND VPWR VPWR rdata[8] sky130_fd_sc_hd__buf_2
X_2936_ _0524_ _0771_ _0523_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2867_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\] _0702_ VGND VGND VPWR VPWR _0703_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1818_ _1581_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[56\] _1502_ _1504_
+ _1506_ VGND VGND VPWR VPWR _1507_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2798_ _0619_ _0623_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3419_ _1247_ _1250_ _1243_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1850__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3768__RESET_B net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1993__S net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4002__197 VGND VGND VPWR VPWR _4002__197/HI net197 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_19_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3770_ clknet_leaf_9_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[17\] net158
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_66_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2064__S net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2721_ _0499_ _0506_ _0509_ _0555_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2652_ _0485_ _0486_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__or2_2
X_2583_ _1595_ _1633_ _0420_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[0\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout119 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[26\] VGND VGND VPWR VPWR net119
+ sky130_fd_sc_hd__clkbuf_4
Xfanout108 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR net108
+ sky130_fd_sc_hd__buf_2
X_3204_ _1035_ _1036_ _1038_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__a21o_1
X_3135_ _1603_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[36\] _0968_ _0969_
+ _0970_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3066_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[16\] _0848_ VGND VGND VPWR VPWR
+ _0902_ sky130_fd_sc_hd__nor2_1
X_2017_ net287 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] net95 VGND
+ VGND VPWR VPWR _0163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2763__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3968_ clknet_leaf_24_CLK _0260_ net145 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3585__A1 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2919_ _0630_ _0633_ _0641_ _0642_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__and4_1
XFILLER_0_18_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3899_ clknet_leaf_9_CLK _0225_ net158 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__3861__RESET_B net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_24_CLK_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1899__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_39_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout73_A _1540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1988__S net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2673__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3949__RESET_B net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3000__C _0798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2059__S net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1898__S net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3822_ clknet_leaf_20_CLK _0148_ net164 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3753_ clknet_leaf_12_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[0\] net161
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3684_ clknet_leaf_41_CLK _0044_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\]
+ sky130_fd_sc_hd__dfrtp_4
X_2704_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[37\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\]
+ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__and2b_1
XFILLER_0_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2635_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\]
+ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2566_ net69 _0406_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__nand2_1
XANTENNA__2758__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2497_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[3\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[4\]
+ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\] _0354_ VGND VGND VPWR VPWR _0362_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3118_ _1624_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[57\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[56\]
+ _1622_ _0953_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__o221a_1
XFILLER_0_97_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3994__189 VGND VGND VPWR VPWR _3994__189/HI net189 sky130_fd_sc_hd__conb_1
X_3049_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[4\] _0875_ _0877_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[3\]
+ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__o22a_1
XANTENNA__2058__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3825__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout76_X net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_100_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2049__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout90 _1544_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2420_ _1566_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[16\] _0288_ _0289_
+ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2351_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] _1754_ _1713_ VGND VGND VPWR
+ VPWR _1757_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_71_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2282_ _1553_ net126 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\] _1558_
+ _1703_ VGND VGND VPWR VPWR _1704_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3805_ clknet_leaf_7_CLK _0131_ net156 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1997_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.rollover_flag myPWM.g_pwm_channel\[1\].CHANNEL.data_mod\[0\]
+ VGND VGND VPWR VPWR _1541_ sky130_fd_sc_hd__nand2_2
X_3736_ clknet_leaf_2_CLK _0096_ net138 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3667_ clknet_leaf_24_CLK _0027_ net144 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_3598_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[10\] _1401_ _1404_ _1405_ _1398_
+ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__o2111a_1
X_2618_ _1630_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[30\] _0441_ _0442_
+ _0454_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_11_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2549_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] _0395_ VGND VGND VPWR VPWR
+ _0396_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2451__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1962__B1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input53_A wdata[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1920_ net314 net49 net78 VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1851_ net329 net48 net82 VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__mux2_1
XANTENNA__2072__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3521_ _1132_ _1282_ _1321_ VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__nand3_1
XFILLER_0_24_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3452_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\]
+ _1286_ VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__o21ai_2
X_3383_ net122 _1175_ _1176_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[14\] VGND VGND
+ VPWR VPWR _1218_ sky130_fd_sc_hd__a22o_1
X_2403_ _1570_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[19\] VGND VGND VPWR
+ VPWR _0273_ sky130_fd_sc_hd__xnor2_1
X_2334_ net123 _1742_ _1744_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[12\]
+ sky130_fd_sc_hd__o21a_1
X_2265_ _1561_ net124 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\] _1594_
+ VGND VGND VPWR VPWR _1687_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_68_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4004_ net199 VGND VGND VPWR VPWR rdata[27] sky130_fd_sc_hd__buf_2
X_2196_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] VGND VGND VPWR VPWR
+ _1618_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2771__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3719_ clknet_leaf_33_CLK _0079_ net139 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3107__A myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xhold22 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[18\] VGND VGND VPWR VPWR net226
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[11\] VGND VGND VPWR VPWR net215
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[43\] VGND VGND VPWR VPWR net259
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[24\] VGND VGND VPWR VPWR net237
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[40\] VGND VGND VPWR VPWR net248
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[44\] VGND VGND VPWR VPWR net303
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold66 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[20\] VGND VGND VPWR VPWR net270
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold77 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[63\] VGND VGND VPWR VPWR net281
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[62\] VGND VGND VPWR VPWR net292
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1996__S net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input56_X net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2856__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2050_ net277 net42 net86 VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2067__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2952_ _0486_ _0492_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__and2_1
X_1903_ net223 net62 net79 VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2883_ net113 _0678_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__or2_1
X_1834_ net317 _1521_ _1522_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.pwm_next
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2654__A_N myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3504_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] _1336_ _1337_ _1335_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[28\]
+ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__a32oi_1
XFILLER_0_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3435_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[24\] _1268_ _1269_ net120 VGND VGND
+ VPWR VPWR _1270_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3366_ _1035_ _1036_ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__nor2_1
XANTENNA__2351__B1 _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2317_ net71 _1731_ _1732_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[7\]
+ sky130_fd_sc_hd__nor3_1
X_3297_ _1130_ _1131_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__nand2_2
X_2248_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[33\] VGND VGND VPWR VPWR
+ _1670_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2179_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[3\] VGND VGND VPWR VPWR _1601_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2406__B2 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput67 net67 VGND VGND VPWR VPWR pwm_out[0] sky130_fd_sc_hd__buf_2
XANTENNA_input16_A addr[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4007__202 VGND VGND VPWR VPWR _4007__202/HI net202 sky130_fd_sc_hd__conb_1
XFILLER_0_22_443 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3220_ _1021_ _1054_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__nor2_1
XANTENNA__2586__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3151_ _0942_ _0951_ _0952_ _0986_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__and4b_1
X_2102_ _1547_ net337 net73 VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__a21o_1
X_3082_ _0600_ _0607_ _0913_ _0599_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__a31o_1
X_2033_ net291 net34 net87 VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__mux2_1
X_3984_ net179 VGND VGND VPWR VPWR rdata[7] sky130_fd_sc_hd__buf_2
X_2935_ _0526_ _0770_ _0527_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2866_ _0513_ _0701_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__xor2_1
XFILLER_0_72_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1817_ _1585_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[58\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[57\]
+ _1583_ _1505_ VGND VGND VPWR VPWR _1506_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2797_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[31\] _0632_ VGND VGND VPWR VPWR
+ _0633_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3418_ _1219_ _1236_ _1237_ _1252_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__and4_1
X_3349_ _1075_ _1183_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__xnor2_1
XANTENNA_input8_A addr[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3828__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1846__Y _1534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3030__A net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2720_ _0512_ _0549_ _0551_ _0555_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2651_ _0485_ _0486_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2080__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2582_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[0\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.count_enable
+ _0349_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_74_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout109 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR net109
+ sky130_fd_sc_hd__buf_2
XFILLER_0_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3203_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[34\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[2\]
+ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__and2b_1
X_3134_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[37\]
+ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__and2b_1
X_3065_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[14\] _0853_ _0900_ net111 VGND VGND
+ VPWR VPWR _0901_ sky130_fd_sc_hd__a22oi_1
X_2016_ net226 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] net95 VGND
+ VGND VPWR VPWR _0162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout153_A net154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3967_ clknet_leaf_25_CLK _0259_ net147 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2918_ _0744_ _0747_ _0749_ net106 _0745_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__a221o_1
X_3898_ clknet_leaf_12_CLK _0224_ net159 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[47\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2849_ _0519_ _0533_ _0537_ _0540_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold130 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[50\] VGND VGND VPWR VPWR net334
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2075__S net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3821_ clknet_leaf_22_CLK _0147_ net162 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3752_ clknet_leaf_2_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.rollover_flag_c net153
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.rollover_flag sky130_fd_sc_hd__dfrtp_1
X_3683_ clknet_leaf_42_CLK _0043_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\]
+ sky130_fd_sc_hd__dfrtp_4
X_2703_ _1604_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[38\] VGND VGND VPWR
+ VPWR _0539_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2634_ _0468_ _0469_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__nand2_2
XFILLER_0_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2565_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[27\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\]
+ _0403_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2496_ _0361_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[4\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3117_ _1627_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[59\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[58\]
+ _1626_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__o22a_1
X_3048_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[3\] _0877_ _0878_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[2\]
+ _0883_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1999__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3956__CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout91 _1544_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_2
XFILLER_0_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout80 _1537_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_2
XFILLER_0_64_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1980__A1 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2350_ net122 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[16\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\]
+ _1749_ VGND VGND VPWR VPWR _1756_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_71_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2281_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] _1559_ _1582_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[25\]
+ VGND VGND VPWR VPWR _1703_ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_23_CLK_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_38_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3804_ clknet_leaf_8_CLK _0130_ net157 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1996_ net309 net58 net73 VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3735_ clknet_leaf_37_CLK _0095_ net138 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[48\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3666_ clknet_leaf_24_CLK _0026_ net144 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__1971__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3597_ _1560_ _1400_ _1409_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[7\] _1427_
+ VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2617_ _0417_ _0443_ _0446_ _0453_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2548_ _0351_ _0394_ _0395_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[22\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__3661__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2479_ _0320_ _0325_ _0343_ _0347_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__or4_1
XFILLER_0_97_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3836__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload0 clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__2679__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input46_A wdata[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3467__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3933__RESET_B net144 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1850_ net327 net47 net82 VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3520_ net119 _1353_ _1354_ VGND VGND VPWR VPWR _1355_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_24_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3451_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\]
+ _1068_ _1285_ _1066_ VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__a221o_1
XANTENNA__2589__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3382_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[14\] _1176_ _1180_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\]
+ VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__o22a_1
X_2402_ _1555_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[7\] VGND VGND VPWR
+ VPWR _0272_ sky130_fd_sc_hd__xnor2_1
X_2333_ net123 _1742_ _1712_ VGND VGND VPWR VPWR _1744_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2264_ _1683_ _1684_ _1685_ _1682_ VGND VGND VPWR VPWR _1686_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4003_ net198 VGND VGND VPWR VPWR rdata[26] sky130_fd_sc_hd__buf_2
X_2195_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[17\] VGND VGND VPWR VPWR
+ _1617_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1979_ net316 net39 net75 VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1944__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3718_ clknet_leaf_41_CLK _0078_ net130 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3649_ clknet_leaf_43_CLK _0009_ net128 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold12 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[41\] VGND VGND VPWR VPWR net216
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[13\] VGND VGND VPWR VPWR net227
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[9\] VGND VGND VPWR VPWR net260
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[6\] VGND VGND VPWR VPWR net238
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[54\] VGND VGND VPWR VPWR net249
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[17\] VGND VGND VPWR VPWR net271
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[59\] VGND VGND VPWR VPWR net282
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold89 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[19\] VGND VGND VPWR VPWR net293
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2121__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2202__A myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_input49_X net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3612__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_69_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2951_ _0763_ _0767_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__nand2b_1
XANTENNA__2083__S net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3612__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1902_ net217 net61 net79 VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__mux2_1
X_2882_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[11\] _0717_ VGND VGND VPWR VPWR
+ _0718_ sky130_fd_sc_hd__nand2_1
X_1833_ myPWM.g_pwm_channel\[1\].CHANNEL.polarity _1521_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable
+ VGND VGND VPWR VPWR _1522_ sky130_fd_sc_hd__o21ai_1
XANTENNA__1926__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3503_ _1336_ _1337_ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3434_ _1135_ _1259_ VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__xnor2_1
XANTENNA__3208__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _1549_ _1199_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2316_ net125 _1727_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[7\] VGND VGND VPWR
+ VPWR _1732_ sky130_fd_sc_hd__a21oi_1
X_3296_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[57\]
+ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__nand2_2
X_2247_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[34\] VGND VGND VPWR VPWR
+ _1669_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_69_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2178_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[3\] VGND VGND VPWR VPWR
+ _1600_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_36_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1917__A1 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1845__B net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2590__B2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout96_A _1541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput68 net68 VGND VGND VPWR VPWR pwm_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_98_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1908__A1 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3150_ net108 _1639_ _0943_ _0954_ _0985_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__o2111a_1
XANTENNA__2078__S net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2101_ myPWM.g_pwm_channel\[0\].CHANNEL.alignment net56 _1545_ VGND VGND VPWR VPWR
+ _0243_ sky130_fd_sc_hd__mux2_1
X_3081_ _1626_ _0916_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__xnor2_1
X_2032_ _1547_ net336 net85 VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3983_ net178 VGND VGND VPWR VPWR rdata[6] sky130_fd_sc_hd__buf_2
XFILLER_0_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2934_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[32\] _0693_ _0692_ VGND
+ VGND VPWR VPWR _0770_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2865_ _0516_ _0518_ _0541_ _0510_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1816_ _1581_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[56\] net120 _1653_
+ VGND VGND VPWR VPWR _1505_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_0_CLK_X clknet_0_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2796_ _0628_ _0631_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3417_ _1243_ _1244_ _1247_ _1251_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__and4b_1
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3348_ _1078_ _1170_ _1087_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3279_ _1113_ VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3844__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout99_X net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2650_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[13\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[45\]
+ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2581_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[13\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[13\]
+ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_74_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3202_ _1035_ _1036_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3133_ _1603_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[36\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[35\]
+ _1601_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__o22a_1
X_3064_ _0495_ _0899_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2015_ net271 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[17\] net95 VGND
+ VGND VPWR VPWR _0161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3966_ clknet_leaf_26_CLK _0258_ net147 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_2917_ _0744_ _0750_ _0751_ _0752_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__and4_1
XFILLER_0_92_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3897_ clknet_leaf_24_CLK _0223_ net159 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[46\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2848_ net116 _0683_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2779_ _1625_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[58\] VGND VGND VPWR
+ VPWR _0615_ sky130_fd_sc_hd__nor2_1
XANTENNA__3664__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold131 myPWM.g_pwm_channel\[0\].CHANNEL.data_mod\[0\] VGND VGND VPWR VPWR net335
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout101_X net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold120 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[25\] VGND VGND VPWR VPWR net324
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2300__A net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3839__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_10_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3820_ clknet_leaf_23_CLK _0146_ net160 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_3751_ clknet_leaf_40_CLK _0111_ net130 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_mod\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2702_ _0537_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__inv_2
XANTENNA__2091__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3682_ clknet_leaf_42_CLK _0042_ net128 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_40_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2633_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\]
+ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2564_ net106 _0403_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\] VGND VGND VPWR
+ VPWR _0406_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3699__RESET_B net144 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2495_ net70 _0360_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3116_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[22\] _1637_ _1638_ net107 VGND VGND
+ VPWR VPWR _0952_ sky130_fd_sc_hd__o22a_1
X_3047_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[2\] _0878_ _0880_ _0882_ VGND VGND
+ VPWR VPWR _0883_ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2463__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3659__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout149_X net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3949_ clknet_leaf_39_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[26\]
+ net132 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[26\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_21_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2684__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_450 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout70 _0350_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_2
Xfanout81 _1534_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_4
XFILLER_0_36_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout92 _1544_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_4
XFILLER_0_101_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2280_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] _1563_ _1592_ net117
+ _1701_ VGND VGND VPWR VPWR _1702_ sky130_fd_sc_hd__o221a_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3485__A2 _1312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2086__S net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Left_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3803_ clknet_leaf_8_CLK _0129_ net157 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1995_ net279 net57 net73 VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__mux2_1
X_3734_ clknet_leaf_40_CLK _0094_ net139 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_41_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3665_ clknet_leaf_25_CLK _0025_ net147 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_2616_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] _0398_ _0447_ _0449_
+ _0452_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_42_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload40 clknet_leaf_22_CLK VGND VGND VPWR VPWR clkload40/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_93_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3596_ _1398_ _1402_ _1406_ _1430_ net124 VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__a32o_1
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2547_ net107 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[22\] _0390_ VGND VGND VPWR
+ VPWR _0395_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2478_ _0322_ _0323_ _0344_ _0346_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__or4_1
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2785__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_50_Left_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload1 clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout81_X net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2911__A1 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_input39_A wdata[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2103__B_N net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3984__179 VGND VGND VPWR VPWR _3984__179/HI net179 sky130_fd_sc_hd__conb_1
XFILLER_0_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3450_ _1059_ _1065_ _1284_ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__a21o_1
X_3381_ _1214_ _1215_ _1181_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__a21o_1
X_2401_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[0\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[0\]
+ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2332_ _1743_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[11\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_20_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2263_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[17\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\]
+ VGND VGND VPWR VPWR _1685_ sky130_fd_sc_hd__xor2_1
X_4002_ net197 VGND VGND VPWR VPWR rdata[25] sky130_fd_sc_hd__buf_2
X_2194_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[16\] VGND VGND VPWR VPWR _1616_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_46_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1978_ net252 net38 net76 VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__mux2_1
X_3717_ clknet_leaf_42_CLK _0077_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3648_ clknet_leaf_43_CLK _0008_ net133 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3579_ _1031_ _1296_ VGND VGND VPWR VPWR _1414_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold13 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[37\] VGND VGND VPWR VPWR net217
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[12\] VGND VGND VPWR VPWR net228
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[47\] VGND VGND VPWR VPWR net250
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[40\] VGND VGND VPWR VPWR net239
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[42\] VGND VGND VPWR VPWR net261
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[62\] VGND VGND VPWR VPWR net272
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[46\] VGND VGND VPWR VPWR net283
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3847__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_22_CLK_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_37_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1871__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2950_ _0763_ _0782_ _0784_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_57_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1901_ net212 net60 net79 VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__mux2_1
X_2881_ _0500_ _0716_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1832_ _1280_ _1456_ _1457_ _1520_ VGND VGND VPWR VPWR _1521_ sky130_fd_sc_hd__a31o_2
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3502_ _0995_ _0996_ _1326_ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_77_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3433_ _1122_ _1132_ VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[33\]
+ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3224__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2315_ net125 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[7\] _1727_ VGND VGND VPWR
+ VPWR _1731_ sky130_fd_sc_hd__and3_1
X_3295_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[57\]
+ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2246_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[35\] VGND VGND VPWR VPWR
+ _1668_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2177_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[2\] VGND VGND VPWR VPWR _1599_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_467 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1853__A1 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2100_ net339 net45 _1545_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__mux2_1
X_3080_ _0914_ _0915_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_6_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2031_ net12 net1 net23 _1542_ VGND VGND VPWR VPWR _1543_ sky130_fd_sc_hd__nor4b_2
XANTENNA__2094__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3982_ net177 VGND VGND VPWR VPWR rdata[5] sky130_fd_sc_hd__buf_2
XANTENNA__3597__A1 _1560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2933_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[32\] _0693_ VGND VGND VPWR
+ VPWR _0769_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2864_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\] _0686_ VGND VGND VPWR VPWR _0700_
+ sky130_fd_sc_hd__or2_1
X_1815_ _1591_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[61\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[59\]
+ _1587_ VGND VGND VPWR VPWR _1504_ sky130_fd_sc_hd__a2bb2o_1
X_2795_ _1631_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[63\] VGND VGND VPWR
+ VPWR _0631_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3219__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3416_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[16\] _1249_ _1250_ VGND VGND VPWR
+ VPWR _1251_ sky130_fd_sc_hd__o21ba_1
X_3347_ _1078_ _1170_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__xnor2_1
X_3278_ _1098_ _1110_ _1112_ _1107_ _1109_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2229_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[59\] VGND VGND VPWR VPWR
+ _1651_ sky130_fd_sc_hd__inv_2
XANTENNA__1901__S net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2260__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2260__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2012__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input21_A addr[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2251__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2003__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2580_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[12\]
+ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_74_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2089__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3201_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[33\]
+ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__nand2b_1
X_3132_ _1601_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[35\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[34\]
+ _1599_ _0967_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3063_ _0496_ _0852_ _0497_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__a21boi_1
X_2014_ net284 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] net94 VGND
+ VGND VPWR VPWR _0160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3965_ clknet_leaf_26_CLK _0257_ net148 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3896_ clknet_leaf_15_CLK _0222_ net166 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2916_ net106 _0749_ _0747_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2847_ _0516_ _0548_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2778_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] _1635_ _0613_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\]
+ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__a22o_1
Xhold110 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[55\] VGND VGND VPWR VPWR net314
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold121 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[27\] VGND VGND VPWR VPWR net325
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold132 myPWM.g_pwm_channel\[1\].CHANNEL.data_mod\[1\] VGND VGND VPWR VPWR net336
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3680__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3750_ clknet_leaf_41_CLK _0110_ net130 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2701_ _0535_ _0536_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_495 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3681_ clknet_leaf_43_CLK _0041_ net128 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2632_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\]
+ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2563_ net106 _0403_ _0405_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[27\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2494_ _0358_ _0359_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3115_ _1622_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[56\] _1636_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\]
+ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_65_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3046_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[0\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[1\]
+ _0769_ _0879_ _0881_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__o41a_1
XFILLER_0_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2463__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3948_ clknet_leaf_39_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[25\]
+ net131 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_21_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3675__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3879_ clknet_leaf_4_CLK _0205_ net150 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_2_1__f_CLK_X clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout71_A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout71 net72 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_2
Xfanout82 _1534_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_4
Xfanout93 _1544_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_2
XFILLER_0_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3317__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3802_ clknet_leaf_9_CLK _0128_ net157 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1994_ net323 net55 net73 VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__mux2_1
X_3733_ clknet_leaf_34_CLK _0093_ net139 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3664_ clknet_leaf_28_CLK _0024_ net147 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkload30 clknet_leaf_11_CLK VGND VGND VPWR VPWR clkload30/Y sky130_fd_sc_hd__inv_8
Xclkload41 clknet_leaf_23_CLK VGND VGND VPWR VPWR clkload41/X sky130_fd_sc_hd__clkbuf_8
X_2615_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] _0398_ _0451_ VGND
+ VGND VPWR VPWR _0452_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3595_ _1075_ _1429_ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2546_ net107 _0390_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[22\] VGND VGND VPWR
+ VPWR _0394_ sky130_fd_sc_hd__a21oi_1
X_2477_ _1604_ net116 _1612_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[13\] _0345_
+ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3029_ net115 _0864_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_54_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2306__A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload2 clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clkload2/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout74_X net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2675__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2427__B2 _1592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2400_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable _0270_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[0\]
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[0\] sky130_fd_sc_hd__mux2_1
X_3380_ net123 _1178_ _1184_ net124 VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2331_ net71 _1741_ _1742_ VGND VGND VPWR VPWR _1743_ sky130_fd_sc_hd__or3_1
XANTENNA__3942__RESET_B net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2262_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] net119 VGND VGND VPWR
+ VPWR _1684_ sky130_fd_sc_hd__or2_1
X_4001_ net196 VGND VGND VPWR VPWR rdata[24] sky130_fd_sc_hd__buf_2
XANTENNA__2097__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2193_ net111 VGND VGND VPWR VPWR _1615_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1977_ net228 net37 net76 VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3716_ clknet_leaf_42_CLK _0076_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_476 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3647_ clknet_leaf_43_CLK _0007_ net128 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3578_ _1196_ _1297_ VGND VGND VPWR VPWR _1413_ sky130_fd_sc_hd__xnor2_1
XANTENNA__3683__RESET_B net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2529_ net111 _0380_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[16\] VGND VGND VPWR
+ VPWR _0383_ sky130_fd_sc_hd__a21oi_1
XANTENNA__1904__S net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold14 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[11\] VGND VGND VPWR VPWR net218
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[5\] VGND VGND VPWR VPWR net240
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[17\] VGND VGND VPWR VPWR net251
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[16\] VGND VGND VPWR VPWR net229
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[23\] VGND VGND VPWR VPWR net262
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[7\] VGND VGND VPWR VPWR net273
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input51_A wdata[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1900_ net210 net59 net79 VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__mux2_1
X_2880_ _0504_ _0681_ _0560_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_72_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1831_ _1594_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[63\] _1671_ _1513_
+ _1519_ VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_37_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3773__Q myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_25_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3501_ _0996_ _1326_ _0995_ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_77_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3432_ _1585_ _1266_ VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[33\]
+ VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__and2_1
X_2314_ _1730_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[6\]
+ sky130_fd_sc_hd__inv_2
X_3294_ _1126_ _1127_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__nand2_1
X_2245_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[36\] VGND VGND VPWR VPWR
+ _1667_ sky130_fd_sc_hd__inv_2
XANTENNA__2639__B2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2639__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2176_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\] VGND VGND VPWR VPWR
+ _1598_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout169_A net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3948__Q myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_87_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout124_X net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3683__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input54_X net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2030_ net26 net27 net66 _1531_ VGND VGND VPWR VPWR _1542_ sky130_fd_sc_hd__and4b_1
XFILLER_0_69_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3981_ net176 VGND VGND VPWR VPWR rdata[4] sky130_fd_sc_hd__buf_2
X_2932_ _1602_ _1649_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2863_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\] _0686_ _0687_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[4\]
+ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__a22o_1
X_1814_ net118 _1651_ VGND VGND VPWR VPWR _1503_ sky130_fd_sc_hd__nor2_1
X_2794_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\] _0629_ VGND VGND VPWR VPWR
+ _0630_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3235__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3415_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] _1246_ _1249_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[16\]
+ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3346_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[12\] _1178_ _1180_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\]
+ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__a22o_1
X_3277_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] _1654_ _1111_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[17\]
+ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2228_ myPWM.g_pwm_channel\[0\].CHANNEL.polarity VGND VGND VPWR VPWR _1650_ sky130_fd_sc_hd__inv_2
X_2159_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[24\] VGND VGND VPWR VPWR _1581_
+ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_21_CLK_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3678__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[24\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2260__A2 _1560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_36_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input14_A addr[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3200_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[2\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[34\]
+ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__xnor2_2
X_3131_ _1599_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[34\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[33\]
+ _1597_ _0966_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__o221a_1
X_3062_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[14\] _0853_ _0858_ _0897_ VGND VGND
+ VPWR VPWR _0898_ sky130_fd_sc_hd__a2bb2o_1
X_2013_ net332 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\] net96 VGND
+ VGND VPWR VPWR _0159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3964_ clknet_leaf_27_CLK _0256_ net148 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_3895_ clknet_leaf_16_CLK _0221_ net166 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[44\]
+ sky130_fd_sc_hd__dfrtp_2
X_2915_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[24\] _0746_ _0745_ VGND VGND VPWR
+ VPWR _0751_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_45_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2846_ _0504_ _0681_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2777_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[59\] _0597_ VGND VGND VPWR
+ VPWR _0613_ sky130_fd_sc_hd__nor2_1
Xhold100 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[58\] VGND VGND VPWR VPWR net304
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold111 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[56\] VGND VGND VPWR VPWR net315
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[10\] VGND VGND VPWR VPWR net326
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 myPWM.g_pwm_channel\[1\].CHANNEL.data_mod\[0\] VGND VGND VPWR VPWR net337
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2140__Y _1562_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input6_A addr[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3329_ _0998_ _1139_ _1143_ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__and3_1
XANTENNA__1912__S net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3258__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2309__A net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1992__A1 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2700_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[37\]
+ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__and2_1
XANTENNA__1983__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3680_ clknet_leaf_43_CLK _0040_ net133 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2631_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] _1636_ VGND VGND VPWR
+ VPWR _0467_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2562_ net106 _0403_ net69 VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2493_ _1603_ _0356_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3114_ net108 _1639_ _0948_ _0949_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__a211o_1
X_3045_ _0528_ _0770_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_419 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout151_A net154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3947_ clknet_leaf_39_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[24\]
+ net131 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[24\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1974__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3878_ clknet_leaf_4_CLK _0204_ net152 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_21_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2829_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] _0660_ _0664_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[16\]
+ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__a22oi_1
XANTENNA__1907__S net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_3__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_2_3__leaf_CLK sky130_fd_sc_hd__clkbuf_16
Xfanout72 _1712_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout83 _1534_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_4
XFILLER_0_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout94 _1541_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_4
XANTENNA__1965__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3801_ clknet_leaf_12_CLK _0127_ net159 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1993_ net311 net54 net73 VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3732_ clknet_leaf_24_CLK _0092_ net145 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[45\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload20 clknet_leaf_34_CLK VGND VGND VPWR VPWR clkload20/Y sky130_fd_sc_hd__clkinv_2
X_3663_ clknet_leaf_26_CLK _0023_ net147 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload31 clknet_leaf_12_CLK VGND VGND VPWR VPWR clkload31/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2614_ _1618_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[19\] _0393_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\]
+ _0450_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__o221a_1
Xclkload42 clknet_leaf_24_CLK VGND VGND VPWR VPWR clkload42/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__3227__B myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[46\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3594_ _1078_ _1399_ _1076_ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2545_ _0393_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[21\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_76_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2476_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] _1611_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\]
+ _1599_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_76_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3028_ _0555_ _0782_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_54_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout154_X net154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload3 clknet_leaf_0_CLK VGND VGND VPWR VPWR clkload3/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2124__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3328__A net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2330_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[9\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[10\]
+ net124 _1734_ VGND VGND VPWR VPWR _1742_ sky130_fd_sc_hd__and4_1
X_2261_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] net119 VGND VGND VPWR
+ VPWR _1683_ sky130_fd_sc_hd__nand2_1
X_4000_ net195 VGND VGND VPWR VPWR rdata[23] sky130_fd_sc_hd__buf_2
XANTENNA__2115__A1 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2192_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[15\] VGND VGND VPWR VPWR
+ _1614_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1976_ net215 net36 net76 VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3715_ clknet_leaf_42_CLK _0075_ net128 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3238__A _1562_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3646_ clknet_leaf_44_CLK _0006_ net133 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3577_ _1046_ _1299_ VGND VGND VPWR VPWR _1412_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2528_ net111 _0380_ _0382_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[15\]
+ sky130_fd_sc_hd__a21oi_1
Xhold37 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[31\] VGND VGND VPWR VPWR net241
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[63\] VGND VGND VPWR VPWR net230
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] _1627_ _1628_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\]
+ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__o22a_1
Xhold15 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[43\] VGND VGND VPWR VPWR net219
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2106__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold48 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[13\] VGND VGND VPWR VPWR net252
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[44\] VGND VGND VPWR VPWR net263
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3652__RESET_B net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1920__S net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2317__A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2593__B2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input44_A wdata[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3990__185 VGND VGND VPWR VPWR _3990__185/HI net185 sky130_fd_sc_hd__conb_1
XFILLER_0_57_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1830_ _1510_ _1514_ _1517_ _1518_ _1502_ VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__a41o_1
XFILLER_0_44_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3500_ _1326_ _1334_ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3431_ _1260_ _1265_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_90_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ _1040_ _1196_ VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2313_ net125 _1727_ _1729_ VGND VGND VPWR VPWR _1730_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_29_Left_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3293_ _1126_ _1127_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__and2_1
X_2244_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[37\] VGND VGND VPWR VPWR
+ _1666_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2175_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[1\] VGND VGND VPWR VPWR _1597_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_38_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1959_ net295 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[61\] net98 VGND
+ VGND VPWR VPWR _0108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout117_X net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3629_ _1459_ _1462_ _1463_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1915__S net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_40_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_40_CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA_input47_X net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3980_ net175 VGND VGND VPWR VPWR rdata[3] sky130_fd_sc_hd__buf_2
XANTENNA__2254__B1 _1592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2931_ _0500_ _0502_ _0766_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[44\]
+ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] VGND VGND VPWR VPWR _0767_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_57_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2862_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[4\] _0687_ _0689_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[3\]
+ _0697_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__o221a_1
X_1813_ _1594_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[63\] VGND VGND VPWR
+ VPWR _1502_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_13_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2793_ _0462_ _0627_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__xnor2_1
XANTENNA__2557__A1 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_25_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3414_ _1238_ _1248_ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3506__B1 _1671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_31_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_31_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3345_ _1065_ _1179_ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3276_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[49\] _1105_ VGND VGND VPWR
+ VPWR _1111_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2227_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[36\] VGND VGND VPWR VPWR
+ _1649_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2138__Y _1560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2158_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] VGND VGND VPWR VPWR
+ _1580_ sky130_fd_sc_hd__inv_2
X_2089_ net266 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[55\] net90 VGND
+ VGND VPWR VPWR _0232_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout94_A _1541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_CLK clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_22_CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__3161__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_CLK clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_13_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_74_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3130_ _1597_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[33\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[32\]
+ _1595_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3996__191 VGND VGND VPWR VPWR _3996__191/HI net191 sky130_fd_sc_hd__conb_1
X_3061_ _0890_ _0894_ _0896_ _0857_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2012_ net316 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] net96 VGND
+ VGND VPWR VPWR _0158_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2778__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3963_ clknet_leaf_26_CLK _0255_ net148 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3894_ clknet_leaf_17_CLK _0220_ net168 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[43\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_70_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2778__B2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2914_ net106 _0749_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__or2_1
X_2845_ _0507_ _0556_ _0558_ _0508_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__a31o_1
Xhold101 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[53\] VGND VGND VPWR VPWR net305
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2776_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[59\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\]
+ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__and2b_1
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3246__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold134 myPWM.g_pwm_channel\[0\].CHANNEL.data_mod\[1\] VGND VGND VPWR VPWR net338
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[21\] VGND VGND VPWR VPWR net327
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[14\] VGND VGND VPWR VPWR net316
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2150__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3328_ net117 _1161_ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3259_ _1058_ _1084_ _1093_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_68_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout97_X net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2457__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_2_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_2_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2630_ _0465_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2561_ _0403_ _0404_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[26\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_20_CLK_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2492_ _1603_ _0356_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_35_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3113_ net107 _1638_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__and2_1
X_3044_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[0\] _0769_ _0879_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[1\]
+ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__o31a_1
XFILLER_0_77_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3946_ clknet_leaf_39_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[23\]
+ net131 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout144_A net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3877_ clknet_leaf_5_CLK _0203_ net152 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_21_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2828_ _0570_ _0577_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__xor2_1
XFILLER_0_14_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2759_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[60\]
+ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__or2_1
XANTENNA__1923__S net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout73 _1540_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_4
Xfanout95 _1541_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_2
XFILLER_0_36_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout84 _1534_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_2
XFILLER_0_101_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3800_ clknet_leaf_12_CLK _0126_ net159 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3770__RESET_B net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1992_ net325 net53 net73 VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__mux2_1
X_3731_ clknet_leaf_25_CLK _0091_ net145 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[44\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_70_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_306 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload10 clknet_leaf_41_CLK VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__inv_8
X_3662_ clknet_leaf_27_CLK _0022_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_3593_ _1560_ _1400_ VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__nor2_1
Xclkload32 clknet_leaf_13_CLK VGND VGND VPWR VPWR clkload32/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2613_ _1614_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[15\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[17\]
+ _1617_ _0418_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__a221oi_1
Xclkload21 clknet_leaf_35_CLK VGND VGND VPWR VPWR clkload21/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_11_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2544_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[21\] _0390_ _0392_ VGND VGND VPWR
+ VPWR _0393_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_93_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2475_ _1617_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] _1631_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[31\]
+ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_76_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3027_ _0860_ _0861_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[9\] VGND VGND VPWR
+ VPWR _0863_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_54_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3858__RESET_B net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3929_ clknet_leaf_35_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[6\] net141
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[6\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__1918__S net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload4 clknet_leaf_1_CLK VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_61_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3321__A1 _1592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1883__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1895__Y _1537_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2060__A1 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2260_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] _1560_ _1574_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\]
+ _1681_ VGND VGND VPWR VPWR _1682_ sky130_fd_sc_hd__a221o_1
XANTENNA__3201__A_N myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2191_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[14\] VGND VGND VPWR VPWR _1613_
+ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_2_2__f_CLK_A clknet_0_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1975_ net253 net35 net75 VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2051__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2423__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3714_ clknet_leaf_43_CLK _0074_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3645_ clknet_leaf_44_CLK _0005_ net133 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3576_ _1025_ _1410_ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2527_ net111 _0380_ net69 VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__o21ai_1
XANTENNA__3254__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2458_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] _1610_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\]
+ _1613_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__o22a_1
XFILLER_0_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold16 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[4\] VGND VGND VPWR VPWR net220
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[38\] VGND VGND VPWR VPWR net242
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[32\] VGND VGND VPWR VPWR net231
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[10\] VGND VGND VPWR VPWR net253
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2389_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[28\] VGND VGND VPWR VPWR
+ _1783_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2042__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input37_A wdata[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1856__A1 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2281__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2033__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3430_ _1128_ _1141_ _1258_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3361_ _1027_ _1028_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__nand2_2
XFILLER_0_0_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2312_ net125 _1727_ _1713_ VGND VGND VPWR VPWR _1729_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3292_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[59\]
+ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2243_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[38\] VGND VGND VPWR VPWR
+ _1665_ sky130_fd_sc_hd__inv_2
X_2174_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\] VGND VGND VPWR VPWR
+ _1596_ sky130_fd_sc_hd__inv_2
XANTENNA__1847__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2153__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__2024__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1958_ net313 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[60\] net98 VGND
+ VGND VPWR VPWR _0107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1889_ net308 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] net102 VGND
+ VGND VPWR VPWR _0041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3628_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[14\] _1658_ VGND VGND VPWR VPWR
+ _1463_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3559_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[12\] _1391_ _1393_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\]
+ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__a22oi_1
XANTENNA__1931__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2002__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkload2_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2254__B2 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2254__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2930_ _0765_ _0503_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_84_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2006__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2861_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[3\] _0689_ _0691_ _0696_ VGND VGND
+ VPWR VPWR _0697_ sky130_fd_sc_hd__a22o_1
X_1812_ _1490_ _1491_ _1492_ _1498_ _1500_ VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_13_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2792_ _1630_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[62\] _0624_ _0626_
+ _0462_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__a221oi_2
XTAP_TAPCELL_ROW_41_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_584 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3413_ _1094_ _1101_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__and2_1
XANTENNA__3506__A1 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3344_ _1089_ _1172_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__nor2_1
X_3275_ _1570_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[51\] VGND VGND VPWR
+ VPWR _1110_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2226_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[40\] VGND VGND VPWR VPWR
+ _1648_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2157_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\] VGND VGND VPWR VPWR _1579_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2088_ net321 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[54\] net90 VGND
+ VGND VPWR VPWR _0231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1926__S net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout87_A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3060_ net112 _0855_ _0892_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[11\] _0895_
+ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__o221ai_1
X_2011_ net252 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] net97 VGND
+ VGND VPWR VPWR _0157_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_66_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3962_ clknet_leaf_29_CLK _0254_ net149 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_3893_ clknet_leaf_17_CLK _0219_ net168 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[42\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_73_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2913_ _0597_ _0748_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2844_ net113 _0678_ _0679_ net112 VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_9_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2431__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2775_ _0478_ _0586_ _0592_ _0610_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_96_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold124 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[51\] VGND VGND VPWR VPWR net328
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 myPWM.g_pwm_channel\[1\].CHANNEL.polarity VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 myPWM.g_pwm_channel\[0\].CHANNEL.polarity VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[60\] VGND VGND VPWR VPWR net306
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_84_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3327_ _1594_ _1157_ _1158_ VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__and3_1
XANTENNA__3262__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3258_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] _1656_ _1071_ _1088_
+ _1092_ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__a221o_1
X_3189_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[38\]
+ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__nor2_1
X_2209_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\] VGND VGND VPWR VPWR
+ _1631_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2606__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_93_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2393__B1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2560_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[26\] _0401_ net69 VGND VGND VPWR
+ VPWR _0404_ sky130_fd_sc_hd__o21ai_1
X_2491_ net70 _0356_ _0357_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[3\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_50_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3112_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[20\] _1639_ _0946_ _0947_ VGND VGND
+ VPWR VPWR _0948_ sky130_fd_sc_hd__o22a_1
X_3043_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[32\] _0693_ VGND VGND VPWR
+ VPWR _0879_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3945_ clknet_leaf_39_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[22\]
+ net131 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[22\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_85_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2620__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3876_ clknet_leaf_4_CLK _0202_ net150 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2827_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] _0660_ _0662_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\]
+ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__o22a_1
X_2758_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[60\]
+ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2689_ _0522_ _0523_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__or2_1
XANTENNA__2100__S _1545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout74 _1540_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout96 _1541_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_4
Xfanout85 net89 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_4
XANTENNA__3167__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2010__S net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1991_ net280 net52 net73 VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3730_ clknet_leaf_25_CLK _0090_ net147 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[43\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_51_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_446 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3661_ clknet_leaf_26_CLK _0021_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkload33 clknet_leaf_14_CLK VGND VGND VPWR VPWR clkload33/Y sky130_fd_sc_hd__clkinv_8
X_3592_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[8\] _1403_ VGND VGND VPWR VPWR _1427_
+ sky130_fd_sc_hd__or2_1
Xclkload11 clknet_leaf_42_CLK VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__inv_4
X_2612_ _1618_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[19\] _0393_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\]
+ _0448_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__a221o_1
Xclkload22 clknet_leaf_2_CLK VGND VGND VPWR VPWR clkload22/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2543_ net107 _0390_ net70 VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2474_ _0308_ _0318_ _0329_ _0342_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__or4_1
XFILLER_0_76_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3026_ _0860_ _0861_ net114 VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_54_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3928_ clknet_leaf_34_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[5\] net141
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\] sky130_fd_sc_hd__dfrtp_4
Xclkload5 clknet_leaf_36_CLK VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_34_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3827__RESET_B net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3859_ clknet_leaf_20_CLK _0185_ net164 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1934__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_34_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2005__S net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2348__B1 _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2190_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[13\] VGND VGND VPWR VPWR
+ _1612_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1974_ net260 net65 net76 VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3713_ clknet_leaf_43_CLK _0073_ net133 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3644_ clknet_leaf_0_CLK _0004_ net134 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3575_ _1046_ _1299_ _1043_ VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__a21oi_1
X_2526_ _0380_ _0381_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[14\]
+ sky130_fd_sc_hd__nor2_1
X_2457_ _1602_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[4\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[25\]
+ _1624_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__o22a_1
Xhold28 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[2\] VGND VGND VPWR VPWR net232
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold17 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[6\] VGND VGND VPWR VPWR net221
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[41\] VGND VGND VPWR VPWR net243
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2388_ _1781_ _1782_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[28\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__2511__B1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3270__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3009_ _0577_ _0792_ _0576_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout72_X net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2502__B1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3749__RESET_B net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2693__A_N myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3360_ _1042_ _1046_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__xnor2_1
X_2311_ _1728_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[5\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3291_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[59\]
+ VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2242_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[39\] VGND VGND VPWR VPWR
+ _1664_ sky130_fd_sc_hd__inv_2
X_2173_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[0\] VGND VGND VPWR VPWR _1595_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1957_ net299 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[59\] net98 VGND
+ VGND VPWR VPWR _0106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1888_ net234 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] net103 VGND
+ VGND VPWR VPWR _0040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3627_ _1460_ _1461_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3558_ _1065_ _1392_ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_8_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2509_ _0351_ _0369_ _0370_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__or3_1
X_3489_ _1124_ _1126_ _1123_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_11_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3451__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2860_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[2\] _0690_ _0694_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[1\]
+ _0695_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1811_ _1484_ _1485_ _1487_ _1488_ _1499_ VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__o221a_1
XFILLER_0_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2791_ _1630_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[62\] _0624_ _0626_
+ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3412_ net121 _1242_ _1246_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] VGND VGND
+ VPWR VPWR _1247_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3343_ _1172_ _1177_ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3274_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\]
+ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__and2b_1
XFILLER_0_84_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2225_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[42\] VGND VGND VPWR VPWR
+ _1647_ sky130_fd_sc_hd__inv_2
X_2156_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] VGND VGND VPWR VPWR
+ _1578_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2087_ net305 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[53\] net91 VGND
+ VGND VPWR VPWR _0230_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout167_A net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2164__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2989_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\] _0819_ VGND VGND VPWR VPWR
+ _0825_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2170__Y _1592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2330__C net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3980__175 VGND VGND VPWR VPWR _3980__175/HI net175 sky130_fd_sc_hd__conb_1
XANTENNA__1942__S net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1995__A1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2013__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input52_X net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1852__S net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2010_ net228 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\] net97 VGND
+ VGND VPWR VPWR _0156_ sky130_fd_sc_hd__mux2_1
XANTENNA__3764__RESET_B net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3424__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3961_ clknet_leaf_26_CLK _0253_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2912_ _0601_ _0739_ _0612_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__a21oi_1
XANTENNA__1986__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3892_ clknet_leaf_19_CLK _0218_ net167 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[41\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2843_ _0491_ _0671_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2774_ _0602_ _0605_ _0609_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__nand3_1
XFILLER_0_53_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold114 myPWM.g_pwm_channel\[1\].CHANNEL.pwm_next VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[1\] VGND VGND VPWR VPWR net307
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold125 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[22\] VGND VGND VPWR VPWR net329
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 myPWM.g_pwm_channel\[1\].CHANNEL.alignment VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__dlygate4sd3_1
X_3326_ _1153_ _1156_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__xnor2_1
XANTENNA__1910__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3257_ _1090_ _1091_ _1070_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__o21a_1
X_3188_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[38\]
+ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__and2_1
X_2208_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] VGND VGND VPWR VPWR
+ _1630_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2139_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[11\] VGND VGND VPWR VPWR
+ _1561_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1977__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1937__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1901__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input12_A addr[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2008__S net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1968__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1847__S net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2490_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[3\] _0354_ VGND VGND VPWR VPWR _0357_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_49_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3363__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3111_ net109 _1640_ _0940_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__o21a_1
X_3042_ _0524_ _0771_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3944_ clknet_leaf_39_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[21\]
+ net131 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3875_ clknet_leaf_5_CLK _0201_ net152 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_2826_ _0484_ _0661_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2757_ _0586_ _0591_ _0478_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2688_ _0522_ _0523_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input4_A addr[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3309_ _1139_ _1143_ _0998_ VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout86 net89 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_4
Xfanout97 _1541_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_2
XFILLER_0_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout75 _1540_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_4
XANTENNA__1894__C net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3986__181 VGND VGND VPWR VPWR _3986__181/HI net181 sky130_fd_sc_hd__conb_1
XFILLER_0_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3324__B1 _1594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_8_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1990_ net324 net51 net73 VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2262__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3660_ clknet_leaf_29_CLK _0020_ net143 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkload34 clknet_leaf_15_CLK VGND VGND VPWR VPWR clkload34/Y sky130_fd_sc_hd__clkinv_4
X_3591_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[7\] _1409_ _1423_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[6\]
+ VGND VGND VPWR VPWR _1426_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2611_ _1614_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[15\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[17\]
+ _1617_ _0419_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_35_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload12 clknet_leaf_44_CLK VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload23 clknet_leaf_3_CLK VGND VGND VPWR VPWR clkload23/Y sky130_fd_sc_hd__inv_6
XFILLER_0_23_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2542_ _0390_ _0391_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[20\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_93_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2473_ _1598_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[2\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\]
+ _1627_ _0310_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__a221o_1
XANTENNA__2118__A1 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3025_ _0555_ _0782_ _0509_ _0554_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_92_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2437__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3927_ clknet_leaf_34_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[4\] net141
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[4\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_34_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3858_ clknet_leaf_20_CLK _0184_ net168 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[39\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload6 clknet_leaf_37_CLK VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__clkinv_8
X_2809_ _0630_ _0633_ _0644_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__and3_1
X_3789_ clknet_leaf_22_CLK _0115_ net162 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2109__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2111__S net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1950__S net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3178__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2021__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1860__S net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1973_ net301 net64 net75 VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__mux2_1
XANTENNA__2704__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3712_ clknet_leaf_43_CLK _0072_ net128 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3643_ clknet_leaf_0_CLK _0003_ net134 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_3574_ _1054_ _1408_ VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__xnor2_1
XANTENNA__3960__RESET_B net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2525_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[14\] _0379_ _0350_ VGND VGND VPWR
+ VPWR _0381_ sky130_fd_sc_hd__o21ai_1
X_2456_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\]
+ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__xor2_1
Xhold18 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[56\] VGND VGND VPWR VPWR net222
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[12\] VGND VGND VPWR VPWR net233
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2387_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[28\] _1779_ _1713_ VGND VGND VPWR
+ VPWR _1782_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2275__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3008_ _0484_ _0841_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1945__S net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2508__C net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2016__S net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1855__S net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_43_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_43_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2310_ net71 _1726_ _1727_ VGND VGND VPWR VPWR _1728_ sky130_fd_sc_hd__or3_1
X_3290_ _1123_ _1124_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__nor2_2
XFILLER_0_20_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2241_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[41\] VGND VGND VPWR VPWR
+ _1663_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2172_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] VGND VGND VPWR VPWR _1594_
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1956_ net304 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[58\] net99 VGND
+ VGND VPWR VPWR _0105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1887_ net257 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[25\] net102 VGND
+ VGND VPWR VPWR _0039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3626_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\] _1659_ _1660_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[12\]
+ VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_34_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_34_CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__2450__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3557_ _1061_ _1309_ _1059_ VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_8_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2508_ net116 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\] net115 _0362_ VGND VGND
+ VPWR VPWR _0370_ sky130_fd_sc_hd__and4_1
X_3488_ _1282_ _1321_ _1322_ _1135_ _1132_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__a2111oi_2
XANTENNA__3281__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2439_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\]
+ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_33_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_25_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_25_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_76_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input42_A wdata[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3191__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2487__B1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1810_ _1494_ _1495_ _1496_ VGND VGND VPWR VPWR _1499_ sky130_fd_sc_hd__or3b_1
XFILLER_0_38_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2790_ _1630_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[62\] _0625_ VGND
+ VGND VPWR VPWR _0626_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_16_CLK clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_16_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3411_ _1105_ _1245_ VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__xnor2_1
X_3342_ _1171_ _1088_ _1061_ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3273_ _1101_ _1105_ _1107_ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__or3b_1
X_2224_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[43\] VGND VGND VPWR VPWR
+ _1646_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2155_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[22\] VGND VGND VPWR VPWR _1577_
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2086_ net276 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\] net91 VGND
+ VGND VPWR VPWR _0229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_444 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2988_ _0812_ _0822_ _0823_ myPWM.g_pwm_channel\[0\].CHANNEL.alignment VGND VGND
+ VPWR VPWR _0824_ sky130_fd_sc_hd__and4b_1
XFILLER_0_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1939_ net216 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[41\] net101 VGND
+ VGND VPWR VPWR _0088_ sky130_fd_sc_hd__mux2_1
XANTENNA__2180__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout115_X net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2953__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3609_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[16\] _1382_ _1442_ net122 VGND VGND
+ VPWR VPWR _1444_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2683__A_N myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3186__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input45_X net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_5_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_5_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_18_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3960_ clknet_leaf_29_CLK _0252_ net149 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2911_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] _0742_ _0746_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[24\]
+ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__a22o_1
X_3891_ clknet_leaf_20_CLK _0217_ net164 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[40\]
+ sky130_fd_sc_hd__dfrtp_4
X_2842_ _0488_ _0670_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2773_ _0607_ _0608_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__nand2_2
XFILLER_0_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2396__C1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold115 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[29\] VGND VGND VPWR VPWR net319
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[27\] VGND VGND VPWR VPWR net308
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[48\] VGND VGND VPWR VPWR net330
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3325_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] _1149_ _1150_ _1159_ VGND VGND
+ VPWR VPWR _1160_ sky130_fd_sc_hd__o31a_1
X_3256_ _1063_ _1089_ _1069_ _1062_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__o211a_1
X_2207_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\] VGND VGND VPWR VPWR _1629_
+ sky130_fd_sc_hd__inv_2
X_3187_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] _1665_ VGND VGND VPWR
+ VPWR _1022_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2138_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[10\] VGND VGND VPWR VPWR _1560_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2069_ net258 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[35\] net92 VGND
+ VGND VPWR VPWR _0212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2114__S net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1953__S net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout92_A _1544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3351__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2024__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1863__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3110_ _0943_ _0945_ _0942_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3041_ _0688_ _0772_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__xnor2_1
X_3943_ clknet_leaf_38_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[20\]
+ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3874_ clknet_leaf_6_CLK _0200_ net155 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2825_ _0571_ _0574_ _0577_ _0582_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2756_ _0478_ _0591_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__and2_1
X_2687_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[3\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[35\]
+ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3308_ _1120_ _1121_ _1137_ _1142_ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__o31a_1
X_3239_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\] _1660_ VGND VGND VPWR
+ VPWR _1074_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_57_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2109__S net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1948__S net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2633__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout76 _1540_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_2
Xfanout98 _1538_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_4
XFILLER_0_24_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout87 net89 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_20_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3227__A_N myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout95_X net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1886__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[24\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2019__S net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1858__S net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2063__A1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload35 clknet_leaf_16_CLK VGND VGND VPWR VPWR clkload35/Y sky130_fd_sc_hd__inv_8
Xclkload24 clknet_leaf_5_CLK VGND VGND VPWR VPWR clkload24/Y sky130_fd_sc_hd__inv_6
X_3590_ _1421_ _1422_ _1424_ VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__o21a_1
X_2610_ _1621_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[24\] VGND VGND VPWR
+ VPWR _0447_ sky130_fd_sc_hd__xnor2_1
Xclkload13 clknet_leaf_25_CLK VGND VGND VPWR VPWR clkload13/X sky130_fd_sc_hd__clkbuf_8
X_2541_ net108 _0389_ net70 VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2472_ _1620_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[21\] _0312_ _0331_ _0340_
+ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__a2111o_1
XANTENNA__2718__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3024_ _0782_ _0783_ _0764_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2054__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3926_ clknet_leaf_34_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[3\] net139
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[3\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_34_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3857_ clknet_leaf_21_CLK _0183_ net163 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload7 clknet_leaf_38_CLK VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_41_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2808_ _0641_ _0642_ _0643_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__and3b_1
X_3788_ clknet_leaf_23_CLK _0114_ net160 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3554__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_2739_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[17\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[49\]
+ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2628__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[24\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2045__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2363__A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3194__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1859__A1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2284__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2036__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1972_ net275 net63 net75 VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3711_ clknet_leaf_43_CLK _0071_ net133 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3642_ clknet_leaf_0_CLK _0002_ net134 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_3573_ _1019_ _1407_ _1020_ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2524_ net113 net112 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[14\] _0375_ VGND VGND
+ VPWR VPWR _0380_ sky130_fd_sc_hd__and4_1
X_2455_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[16\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[16\]
+ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__xor2_1
X_2386_ net118 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[28\] _1776_ VGND VGND VPWR
+ VPWR _1781_ sky130_fd_sc_hd__and3_1
Xhold19 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[38\] VGND VGND VPWR VPWR net223
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3007_ _0481_ _0842_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2027__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3909_ clknet_leaf_5_CLK _0235_ net154 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[58\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_7_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2122__S net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1961__S net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3670__RESET_B net144 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2358__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2266__B2 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3189__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2018__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1871__S net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2240_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[42\] VGND VGND VPWR VPWR
+ _1662_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2171_ net117 VGND VGND VPWR VPWR _1593_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2257__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_73_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1955_ net310 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[57\] net98 VGND
+ VGND VPWR VPWR _0104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3509__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_1886_ net207 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[24\] net102 VGND
+ VGND VPWR VPWR _0038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3625_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[14\] _1658_ _1659_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\]
+ _1459_ VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__o221a_1
XFILLER_0_31_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3556_ _1061_ _1309_ VGND VGND VPWR VPWR _1391_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_8_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout105_A _1535_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2507_ net115 _0367_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__nor2_1
X_3487_ _1125_ _1128_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__nand2_1
X_2438_ _0297_ _0306_ _0307_ _0268_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.rollover_flag_c
+ sky130_fd_sc_hd__and4b_1
X_2369_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\] _1767_ VGND VGND VPWR VPWR
+ _1769_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2117__S net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1956__S net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input35_A wdata[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2027__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1866__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2411__B2 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3939__RESET_B net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3410_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[17\] _1655_ _1238_ VGND
+ VGND VPWR VPWR _1245_ sky130_fd_sc_hd__a21oi_1
X_3341_ _1069_ _1173_ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3272_ _1098_ _1104_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__and2_1
X_2223_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[44\] VGND VGND VPWR VPWR
+ _1645_ sky130_fd_sc_hd__inv_2
X_2154_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND VPWR VPWR
+ _1576_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2085_ net328 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[51\] net91 VGND
+ VGND VPWR VPWR _0228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2987_ _0813_ _0814_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\] VGND VGND VPWR
+ VPWR _0823_ sky130_fd_sc_hd__or3b_1
XFILLER_0_8_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2461__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_1938_ net239 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[40\] net100 VGND
+ VGND VPWR VPWR _0087_ sky130_fd_sc_hd__mux2_1
X_1869_ net273 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] net104 VGND
+ VGND VPWR VPWR _0021_ sky130_fd_sc_hd__mux2_1
XANTENNA__2953__A2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3608_ net122 _1442_ _1438_ _1564_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3539_ _1118_ _1319_ _1320_ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__nand3_1
XANTENNA__3292__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2636__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_17_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input38_X net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload0_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2910_ _0593_ _0605_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__xnor2_1
X_3890_ clknet_leaf_18_CLK _0216_ net168 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[39\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_85_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2841_ _0673_ _0676_ _1613_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__a21oi_1
XANTENNA__3773__RESET_B net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2772_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[58\]
+ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_44_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold116 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[18\] VGND VGND VPWR VPWR net320
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold105 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[31\] VGND VGND VPWR VPWR net309
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold127 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[61\] VGND VGND VPWR VPWR net331
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3324_ _1157_ _1158_ _1594_ VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__a21o_1
X_3255_ _1565_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[47\] VGND VGND VPWR
+ VPWR _1090_ sky130_fd_sc_hd__nor2_1
X_2206_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] VGND VGND VPWR VPWR
+ _1628_ sky130_fd_sc_hd__inv_2
X_3186_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[39\]
+ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__xor2_2
X_2137_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[9\] VGND VGND VPWR VPWR _1559_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2456__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Left_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2068_ net255 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[34\] net92 VGND
+ VGND VPWR VPWR _0211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2387__B1 _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_62_Left_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout85_A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2366__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2614__B2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_80_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2532__C myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_49_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2040__S net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2550__B1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3040_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[4\] _0875_ VGND VGND VPWR VPWR _0876_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_81_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3942_ clknet_leaf_38_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[19\]
+ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[19\] sky130_fd_sc_hd__dfrtp_1
X_3873_ clknet_leaf_6_CLK _0199_ net155 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2824_ _0574_ _0659_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2755_ _0473_ _0476_ _0589_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__or3_1
X_2686_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[3\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[35\]
+ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3307_ _1125_ _1128_ _1141_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__or3_1
XANTENNA__2541__B1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3238_ _1562_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[44\] VGND VGND VPWR
+ VPWR _1073_ sky130_fd_sc_hd__nor2_1
X_3169_ _1000_ _1002_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__nand2_1
XANTENNA__2186__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout88 _1543_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_2
XFILLER_0_9_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout77 _1537_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_4
Xfanout99 _1538_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_20_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout88_X net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2035__S net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload25 clknet_leaf_6_CLK VGND VGND VPWR VPWR clkload25/Y sky130_fd_sc_hd__clkinv_2
Xclkload14 clknet_leaf_26_CLK VGND VGND VPWR VPWR clkload14/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__1874__S net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload36 clknet_leaf_17_CLK VGND VGND VPWR VPWR clkload36/Y sky130_fd_sc_hd__inv_8
XFILLER_0_11_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2540_ net110 net109 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[20\] _0385_ VGND VGND
+ VPWR VPWR _0390_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_93_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2471_ _0311_ _0337_ _0338_ _0339_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__or4_1
XFILLER_0_50_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3023_ _0513_ _0781_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_54_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3251__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3925_ clknet_leaf_33_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[2\] net139
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[2\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_62_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload8 clknet_leaf_39_CLK VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_33_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3856_ clknet_leaf_21_CLK _0182_ net163 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3787_ clknet_leaf_20_CLK _0113_ net167 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2807_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\] _0634_ VGND VGND VPWR VPWR
+ _0643_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2738_ _0572_ _0573_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__nand2_2
XFILLER_0_41_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2669_ _0500_ _0504_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1813__A _1594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2293__A2 myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1959__S net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2475__A2_N myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input65_A wdata[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1869__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3710_ clknet_leaf_0_CLK _0070_ net136 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[55\]
+ sky130_fd_sc_hd__dfrtp_1
X_1971_ net221 net62 net75 VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3641_ clknet_leaf_1_CLK _0001_ net134 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_3572_ _1299_ _1300_ _1302_ _1023_ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2523_ _0351_ _0378_ _0379_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[13\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_11_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2454_ _1595_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[0\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[3\]
+ _1601_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__a22o_1
X_2385_ _1780_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[27\]
+ sky130_fd_sc_hd__inv_2
Xinput1 addr[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_67_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2275__A2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_3006_ _0484_ _0841_ _0483_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3908_ clknet_leaf_3_CLK _0234_ net151 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[57\]
+ sky130_fd_sc_hd__dfrtp_2
X_3839_ clknet_leaf_6_CLK _0165_ net155 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3295__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3463__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2374__A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3798__RESET_B net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2170_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\] VGND VGND VPWR VPWR
+ _1592_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2257__A2 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1954_ net315 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[56\] net98 VGND
+ VGND VPWR VPWR _0103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2731__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3624_ net122 _1657_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__nand2_1
X_1885_ net312 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] net102 VGND
+ VGND VPWR VPWR _0037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3555_ _1387_ _1388_ _1389_ VGND VGND VPWR VPWR _1390_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_8_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3486_ _1319_ _1320_ _1283_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_11_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2506_ _0351_ _0367_ _0368_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[7\]
+ sky130_fd_sc_hd__nor3_1
X_2437_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[31\]
+ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2368_ _1768_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[22\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_47_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2299_ _1719_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[2\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_79_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1972__S net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout70_X net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input28_A addr[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2043__S net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1882__S net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3340_ _1070_ _1174_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1922__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3271_ _1105_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__inv_2
XANTENNA__2279__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2222_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[45\] VGND VGND VPWR VPWR
+ _1644_ sky130_fd_sc_hd__inv_2
X_2153_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] VGND VGND VPWR VPWR _1575_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2084_ net334 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[50\] net91 VGND
+ VGND VPWR VPWR _0227_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_6_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1989__A1 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2986_ _0812_ _0821_ _0814_ _0815_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__or4b_1
XFILLER_0_8_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1937_ net289 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[39\] net100 VGND
+ VGND VPWR VPWR _0086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1868_ net238 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\] net104 VGND
+ VGND VPWR VPWR _0020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3607_ _1070_ _1441_ VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1799_ _1575_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[53\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\]
+ _1573_ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__o22a_1
X_3538_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[22\] _1369_ _1372_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\]
+ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__o22a_1
XANTENNA__1913__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3469_ _1019_ _1054_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1967__S net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1904__A1 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2038__S net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1877__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2840_ _0489_ _0672_ _0498_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2396__A1 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2771_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[58\]
+ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold117 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[54\] VGND VGND VPWR VPWR net321
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold106 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[57\] VGND VGND VPWR VPWR net310
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold128 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[15\] VGND VGND VPWR VPWR net332
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3323_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[63\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\]
+ VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__nand2b_1
X_3254_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] _1659_ VGND VGND VPWR
+ VPWR _1089_ sky130_fd_sc_hd__and2_1
X_2205_ net106 VGND VGND VPWR VPWR _1627_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3185_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[39\]
+ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__nand2_1
X_4001__196 VGND VGND VPWR VPWR _4001__196/HI net196 sky130_fd_sc_hd__conb_1
X_2136_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[8\] VGND VGND VPWR VPWR _1558_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout165_A net169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2067_ net247 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[33\] net92 VGND
+ VGND VPWR VPWR _0210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1831__B1 _1671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2969_ _0761_ _0800_ _0804_ _0609_ _0605_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_29_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout78_A _1537_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2647__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input50_X net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3941_ clknet_leaf_38_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[18\]
+ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3872_ clknet_leaf_6_CLK _0198_ net155 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2823_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[17\] _1642_ _0571_ _0577_
+ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__a22o_1
X_2754_ _0587_ _0588_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2685_ _1600_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[35\] VGND VGND VPWR
+ VPWR _0521_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3306_ _1584_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[58\] _1140_ _1582_
+ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__o22a_1
X_3237_ _1562_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[44\] VGND VGND VPWR
+ VPWR _1072_ sky130_fd_sc_hd__nand2_1
X_3168_ _1000_ _1002_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__and2_1
X_2119_ net233 net37 net84 VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout168_X net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3099_ _1629_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[61\] VGND VGND VPWR
+ VPWR _0935_ sky130_fd_sc_hd__nand2_1
XANTENNA__3298__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout78 _1537_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1980__S net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input10_A addr[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_31_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3993__188 VGND VGND VPWR VPWR _3993__188/HI net188 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_56_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload26 clknet_leaf_7_CLK VGND VGND VPWR VPWR clkload26/Y sky130_fd_sc_hd__inv_6
XFILLER_0_23_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload15 clknet_leaf_27_CLK VGND VGND VPWR VPWR clkload15/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_35_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload37 clknet_leaf_18_CLK VGND VGND VPWR VPWR clkload37/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__2051__S net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2470_ _1608_ net115 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] _1626_
+ _0324_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__a221o_1
XANTENNA__1890__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3022_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[13\] _0855_ _0857_ VGND VGND VPWR
+ VPWR _0858_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3924_ clknet_leaf_33_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[1\] net140
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3855_ clknet_leaf_21_CLK _0181_ net163 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[36\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload9 clknet_leaf_40_CLK VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_6_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2806_ _0639_ _0640_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\] VGND VGND VPWR
+ VPWR _0642_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout128_A net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3786_ clknet_leaf_24_CLK _0112_ net159 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2737_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[50\]
+ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2668_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[11\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[43\]
+ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__xor2_4
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2599_ _1598_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[2\] _0433_ _0435_
+ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__a211o_1
XANTENNA_input2_A addr[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1975__S net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input58_A wdata[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2046__S net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1970_ net278 net61 net75 VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1885__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3640_ clknet_leaf_1_CLK _0000_ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_3571_ _1404_ _1405_ VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2522_ net113 net112 _0375_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2453_ _1617_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] _1621_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[24\]
+ _0321_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__a221o_1
X_2384_ net72 _1778_ _1779_ VGND VGND VPWR VPWR _1780_ sky130_fd_sc_hd__or3_1
Xinput2 addr[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_67_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3005_ _0792_ _0793_ _0794_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3907_ clknet_leaf_5_CLK _0233_ net154 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[56\]
+ sky130_fd_sc_hd__dfrtp_2
X_3838_ clknet_leaf_7_CLK _0164_ net156 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_37_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_37_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3769_ clknet_leaf_14_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[16\]
+ net165 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_14_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_28_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3999__194 VGND VGND VPWR VPWR _3999__194/HI net194 sky130_fd_sc_hd__conb_1
XFILLER_0_88_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3767__RESET_B net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1953_ net314 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\] net98 VGND
+ VGND VPWR VPWR _0102_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_19_CLK clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_19_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1884_ net329 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] net103 VGND
+ VGND VPWR VPWR _0036_ sky130_fd_sc_hd__mux2_1
X_3623_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[15\] _1657_ VGND VGND VPWR VPWR
+ _1458_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3554_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] _1379_ _1380_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[18\]
+ VGND VGND VPWR VPWR _1389_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3485_ _1287_ _1312_ _1314_ _1104_ _1098_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2505_ net116 _0362_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\] VGND VGND VPWR
+ VPWR _0368_ sky130_fd_sc_hd__a21oi_1
X_2436_ _1590_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[29\] _0305_ VGND
+ VGND VPWR VPWR _0306_ sky130_fd_sc_hd__o21ba_1
X_2367_ net72 _1766_ _1767_ VGND VGND VPWR VPWR _1768_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2298_ net71 _1717_ _1718_ VGND VGND VPWR VPWR _1719_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3270_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[50\]
+ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__xor2_4
X_2221_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[48\] VGND VGND VPWR VPWR
+ _1643_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_8_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_8_CLK sky130_fd_sc_hd__clkbuf_8
X_2152_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] VGND VGND VPWR VPWR
+ _1574_ sky130_fd_sc_hd__inv_2
X_2083_ net277 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[49\] net91 VGND
+ VGND VPWR VPWR _0226_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2985_ _0818_ _0820_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__nand2_1
X_1936_ net223 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[38\] net100 VGND
+ VGND VPWR VPWR _0085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1867_ net240 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\] net104 VGND
+ VGND VPWR VPWR _0019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3606_ _1068_ _1437_ _1066_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__a21oi_1
X_1798_ _1484_ _1486_ VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__nand2_1
Xinput60 wdata[4] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_2
X_4006__201 VGND VGND VPWR VPWR _4006__201/HI net201 sky130_fd_sc_hd__conb_1
X_3537_ _1003_ _1371_ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__xnor2_1
X_3468_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[39\]
+ _1023_ _1302_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__a211o_1
X_3399_ _1232_ _1233_ _1231_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__and3b_1
X_2419_ _1568_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[18\] VGND VGND VPWR
+ VPWR _0289_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2929__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1983__S net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input40_A wdata[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2054__S net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2770_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[58\]
+ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__nor2_1
XANTENNA__1893__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold107 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[28\] VGND VGND VPWR VPWR net311
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold129 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[20\] VGND VGND VPWR VPWR net333
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[57\] VGND VGND VPWR VPWR net322
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3322_ _1592_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[62\] _1145_ _1155_
+ _1154_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__a221o_1
X_3253_ _1079_ _1086_ _1087_ _1072_ _1073_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__a221o_1
X_3184_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[39\]
+ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__nor2_1
X_2204_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[26\] VGND VGND VPWR VPWR _1626_
+ sky130_fd_sc_hd__inv_2
X_2135_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\] VGND VGND VPWR VPWR
+ _1557_ sky130_fd_sc_hd__inv_2
X_2066_ net291 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[32\] net92 VGND
+ VGND VPWR VPWR _0209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout158_A net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1831__A1 _1594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2968_ _0597_ _0600_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1919_ net249 net48 net78 VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2899_ net108 _0653_ _0655_ net107 _0733_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1898__A1 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1978__S net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3478__B _1312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_5_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1889__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input43_X net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2049__S net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3940_ clknet_leaf_39_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[17\]
+ net131 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__1888__S net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3871_ clknet_leaf_7_CLK _0197_ net156 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2822_ _0656_ _0657_ _0651_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2753_ _0587_ _0588_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2684_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[36\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\]
+ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_41_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3305_ _1653_ _1135_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3236_ _1061_ _1065_ _1069_ _1070_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__and4bb_1
X_3167_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[54\]
+ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__or2_1
X_3098_ _1629_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[61\] _1635_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\]
+ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__a2bb2o_1
X_2118_ net218 net36 net84 VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2049_ net269 net41 net86 VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__mux2_1
XANTENNA__2057__A1 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout79 _1537_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_4
XFILLER_0_91_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout90_A _1544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2048__A1 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload16 clknet_leaf_28_CLK VGND VGND VPWR VPWR clkload16/Y sky130_fd_sc_hd__inv_6
Xclkload27 clknet_leaf_8_CLK VGND VGND VPWR VPWR clkload27/Y sky130_fd_sc_hd__clkinv_4
Xclkload38 clknet_leaf_19_CLK VGND VGND VPWR VPWR clkload38/Y sky130_fd_sc_hd__inv_8
XFILLER_0_50_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3021_ net112 _0855_ _0856_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[12\] VGND VGND
+ VPWR VPWR _0857_ sky130_fd_sc_hd__a22o_1
XANTENNA__2039__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3923_ clknet_leaf_33_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[0\] net140
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_46_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3854_ clknet_leaf_22_CLK _0180_ net162 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2805_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\] _0639_ _0640_ _0634_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\]
+ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3785_ clknet_leaf_18_CLK net318 net167 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.pwm_out
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2736_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[50\]
+ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2667_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[11\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[43\]
+ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2598_ _1606_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[7\] _0421_ _0422_
+ _0434_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3219_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[40\]
+ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__xor2_2
XFILLER_0_69_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2660__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1991__S net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout93_X net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2992__A2 _0798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3570_ _1395_ _1397_ _1559_ VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__a21o_1
XANTENNA__2062__S net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2521_ net113 _0375_ net112 VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2452_ _1595_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[0\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\]
+ _1605_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__a2bb2o_1
X_2383_ net118 _1776_ VGND VGND VPWR VPWR _1779_ sky130_fd_sc_hd__and2_1
XANTENNA__2298__A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 addr[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_67_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3004_ _0835_ _0838_ _0839_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_39_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3906_ clknet_leaf_6_CLK _0232_ net155 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[55\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3837_ clknet_leaf_7_CLK _0163_ net156 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3768_ clknet_leaf_13_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[15\]
+ net165 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[15\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_clkbuf_leaf_30_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2719_ _0553_ _0554_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__nor2_2
XFILLER_0_100_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3699_ clknet_leaf_25_CLK _0059_ net144 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1986__S net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2390__B myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_25_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2057__S net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2414__B2 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2414__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1952_ net249 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\] net98 VGND
+ VGND VPWR VPWR _0101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1883_ net327 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] net103 VGND
+ VGND VPWR VPWR _0035_ sky130_fd_sc_hd__mux2_1
X_3622_ _1346_ _1453_ _1455_ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3553_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] _1385_ _1386_ net121 _1380_
+ VGND VGND VPWR VPWR _1388_ sky130_fd_sc_hd__o32a_1
X_3484_ _1096_ _1102_ _1318_ _1095_ VGND VGND VPWR VPWR _1319_ sky130_fd_sc_hd__o211a_1
X_2504_ net116 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\] _0362_ VGND VGND VPWR
+ VPWR _0367_ sky130_fd_sc_hd__and3_1
X_2435_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] _1780_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[29\]
+ _1590_ _0304_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__a221o_1
X_2366_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[22\]
+ _1761_ VGND VGND VPWR VPWR _1767_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2297_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\] _1714_ VGND VGND VPWR VPWR _1718_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2102__B1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2491__A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2653__A_N myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3823__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3733__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2220_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[49\] VGND VGND VPWR VPWR
+ _1642_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2151_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR _1573_
+ sky130_fd_sc_hd__inv_2
X_2082_ net269 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\] net91 VGND
+ VGND VPWR VPWR _0225_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2984_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\] _0816_ _0817_ _0819_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\]
+ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__a32o_1
XFILLER_0_8_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1935_ net217 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[37\] net100 VGND
+ VGND VPWR VPWR _0084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1866_ net244 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] net104 VGND
+ VGND VPWR VPWR _0018_ sky130_fd_sc_hd__mux2_1
X_3605_ _1394_ _1436_ _1438_ _1564_ _1439_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__a221o_1
X_1797_ _1577_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[54\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[53\]
+ _1575_ _1485_ VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__a221oi_1
Xinput61 wdata[5] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput50 wdata[24] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_2
X_3536_ _1116_ _1365_ VGND VGND VPWR VPWR _1371_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout103_A _1535_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3467_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[38\]
+ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[37\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\]
+ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__o211a_1
X_3398_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] _1228_ VGND VGND VPWR VPWR
+ _1233_ sky130_fd_sc_hd__or2_1
X_2418_ _0276_ _0279_ _0285_ _0287_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__or4b_1
X_2349_ _1754_ _1755_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[16\]
+ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input33_A nRST VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold108 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[23\] VGND VGND VPWR VPWR net312
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2070__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold119 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[29\] VGND VGND VPWR VPWR net323
+ sky130_fd_sc_hd__dlygate4sd3_1
X_3321_ _1592_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[62\] _1145_ _1155_
+ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3252_ _1561_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[43\] VGND VGND VPWR
+ VPWR _1087_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_13_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3183_ _1578_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[55\] _1014_ _1017_
+ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__o31a_1
X_2203_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND VPWR VPWR
+ _1625_ sky130_fd_sc_hd__inv_2
X_2134_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[7\] VGND VGND VPWR VPWR _1556_ sky130_fd_sc_hd__inv_2
X_2065_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.rollover_flag myPWM.g_pwm_channel\[1\].CHANNEL.data_mod\[1\]
+ VGND VGND VPWR VPWR _1544_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_22_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2967_ _0761_ _0800_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2898_ _0658_ _0732_ _0733_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__and3_1
X_1918_ net290 net47 net78 VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1849_ net333 net46 net81 VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Left_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3519_ _1350_ _1351_ _1587_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1994__S net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input36_X net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3870_ clknet_leaf_7_CLK _0196_ net156 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2292__C myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2821_ net107 _0655_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2752_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[53\]
+ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2683_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[36\]
+ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3304_ _1588_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[60\] _1138_ VGND
+ VGND VPWR VPWR _1139_ sky130_fd_sc_hd__o21a_1
X_3235_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\]
+ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__xnor2_2
XANTENNA__2829__A1 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_3166_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[54\]
+ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout170_A net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3097_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\] _1634_ _0932_ VGND VGND VPWR
+ VPWR _0933_ sky130_fd_sc_hd__o21a_1
X_2117_ net326 net35 net83 VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2048_ net294 net40 net87 VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout69 net70 VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3999_ net194 VGND VGND VPWR VPWR rdata[22] sky130_fd_sc_hd__buf_2
XFILLER_0_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3831__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout83_A _1534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1989__S net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload17 clknet_leaf_30_CLK VGND VGND VPWR VPWR clkload17/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload28 clknet_leaf_9_CLK VGND VGND VPWR VPWR clkload28/Y sky130_fd_sc_hd__clkinv_8
Xclkload39 clknet_leaf_20_CLK VGND VGND VPWR VPWR clkload39/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_23_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1899__S net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3020_ _0487_ _0785_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3922_ clknet_leaf_40_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.rollover_flag_c net130
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.rollover_flag sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3853_ clknet_leaf_23_CLK _0179_ net160 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2804_ _0624_ _0625_ _0638_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3784_ clknet_leaf_2_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[31\] net153
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2735_ _0570_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__inv_2
X_2666_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[11\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[43\]
+ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__or2_1
XANTENNA__2759__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2597_ _1596_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[1\] VGND VGND VPWR
+ VPWR _0434_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3218_ _1557_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[40\] _1052_ _1555_
+ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__o22a_1
X_3149_ net108 _1639_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[48\] _1616_
+ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_53_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_4_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3826__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout86_X net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2520_ net113 _0375_ _0377_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[12\]
+ sky130_fd_sc_hd__a21oi_1
X_2451_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] _1611_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\]
+ _1619_ _0319_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__a221o_1
X_2382_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[27\] _1776_ VGND VGND VPWR VPWR
+ _1778_ sky130_fd_sc_hd__nor2_1
Xinput4 addr[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
XANTENNA__3457__B2 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3003_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] _0831_ _0834_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[22\]
+ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3905_ clknet_leaf_6_CLK _0231_ net156 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[54\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__1929__Y _1538_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3836_ clknet_leaf_8_CLK _0162_ net157 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\]
+ sky130_fd_sc_hd__dfrtp_4
X_3767_ clknet_leaf_13_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[14\]
+ net165 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[14\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2718_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[41\]
+ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_5_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3983__178 VGND VGND VPWR VPWR _3983__178/HI net178 sky130_fd_sc_hd__conb_1
X_3698_ clknet_leaf_25_CLK _0058_ net147 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2649_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[13\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[45\]
+ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2120__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2671__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input63_A wdata[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2111__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1951_ net290 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[53\] net99 VGND
+ VGND VPWR VPWR _0100_ sky130_fd_sc_hd__mux2_1
XANTENNA__2073__S net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1882_ net333 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] net103 VGND
+ VGND VPWR VPWR _0034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3621_ _1345_ _1364_ _1342_ VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__a21oi_1
X_3552_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] _1383_ _1384_ _1382_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[16\]
+ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__a32o_1
XANTENNA__3776__RESET_B net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1925__A1 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2503_ net116 _0362_ _0366_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[6\]
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__3705__RESET_B net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3483_ _1098_ _1104_ _1317_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__or3_1
X_2434_ _1586_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[27\] _0269_ _0302_
+ _0303_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__a2111o_1
X_2365_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[22\] _1764_ VGND VGND VPWR VPWR
+ _1766_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_87_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2296_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[0\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[1\]
+ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable
+ VGND VGND VPWR VPWR _1717_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2772__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_96_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3819_ clknet_leaf_18_CLK _0145_ net167 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1916__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3108__A myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1907__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2857__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2150_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] VGND VGND VPWR VPWR
+ _1572_ sky130_fd_sc_hd__inv_2
X_2081_ net294 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[47\] net92 VGND
+ VGND VPWR VPWR _0224_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2068__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2983_ _0622_ _0808_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1934_ net212 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[36\] net100 VGND
+ VGND VPWR VPWR _0083_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_44_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1865_ net254 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[3\] net104 VGND
+ VGND VPWR VPWR _0017_ sky130_fd_sc_hd__mux2_1
Xinput40 wdata[15] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_2
X_3604_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\] _1393_ VGND VGND VPWR VPWR
+ _1439_ sky130_fd_sc_hd__nor2_1
X_1796_ _1579_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[55\] VGND VGND VPWR
+ VPWR _1485_ sky130_fd_sc_hd__and2_1
Xinput62 wdata[6] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_2
Xinput51 wdata[25] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_2
X_3535_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\] _1368_ _1369_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[22\]
+ VGND VGND VPWR VPWR _1370_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3466_ _1021_ _1054_ _1300_ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2417_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] _1747_ _1753_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\]
+ _0286_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__o221a_1
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3397_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] _1230_ VGND VGND VPWR VPWR
+ _1232_ sky130_fd_sc_hd__nor2_1
XANTENNA__2767__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2348_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[16\] _1752_ _1713_ VGND VGND VPWR
+ VPWR _1755_ sky130_fd_sc_hd__o21ai_1
X_2279_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\]
+ VGND VGND VPWR VPWR _1701_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3989__184 VGND VGND VPWR VPWR _3989__184/HI net184 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_10_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3834__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2677__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input26_A addr[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2250__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold109 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[60\] VGND VGND VPWR VPWR net313
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3320_ _1592_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[62\] _1146_ VGND
+ VGND VPWR VPWR _1155_ sky130_fd_sc_hd__o21a_1
XFILLER_0_95_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3251_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] _1662_ _1085_ VGND
+ VGND VPWR VPWR _1086_ sky130_fd_sc_hd__o21a_1
X_3182_ _1006_ _1015_ _1580_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[56\]
+ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__o2bb2a_1
X_2202_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] VGND VGND VPWR VPWR _1624_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2133_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] VGND VGND VPWR VPWR
+ _1555_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2064_ net281 net58 net85 VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3919__Q myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_2966_ _0761_ _0796_ _0798_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2897_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[22\] _0650_ VGND VGND VPWR VPWR
+ _0733_ sky130_fd_sc_hd__or2_1
X_1917_ net296 net46 net77 VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1848_ net293 net44 net82 VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3518_ _1129_ _1348_ VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__xnor2_1
X_3449_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[46\]
+ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2820_ net108 _0653_ _0655_ net107 VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_5_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2751_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[53\]
+ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__or2_1
XANTENNA__2081__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2682_ _1604_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[38\] VGND VGND VPWR
+ VPWR _0518_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3303_ _1586_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[59\] _1125_ VGND
+ VGND VPWR VPWR _1138_ sky130_fd_sc_hd__or3_1
X_3234_ _1066_ _1067_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__or2_2
X_3165_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[54\]
+ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__nand2_1
X_3096_ _1632_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[63\] VGND VGND VPWR
+ VPWR _0932_ sky130_fd_sc_hd__nand2_1
X_2116_ net214 net65 net84 VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__mux2_1
X_2047_ net283 net39 net87 VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3998_ net193 VGND VGND VPWR VPWR rdata[21] sky130_fd_sc_hd__buf_2
XANTENNA__2780__A _1623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2949_ _0782_ _0784_ _0767_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout76_A _1540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2453__B1 _1621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload29 clknet_leaf_10_CLK VGND VGND VPWR VPWR clkload29/Y sky130_fd_sc_hd__inv_8
Xclkload18 clknet_leaf_31_CLK VGND VGND VPWR VPWR clkload18/Y sky130_fd_sc_hd__inv_6
XFILLER_0_23_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2201__Y _1623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2076__S net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3921_ clknet_leaf_21_CLK _0247_ net163 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.alignment
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3852_ clknet_leaf_21_CLK _0178_ net162 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2803_ _0624_ _0625_ _0638_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__nand3_1
X_3783_ clknet_leaf_12_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[30\]
+ net153 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[30\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2734_ _0552_ _0557_ _0569_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_41_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2665_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[11\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[43\]
+ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__nor2_1
X_2596_ _1604_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[6\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[7\]
+ _1606_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_10_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3217_ _1557_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[40\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[39\]
+ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__a21o_1
X_3148_ _1616_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[48\] _0944_ _0949_
+ _0958_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__a2111o_1
X_3079_ _0607_ _0913_ _0600_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_53_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3842__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout79_X net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3894__RESET_B net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2450_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\]
+ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__xor2_1
XFILLER_0_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2381_ _1776_ _1777_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[26\]
+ sky130_fd_sc_hd__nor2_1
Xinput5 addr[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3002_ net107 _0833_ _0837_ net108 VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_36_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3904_ clknet_leaf_6_CLK _0230_ net156 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[53\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3835_ clknet_leaf_8_CLK _0161_ net157 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_74_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3766_ clknet_leaf_13_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[13\]
+ net165 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2717_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[41\]
+ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__nor2_1
X_3697_ clknet_leaf_25_CLK _0057_ net147 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2648_ _0482_ _0483_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__nand2_2
XANTENNA__3662__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2579_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[20\]
+ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__xor2_1
XFILLER_0_100_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2399__B myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input56_A wdata[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1870__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1950_ net296 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\] net99 VGND
+ VGND VPWR VPWR _0099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1881_ net293 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] net103 VGND
+ VGND VPWR VPWR _0033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3620_ _1352_ _1363_ _1454_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3551_ _1099_ _1381_ _1106_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2502_ net116 _0362_ net70 VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3482_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[50\]
+ _1316_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2433_ _1582_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[25\] VGND VGND VPWR
+ VPWR _0303_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3127__B2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_3_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2364_ _1765_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[21\]
+ sky130_fd_sc_hd__inv_2
X_2295_ _1716_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[1\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3818_ clknet_leaf_23_CLK _0144_ net159 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout129_X net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3749_ clknet_leaf_42_CLK _0109_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[62\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_30_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1852__A1 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap89 _1543_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
XFILLER_0_77_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2203__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input59_X net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_467 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2080_ net283 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[46\] net92 VGND
+ VGND VPWR VPWR _0223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2084__S net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2982_ _0816_ _0817_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\] VGND VGND VPWR
+ VPWR _0818_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3596__B2 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1933_ net210 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[35\] net100 VGND
+ VGND VPWR VPWR _0082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3603_ _1069_ _1437_ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__xnor2_1
Xinput30 addr[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1864_ net232 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\] net104 VGND
+ VGND VPWR VPWR _0016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput41 wdata[16] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
X_1795_ _1579_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[55\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[54\]
+ _1577_ VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__o22a_1
Xinput63 wdata[7] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_2
Xinput52 wdata[26] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_2
XANTENNA__3209__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3534_ _1011_ _1366_ VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__xnor2_1
XANTENNA__2020__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3465_ _1025_ _1045_ VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2416_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] _1747_ _1750_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\]
+ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__o2bb2a_1
X_3396_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] _1228_ _1230_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\]
+ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__a22oi_1
X_2347_ net122 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[16\] _1749_ VGND VGND VPWR
+ VPWR _1754_ sky130_fd_sc_hd__and3_1
XANTENNA__3940__Q myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2278_ _1693_ _1695_ _1697_ _1699_ VGND VGND VPWR VPWR _1700_ sky130_fd_sc_hd__and4_1
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2011__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3667__RESET_B net144 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input19_A addr[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_2_0__f_CLK_X clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2250__B2 _1560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2250__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3029__A net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3250_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] _1662_ _1663_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\]
+ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__a22o_1
XANTENNA__2079__S net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3181_ _1578_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[55\] VGND VGND VPWR
+ VPWR _1016_ sky130_fd_sc_hd__nor2_1
X_2201_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[25\] VGND VGND VPWR VPWR
+ _1623_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2132_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] VGND VGND VPWR VPWR
+ _1554_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2063_ net292 net57 net85 VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2965_ _0799_ _0761_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__and2b_1
XFILLER_0_56_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2896_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] _0649_ VGND VGND VPWR VPWR
+ _0732_ sky130_fd_sc_hd__or2_1
X_1916_ net302 net44 net78 VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1847_ net320 net43 net82 VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3517_ _1587_ _1350_ _1351_ VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3448_ _1003_ _1010_ _1014_ _1119_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__and4_1
X_3379_ _1212_ _1213_ _1185_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3845__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_43_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2750_ _0570_ _0579_ _0585_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__o21a_2
X_2681_ _0513_ _0516_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__and2b_1
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3302_ _1125_ _1128_ _1136_ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__or3b_1
X_3233_ _1066_ _1067_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__nor2_1
X_3164_ _1576_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[54\] VGND VGND VPWR
+ VPWR _0999_ sky130_fd_sc_hd__nor2_1
X_3095_ _0930_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__inv_2
X_2115_ net236 net64 net84 VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__mux2_1
X_2046_ net274 net38 net88 VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout156_A net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3997_ net192 VGND VGND VPWR VPWR rdata[20] sky130_fd_sc_hd__buf_2
XFILLER_0_91_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3941__RESET_B net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2948_ _0500_ _0504_ _0783_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2879_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\] _0682_ _0713_ _0714_ VGND VGND
+ VPWR VPWR _0715_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_32_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_584 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2301__A net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout69_A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload19 clknet_leaf_33_CLK VGND VGND VPWR VPWR clkload19/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input41_X net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3920_ clknet_leaf_21_CLK _0246_ net163 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.polarity
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3851_ clknet_leaf_23_CLK _0177_ net160 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2092__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3782_ clknet_leaf_11_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[29\]
+ net153 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] sky130_fd_sc_hd__dfrtp_4
X_2802_ _0635_ _0636_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__nand2b_1
X_2733_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[16\] _1643_ _0495_ _0568_
+ _0564_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2664_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[44\]
+ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__xor2_2
X_2595_ _0428_ _0431_ _0430_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__or3b_1
XANTENNA__2380__B1 _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3216_ _1021_ _1049_ _1050_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_19_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3147_ _0961_ _0962_ _0964_ _0982_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__o22a_1
XFILLER_0_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3078_ _0601_ _0606_ _0913_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_53_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2435__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2029_ net309 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\] net94 VGND
+ VGND VPWR VPWR _0175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Left_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2206__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2380_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[26\] _1774_ _1713_ VGND VGND VPWR
+ VPWR _1777_ sky130_fd_sc_hd__o21ai_1
Xinput6 addr[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XANTENNA__2087__S net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3001_ _0828_ _0836_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2417__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3903_ clknet_leaf_7_CLK _0229_ net170 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_86_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3834_ clknet_leaf_15_CLK _0160_ net166 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3765_ clknet_leaf_14_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[12\]
+ net165 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2716_ _0512_ _0549_ _0551_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__and3_1
X_3696_ clknet_leaf_25_CLK _0056_ net148 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2647_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\]
+ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__nand2_1
XANTENNA__2353__B1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2578_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[31\] VGND VGND VPWR VPWR
+ _0416_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout91_X net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input49_A wdata[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1880_ net320 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] net102 VGND
+ VGND VPWR VPWR _0032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3550_ _1099_ _1106_ _1381_ VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2501_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[5\] VGND VGND VPWR VPWR
+ _0365_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3481_ _1568_ _1654_ _1099_ VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2432_ _0273_ _0299_ _0300_ _0301_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2363_ net72 _1763_ _1764_ VGND VGND VPWR VPWR _1765_ sky130_fd_sc_hd__or3_1
X_2294_ net71 _1714_ _1715_ VGND VGND VPWR VPWR _1716_ sky130_fd_sc_hd__or3_1
XFILLER_0_79_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3714__RESET_B net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3817_ clknet_leaf_2_CLK _0143_ net153 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_3748_ clknet_leaf_42_CLK _0108_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[61\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_70_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3673__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3679_ clknet_leaf_43_CLK _0039_ net128 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_100_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2981_ _0621_ _0637_ _0809_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__nand3_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1932_ net224 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[34\] net100 VGND
+ VGND VPWR VPWR _0081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1863_ net307 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\] net104 VGND
+ VGND VPWR VPWR _0015_ sky130_fd_sc_hd__mux2_1
X_3602_ _1061_ _1065_ _1309_ _1285_ VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__a31o_1
Xinput20 addr[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_1
Xinput31 addr[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
Xinput42 wdata[17] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
X_1794_ _1479_ _1482_ _1458_ _1464_ VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__o2bb2a_1
Xinput53 wdata[27] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput64 wdata[8] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_0_CLK_A CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3533_ _1014_ _1367_ VGND VGND VPWR VPWR _1368_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3464_ _1031_ _1196_ _1296_ _1298_ VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__a31o_1
X_2415_ _0280_ _0281_ _0282_ _0284_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__or4b_1
XFILLER_0_58_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3225__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3395_ _1003_ _1229_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__xnor2_1
X_2346_ _1753_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[15\]
+ sky130_fd_sc_hd__inv_2
X_2277_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] _1567_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\]
+ _1581_ _1698_ VGND VGND VPWR VPWR _1699_ sky130_fd_sc_hd__o221a_1
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1834__A2 _1521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3668__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2304__A net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout99_A _1538_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_2_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2200_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[24\] VGND VGND VPWR VPWR _1622_
+ sky130_fd_sc_hd__inv_2
X_3180_ _1010_ _1014_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__nor2_1
X_2131_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] VGND VGND VPWR VPWR
+ _1553_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2062_ net331 net55 net85 VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2095__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2964_ _0796_ _0798_ _0799_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_84_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1915_ net211 net43 net78 VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2895_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[19\] _0668_ VGND VGND VPWR VPWR
+ _0731_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1846_ _1533_ net26 net66 VGND VGND VPWR VPWR _1534_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3516_ _1126_ _1349_ _1125_ VGND VGND VPWR VPWR _1351_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout101_A _1538_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3447_ _1008_ _1013_ _1281_ _1012_ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__a31o_1
X_3378_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[10\] _1182_ _1187_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[9\]
+ VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__o22ai_1
XANTENNA__3139__A1_N net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2329_ net124 _1739_ VGND VGND VPWR VPWR _1741_ sky130_fd_sc_hd__nor2_1
XANTENNA__1902__S net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3995__190 VGND VGND VPWR VPWR _3995__190/HI net190 sky130_fd_sc_hd__conb_1
XFILLER_0_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1991__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3496__A1 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input31_A addr[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2680_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[39\]
+ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__xnor2_2
XANTENNA__1982__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3301_ _1132_ _1135_ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__and2_1
X_3232_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[47\]
+ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__nor2_1
X_3163_ _0996_ _0997_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__and2_2
X_3979__174 VGND VGND VPWR VPWR _3979__174/HI net174 sky130_fd_sc_hd__conb_1
X_2114_ net273 net63 net83 VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__mux2_1
X_3094_ _1632_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[63\] _1634_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\]
+ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__a2bb2o_1
X_2045_ net303 net37 net88 VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3996_ net191 VGND VGND VPWR VPWR rdata[19] sky130_fd_sc_hd__buf_2
XANTENNA_fanout149_A net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2947_ _0509_ _0555_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1973__A1 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2878_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\] _0682_ _0711_ net114 VGND VGND
+ VPWR VPWR _0714_ sky130_fd_sc_hd__a22oi_1
XANTENNA__1964__Y _1540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1829_ _1503_ _1509_ _1516_ VGND VGND VPWR VPWR _1518_ sky130_fd_sc_hd__or3b_1
XFILLER_0_13_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout104_X net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3681__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3413__A _1094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2453__A2 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_90_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2699__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3651__RESET_B net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input34_X net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3850_ clknet_leaf_2_CLK _0176_ net153 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_mod\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3781_ clknet_leaf_11_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[28\]
+ net153 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[28\] sky130_fd_sc_hd__dfrtp_4
X_2801_ _0635_ _0636_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2732_ _0489_ _0498_ _0566_ _0567_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__a31o_1
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2663_ _0488_ _0491_ _0495_ _0498_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__nand4_1
XFILLER_0_22_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2594_ _1609_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[9\] VGND VGND VPWR
+ VPWR _0431_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3215_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] _1664_ VGND VGND VPWR
+ VPWR _1050_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3146_ net112 _1644_ _1645_ net113 _0981_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__a221oi_2
X_3077_ _0605_ _0801_ _0802_ _0608_ _0604_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__o311ai_2
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2028_ net279 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\] net94 VGND
+ VGND VPWR VPWR _0174_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3676__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3979_ net174 VGND VGND VPWR VPWR rdata[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_33_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_42_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2031__B net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout81_A _1534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2123__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2114__A1 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput7 addr[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
X_3000_ _0590_ _0796_ _0798_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__nand3_1
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3902_ clknet_leaf_7_CLK _0228_ net156 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[51\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3833_ clknet_leaf_12_CLK _0159_ net161 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_27_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3764_ clknet_leaf_13_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[11\]
+ net165 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__1928__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2715_ _0519_ _0533_ _0550_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__nand3_1
X_3695_ clknet_leaf_27_CLK _0055_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3228__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2132__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2646_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\]
+ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2577_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[31\] _0413_ _0415_ _0351_ VGND VGND
+ VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[31\] sky130_fd_sc_hd__a211oi_2
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2105__A1 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3129_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[37\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\]
+ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_38_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1910__S net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1919__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2592__B2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout84_X net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_1_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2280__B1 _1592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2032__B1 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3480_ _1287_ _1312_ _1314_ VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2500_ net70 _0363_ _0364_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[5\]
+ sky130_fd_sc_hd__and3_1
X_2431_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] _1765_ VGND VGND VPWR
+ VPWR _0301_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_47_Left_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2362_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\]
+ _1760_ VGND VGND VPWR VPWR _1764_ sky130_fd_sc_hd__and3_1
X_2293_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[0\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable
+ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[1\] VGND VGND VPWR VPWR _1715_ sky130_fd_sc_hd__a21oi_1
X_4004__199 VGND VGND VPWR VPWR _4004__199/HI net199 sky130_fd_sc_hd__conb_1
XFILLER_0_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout131_A net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3816_ clknet_leaf_3_CLK _0142_ net151 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_3747_ clknet_leaf_42_CLK _0107_ net128 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_65_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3678_ clknet_leaf_43_CLK _0038_ net133 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2629_ _0463_ _0464_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__and2b_1
XANTENNA__1905__S net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_83_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input61_A wdata[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2500__A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_92_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2980_ _0621_ _0809_ _0637_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1931_ net213 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[33\] net100 VGND
+ VGND VPWR VPWR _0080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1862_ net205 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[0\] net104 VGND
+ VGND VPWR VPWR _0014_ sky130_fd_sc_hd__mux2_1
X_3601_ _1428_ _1431_ _1434_ _1435_ VGND VGND VPWR VPWR _1436_ sky130_fd_sc_hd__o31ai_2
XANTENNA__3774__Q myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xinput10 addr[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
Xinput21 addr[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1793_ _1461_ _1481_ _1480_ _1460_ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__and4b_1
Xinput32 addr[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
Xinput54 wdata[28] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput43 wdata[18] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
X_3532_ _1011_ _1366_ _1008_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__o21ai_1
Xinput65 wdata[9] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_2
X_3463_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[35\]
+ _1196_ _1294_ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__a31o_1
X_2414_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] _1728_ _1730_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\]
+ _0283_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_30_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_30_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3394_ _1115_ _1118_ _1005_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__a21oi_1
X_2345_ net71 _1751_ _1752_ VGND VGND VPWR VPWR _1753_ sky130_fd_sc_hd__or3_1
XFILLER_0_74_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2276_ _1580_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[24\] _1586_ net118 VGND VGND
+ VPWR VPWR _1698_ sky130_fd_sc_hd__o22a_1
XANTENNA__3935__RESET_B net144 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2320__A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_CLK clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_21_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input64_X net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_12_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_12_CLK sky130_fd_sc_hd__clkbuf_8
X_2130_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND VPWR VPWR
+ _1552_ sky130_fd_sc_hd__inv_2
X_2061_ net306 net54 net85 VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2963_ _0466_ _0470_ _0473_ _0589_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_84_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1914_ net267 net42 net78 VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2894_ _0725_ _0727_ _0728_ _0729_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1845_ net12 net1 net23 _1532_ VGND VGND VPWR VPWR _1533_ sky130_fd_sc_hd__or4_2
X_3515_ _1125_ _1126_ _1349_ VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3446_ _1000_ _1116_ _1009_ _1001_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__a211o_1
XFILLER_0_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3377_ _1190_ _1209_ _1210_ _1211_ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__o31a_1
XFILLER_0_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2328_ _1740_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[10\]
+ sky130_fd_sc_hd__inv_2
X_2259_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[14\]
+ VGND VGND VPWR VPWR _1681_ sky130_fd_sc_hd__xor2_1
XFILLER_0_67_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2465__B1 _1623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3679__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input24_A addr[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_1_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3300_ _1133_ _1134_ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3231_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[47\]
+ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__and2_1
X_3162_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[61\]
+ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__or2_1
X_2113_ net238 net62 net83 VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__mux2_1
X_3093_ _0922_ _0926_ _0928_ _0827_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__a31o_1
X_2044_ net259 net36 net88 VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3995_ net190 VGND VGND VPWR VPWR rdata[18] sky130_fd_sc_hd__buf_2
XFILLER_0_57_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2135__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2946_ _0774_ _0775_ _0779_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_20_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2877_ _0707_ _0709_ _0712_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1828_ _1589_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[60\] _1509_ VGND
+ VGND VPWR VPWR _1517_ sky130_fd_sc_hd__or3_1
XFILLER_0_40_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_2_1__f_CLK_A clknet_0_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3429_ net118 _1262_ VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__and2_1
XANTENNA__3950__RESET_B net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_1_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1913__S net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3323__B myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3780_ clknet_leaf_11_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[27\]
+ net154 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[27\] sky130_fd_sc_hd__dfrtp_1
X_2800_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[62\]
+ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__nand2_1
X_2731_ _1614_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\] VGND VGND VPWR
+ VPWR _0567_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2662_ _0496_ _0497_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__nand2_2
XANTENNA__3779__RESET_B net154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3782__Q myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_2593_ _1600_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[3\] _0365_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\]
+ _0429_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__o221a_1
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3214_ _1025_ _1047_ _1022_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3145_ net113 _1645_ _1646_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[11\] _0980_
+ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__o221a_1
XFILLER_0_96_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1891__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3076_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] _0910_ VGND VGND VPWR VPWR
+ _0912_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2027_ net323 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] net94 VGND
+ VGND VPWR VPWR _0173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout161_A net169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3978_ net173 VGND VGND VPWR VPWR rdata[1] sky130_fd_sc_hd__buf_2
XANTENNA__3396__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__3396__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2929_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[42\]
+ _0764_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1908__S net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2966__C _0798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout74_A _1540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3320__A1 _1592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput8 addr[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3901_ clknet_leaf_8_CLK _0227_ net157 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[50\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3832_ clknet_leaf_12_CLK _0158_ net159 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\]
+ sky130_fd_sc_hd__dfrtp_4
X_3763_ clknet_leaf_13_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[10\]
+ net165 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[10\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_30_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2050__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4009__204 VGND VGND VPWR VPWR _4009__204/HI net204 sky130_fd_sc_hd__conb_1
X_2714_ _0517_ _0537_ _0545_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__and3_1
X_3694_ clknet_leaf_26_CLK _0054_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2645_ _0479_ _0480_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__nand2b_2
X_2576_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[31\] _0413_ VGND VGND VPWR VPWR
+ _0415_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3128_ _0963_ _0961_ _0962_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_66_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3059_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[12\] _0856_ VGND VGND VPWR VPWR
+ _0895_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2577__C1 _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2041__A1 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3541__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__3541__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout77_X net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1855__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2280__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2280__B2 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2430_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[17\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[17\]
+ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__xor2_1
X_2361_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] _1761_ VGND VGND VPWR VPWR
+ _1763_ sky130_fd_sc_hd__nor2_1
X_2292_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[0\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[1\]
+ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable VGND VGND VPWR VPWR _1714_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2099__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_41_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2271__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3815_ clknet_leaf_4_CLK _0141_ net150 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2023__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3746_ clknet_leaf_43_CLK _0106_ net128 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[59\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_15_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3677_ clknet_leaf_44_CLK _0037_ net133 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2628_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[24\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[56\]
+ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__nand2_1
X_2559_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[26\]
+ _0399_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1921__S net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2014__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3155__Y _0991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input54_A wdata[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2253__A1 _1570_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1930_ net231 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[32\] net100 VGND
+ VGND VPWR VPWR _0079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1861_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.rollover_flag myPWM.g_pwm_channel\[0\].CHANNEL.data_mod\[0\]
+ VGND VGND VPWR VPWR _1535_ sky130_fd_sc_hd__nand2_2
X_3600_ net123 _1391_ _1430_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] VGND VGND
+ VPWR VPWR _1435_ sky130_fd_sc_hd__o22a_1
XANTENNA__2005__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput11 addr[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput22 addr[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
Xinput33 nRST VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_4
X_1792_ _1560_ net124 _1661_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[42\]
+ VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__or4_1
X_3531_ _1000_ _1116_ _1365_ _1001_ VGND VGND VPWR VPWR _1366_ sky130_fd_sc_hd__a31o_1
Xinput44 wdata[19] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput55 wdata[29] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput66 wen VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_1
XFILLER_0_52_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3462_ _1031_ _1296_ _1030_ VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__a21o_1
X_3393_ _1115_ _1118_ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__xnor2_1
X_2413_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] _1722_ _1735_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\]
+ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_58_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3505__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_2344_ net122 _1749_ VGND VGND VPWR VPWR _1752_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2275_ _1574_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\]
+ _1577_ _1696_ VGND VGND VPWR VPWR _1697_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout127_X net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3729_ clknet_leaf_26_CLK _0089_ net147 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[42\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__1916__S net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2601__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input1_X net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input57_X net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2060_ net282 net53 net85 VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2962_ _0786_ _0787_ _0791_ _0797_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__a31o_2
XFILLER_0_60_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1913_ net330 net41 net78 VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__mux2_1
X_2893_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[15\] _0675_ VGND VGND VPWR VPWR
+ _0729_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1844_ net27 _1531_ VGND VGND VPWR VPWR _1532_ sky130_fd_sc_hd__nand2b_1
XANTENNA__2421__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3514_ _1131_ _1134_ _1347_ _1133_ _1129_ VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__a311o_1
XFILLER_0_4_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3445_ _1168_ _1257_ _1263_ _1274_ _1279_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__a41o_1
XFILLER_0_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3376_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[9\] _1187_ _1189_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[8\]
+ VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__a22oi_1
X_2327_ net71 _1738_ _1739_ VGND VGND VPWR VPWR _1740_ sky130_fd_sc_hd__or3_1
X_2258_ _1673_ _1675_ _1677_ _1679_ VGND VGND VPWR VPWR _1680_ sky130_fd_sc_hd__or4_1
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2465__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2465__B2 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_2189_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\] VGND VGND VPWR VPWR _1611_
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_84_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2331__A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3162__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input17_A addr[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2506__A _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3230_ _1062_ _1064_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__nand2_2
XANTENNA_max_cap89_X net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3161_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[61\]
+ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__nand2_1
X_2112_ net240 net61 net83 VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__mux2_1
X_3092_ _1626_ _0914_ _0915_ _0920_ _0927_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__a311o_1
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2043_ net261 net35 net88 VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3994_ net189 VGND VGND VPWR VPWR rdata[17] sky130_fd_sc_hd__buf_2
X_2945_ _0515_ _0780_ _0514_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2876_ net115 _0706_ _0711_ net114 VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__o22ai_1
X_1827_ net118 _1651_ _1652_ net119 _1515_ VGND VGND VPWR VPWR _1516_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2151__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__3247__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3428_ net118 _1262_ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__or2_1
X_3359_ _1025_ _1047_ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__xnor2_1
XANTENNA_input9_A addr[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2000__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2429__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2236__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[46\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2730_ _0490_ _0565_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2661_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[15\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\]
+ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__nand2_1
X_3985__180 VGND VGND VPWR VPWR _3985__180/HI net180 sky130_fd_sc_hd__conb_1
XANTENNA__3157__A2 _0991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2592_ _1598_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[2\] _0361_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\]
+ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__o22a_1
XFILLER_0_22_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3213_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] _1666_ _1025_ _1022_
+ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3748__RESET_B net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3144_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[11\] _1646_ _1647_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\]
+ _0979_ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__a221o_1
X_3075_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[24\] _0908_ _0910_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\]
+ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2026_ net311 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] net94 VGND
+ VGND VPWR VPWR _0172_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2146__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout154_A net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3977_ net172 VGND VGND VPWR VPWR rdata[0] sky130_fd_sc_hd__buf_2
XFILLER_0_57_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2928_ _0509_ _0554_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2859_ _1595_ _0693_ _0694_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[1\] VGND VGND
+ VPWR VPWR _0695_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_5_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1924__S net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput9 addr[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XANTENNA__3075__B2 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_52_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3900_ clknet_leaf_8_CLK _0226_ net157 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3831_ clknet_leaf_15_CLK _0157_ net166 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3762_ clknet_leaf_13_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[9\] net165
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_0_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3693_ clknet_leaf_29_CLK _0053_ net143 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2713_ _0517_ _0547_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2644_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\]
+ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__nand2_1
X_2575_ _0414_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[30\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3127_ net112 _1644_ _1613_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\]
+ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__3260__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3058_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\] _0871_ _0892_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[11\]
+ _0893_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__a221oi_1
X_2009_ net215 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[11\] net97 VGND
+ VGND VPWR VPWR _0155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2604__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1919__S net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_3__f_CLK_X clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2360_ _1761_ _1762_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[20\]
+ sky130_fd_sc_hd__nor2_1
X_2291_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable _1711_ VGND VGND VPWR VPWR
+ _1713_ sky130_fd_sc_hd__nand2_4
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3814_ clknet_leaf_4_CLK _0140_ net150 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3745_ clknet_leaf_43_CLK _0105_ net133 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[58\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3676_ clknet_leaf_0_CLK _0036_ net135 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3763__RESET_B net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2627_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[24\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[56\]
+ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__nor2_1
X_2558_ _0401_ _0402_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[25\]
+ sky130_fd_sc_hd__nor2_1
X_2489_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[3\] _0354_ VGND VGND VPWR VPWR _0356_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3165__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input47_A wdata[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2509__A _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2253__A2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1860_ net241 net58 net81 VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1791_ net122 _1657_ _1660_ net123 _1463_ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 addr[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_1
Xinput34 wdata[0] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_4
Xinput45 wdata[1] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_2
X_3530_ _1319_ _1320_ _1118_ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__a21o_1
Xinput23 addr[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_1
Xinput56 wdata[2] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3461_ _1034_ _1295_ _1033_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__a21o_1
X_3392_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\] _1226_ VGND VGND VPWR VPWR
+ _1227_ sky130_fd_sc_hd__nor2_1
X_2412_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] _1737_ _1730_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\]
+ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__a2bb2o_1
X_2343_ net122 _1749_ VGND VGND VPWR VPWR _1751_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2274_ _1559_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\]
+ _1551_ VGND VGND VPWR VPWR _1696_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_79_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2154__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1989_ net237 net50 net73 VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3728_ clknet_leaf_25_CLK _0088_ net147 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[41\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_101_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3659_ clknet_leaf_27_CLK _0019_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1932__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2329__A net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1994__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_40_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2003__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2961_ _0481_ _0484_ _0793_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__or3_1
XFILLER_0_84_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1912_ net250 net40 net77 VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1985__A1 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2892_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[16\] _0664_ _0665_ _0663_ VGND VGND
+ VPWR VPWR _0728_ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1843_ _1523_ _1524_ _1525_ _1530_ VGND VGND VPWR VPWR _1531_ sky130_fd_sc_hd__nor4_1
XFILLER_0_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3513_ _1131_ _1134_ _1347_ _1133_ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_73_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3444_ _1168_ _1276_ _1277_ _1278_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__a211o_1
X_3375_ _1556_ _1191_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__and2_1
X_2326_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[9\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[10\]
+ _1734_ VGND VGND VPWR VPWR _1739_ sky130_fd_sc_hd__and3_1
XANTENNA__2149__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_2257_ _1552_ net127 _1572_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] _1678_
+ VGND VGND VPWR VPWR _1679_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2188_ net114 VGND VGND VPWR VPWR _1610_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_84_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1976__A1 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1927__S net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout97_A _1541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1900__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2065__Y _1544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1967__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_89_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3160_ _0993_ _0994_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__and2b_1
Xhold1 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[0\] VGND VGND VPWR VPWR net205
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2111_ net244 net60 net83 VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__mux2_1
X_3091_ _0911_ _0912_ _0916_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[26\] VGND VGND
+ VPWR VPWR _0927_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_55_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2042_ net243 net65 net88 VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3993_ net188 VGND VGND VPWR VPWR rdata[16] sky130_fd_sc_hd__buf_2
X_2944_ _0538_ _0546_ _0774_ _0776_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2875_ _0509_ _0710_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__xor2_1
XFILLER_0_72_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1826_ net119 _1652_ _1653_ net120 _1505_ VGND VGND VPWR VPWR _1515_ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3427_ _1125_ _1261_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3358_ net125 _1192_ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__nand2_1
X_2309_ net127 net126 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\] _1717_ VGND VGND
+ VPWR VPWR _1727_ sky130_fd_sc_hd__and4_1
X_3289_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[60\]
+ VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_28_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2660_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[15\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\]
+ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2591_ _1604_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[6\] _0425_ _0426_
+ _0427_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_10_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3212_ _1027_ _1041_ _1045_ _1026_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2117__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3143_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\] _1647_ _0974_ _0977_ _0978_
+ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3074_ _0609_ _0909_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2025_ net325 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] net94 VGND
+ VGND VPWR VPWR _0171_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3717__RESET_B net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3976_ myPWM.g_pwm_channel\[1\].CHANNEL.pwm_out VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_61_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2927_ _0488_ _0491_ _0762_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2162__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2858_ _0528_ _0529_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__xnor2_1
X_1809_ _1483_ _1494_ _1495_ _1497_ VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__or4_1
X_2789_ _1628_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[61\] VGND VGND VPWR
+ VPWR _0625_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout102_X net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2101__S _1545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2108__A1 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1940__S net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2011__S net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1850__S net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2283__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3830_ clknet_leaf_16_CLK _0156_ net166 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3761_ clknet_leaf_13_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[8\] net161
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2712_ _0518_ _0541_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_30_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3692_ clknet_leaf_28_CLK _0052_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2643_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\]
+ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__nor2_1
X_2574_ _0351_ _0412_ _0413_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__or3_1
XFILLER_0_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3126_ _1615_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\]
+ _1613_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_66_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3057_ _0862_ _0865_ _0871_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\] _0867_
+ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__o221a_1
X_2008_ net253 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] net97 VGND
+ VGND VPWR VPWR _0154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3259__Y _1094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3959_ clknet_leaf_30_CLK _0251_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1935__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3170__B myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2265__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2006__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_42_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_42_CLK sky130_fd_sc_hd__clkbuf_8
X_2290_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable _1711_ VGND VGND VPWR VPWR
+ _1712_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_16_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3813_ clknet_leaf_4_CLK _0139_ net152 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_25_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3744_ clknet_leaf_43_CLK _0104_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[57\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_70_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3675_ clknet_leaf_0_CLK _0035_ net134 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2626_ _0461_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_33_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_33_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2557_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] _0399_ net69 VGND VGND VPWR
+ VPWR _0402_ sky130_fd_sc_hd__o21ai_1
X_2488_ _0354_ _0355_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[2\]
+ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_34_Left_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3109_ _1616_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[48\] _0944_ VGND
+ VGND VPWR VPWR _0945_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_87_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1997__Y _1541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_43_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2406__A1_N myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_CLK clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_24_CLK sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_52_Left_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout82_X net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_439 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1790_ net124 _1661_ _1662_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[10\] _1478_
+ VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput13 addr[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput24 addr[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput35 wdata[10] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_2
Xinput46 wdata[20] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput57 wdata[30] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_15_CLK clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_15_CLK sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_70_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3460_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[32\] _1199_ _1198_ VGND
+ VGND VPWR VPWR _1295_ sky130_fd_sc_hd__a21o_1
X_3391_ _1014_ _1225_ VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__xnor2_1
X_2411_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] _1716_ _1735_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\]
+ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__a2bb2o_1
X_2342_ _1750_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[14\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_20_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2273_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] _1583_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\]
+ _1594_ _1694_ VGND VGND VPWR VPWR _1695_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_550 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1988_ net262 net49 net74 VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3727_ clknet_leaf_27_CLK _0087_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[40\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3658_ clknet_leaf_29_CLK _0018_ net143 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_3589_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\] _1411_ _1423_ net125 VGND VGND
+ VPWR VPWR _1424_ sky130_fd_sc_hd__o22a_1
X_2609_ _0437_ _0438_ _0444_ _0445_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2468__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[24\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2345__A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_4_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_17_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2960_ _0479_ _0483_ _0795_ _0480_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__o211a_1
X_1911_ net209 net39 net79 VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__mux2_1
X_2891_ _0680_ _0721_ _0722_ _0726_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1842_ _1526_ _1527_ _1528_ _1529_ VGND VGND VPWR VPWR _1530_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3512_ _1282_ _1321_ _1132_ VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3443_ _1593_ _1161_ _1162_ _1159_ VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_100_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3374_ _1556_ _1191_ _1207_ _1208_ _1193_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2325_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[9\] _1734_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[10\]
+ VGND VGND VPWR VPWR _1738_ sky130_fd_sc_hd__a21oi_1
X_2256_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] _1556_ _1568_ net121
+ VGND VGND VPWR VPWR _1678_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2187_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] VGND VGND VPWR VPWR
+ _1609_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_84_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout132_X net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1943__S net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3350__B2 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2014__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input62_X net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1853__S net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2110_ net254 net59 net83 VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__mux2_1
Xhold2 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[15\] VGND VGND VPWR VPWR net206
+ sky130_fd_sc_hd__dlygate4sd3_1
X_3090_ _0840_ _0907_ _0923_ _0925_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2041_ net248 net64 net87 VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3992_ net187 VGND VGND VPWR VPWR rdata[15] sky130_fd_sc_hd__buf_2
X_2943_ _0513_ _0515_ _0777_ _0778_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2874_ _0556_ _0558_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__nand2_1
XANTENNA__2080__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[46\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1825_ _1591_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[61\] _1508_ VGND
+ VGND VPWR VPWR _1514_ sky130_fd_sc_hd__or3_1
XFILLER_0_32_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2907__B2 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3426_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] _1651_ _1260_ VGND
+ VGND VPWR VPWR _1261_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3357_ _1021_ _1049_ VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__xnor2_1
X_2308_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\] _1723_ VGND VGND VPWR VPWR _1726_
+ sky130_fd_sc_hd__nor2_1
X_3288_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[60\]
+ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__and2_1
X_2239_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[43\] VGND VGND VPWR VPWR
+ _1661_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1938__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1885__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input22_A addr[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3897__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[46\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2009__S net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1848__S net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2062__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2590_ _1600_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[3\] _0371_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\]
+ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__a22o_1
XANTENNA__3364__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3211_ _1045_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3142_ _1610_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[41\] _0975_ _0976_
+ _0977_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__o221ai_1
XANTENNA__1876__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3073_ _0605_ _0801_ _0802_ _0604_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__o31a_1
XFILLER_0_89_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2024_ net280 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] net94 VGND
+ VGND VPWR VPWR _0170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3975_ myPWM.g_pwm_channel\[0\].CHANNEL.pwm_out VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_1
XANTENNA__2053__A1 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2926_ _0495_ _0498_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2857_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[33\]
+ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1808_ _1567_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\] _1496_ VGND
+ VGND VPWR VPWR _1497_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2788_ _0611_ _0618_ _0623_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3409_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] _1241_ VGND VGND VPWR VPWR
+ _1244_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_5_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1867__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3449__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2044__A1 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3184__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1858__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3760_ clknet_leaf_13_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[7\] net161
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[7\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__2035__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2711_ _0540_ _0545_ _0539_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_30_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3691_ clknet_leaf_29_CLK _0051_ net143 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2642_ _1621_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[56\] _0475_ _0476_
+ _0477_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_78_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2573_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\]
+ _0407_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1849__A1 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3125_ _1615_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\] VGND VGND VPWR
+ VPWR _0961_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3056_ _0500_ _0891_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__xnor2_1
X_2007_ net260 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] net97 VGND VGND
+ VPWR VPWR _0153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3938__RESET_B net144 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3958_ clknet_leaf_33_CLK _0250_ net140 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3889_ clknet_leaf_21_CLK _0215_ net163 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[38\]
+ sky130_fd_sc_hd__dfrtp_2
X_2909_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[26\] _0740_ VGND VGND VPWR VPWR
+ _0745_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2112__S net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1951__S net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2265__B2 _1594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2022__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_CLK CLK VGND VGND VPWR VPWR clknet_0_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_47_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2256__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2008__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3812_ clknet_leaf_5_CLK _0138_ net152 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3743_ clknet_leaf_43_CLK _0103_ net133 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[56\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_55_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3674_ clknet_leaf_1_CLK _0034_ net135 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_70_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2625_ _0459_ _0460_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2556_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] _0399_ VGND VGND VPWR VPWR
+ _0401_ sky130_fd_sc_hd__and2_1
X_2487_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[2\] _0352_ net70 VGND VGND VPWR
+ VPWR _0355_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2168__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3108_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] _1642_ VGND VGND VPWR VPWR
+ _0944_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3772__RESET_B net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3039_ _0538_ _0774_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2107__S net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1946__S net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2631__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2988__D myPWM.g_pwm_channel\[0\].CHANNEL.alignment VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout75_X net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2017__S net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1856__S net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_584 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput36 wdata[11] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_2
Xinput25 addr[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xinput14 addr[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
XANTENNA__2410__B2 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput47 wdata[21] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput58 wdata[31] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_2
XFILLER_0_52_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2410_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] _1725_ _1737_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\]
+ _0272_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__a221o_1
X_3390_ _1011_ _1220_ _1016_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_75_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2341_ _1712_ _1748_ _1749_ VGND VGND VPWR VPWR _1750_ sky130_fd_sc_hd__or3_1
X_2272_ _1551_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\] _1557_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[8\]
+ VGND VGND VPWR VPWR _1694_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_48_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1987_ net288 net48 net74 VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_562 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3726_ clknet_leaf_27_CLK _0086_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[39\]
+ sky130_fd_sc_hd__dfrtp_4
X_3657_ clknet_leaf_30_CLK _0017_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_3588_ _1021_ _1407_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2608_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[16\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[16\]
+ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__xor2_1
X_2539_ _0351_ _0388_ _0389_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[19\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__3282__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2468__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2361__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input52_A wdata[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2459__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2890_ net111 _0675_ _0677_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__a21o_1
X_1910_ net265 net38 net80 VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1841_ net8 net11 net10 net14 VGND VGND VPWR VPWR _1529_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_25_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3511_ _1331_ _1333_ _1344_ VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__nand3_1
XFILLER_0_4_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3442_ _1162_ _1163_ _1166_ _1160_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__and4b_1
XFILLER_0_100_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3373_ net125 _1192_ _1194_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\] VGND VGND
+ VPWR VPWR _1208_ sky130_fd_sc_hd__o22ai_1
X_2324_ _1737_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[9\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_20_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2255_ _1562_ net123 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] _1569_
+ _1676_ VGND VGND VPWR VPWR _1677_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2186_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\] VGND VGND VPWR VPWR
+ _1608_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_84_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3709_ clknet_leaf_0_CLK _0069_ net134 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_95_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2120__S net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4000__195 VGND VGND VPWR VPWR _4000__195/HI net195 sky130_fd_sc_hd__conb_1
XFILLER_0_78_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3187__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2377__B1 _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input55_X net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[24\] VGND VGND VPWR VPWR net207
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2040_ net298 net63 net88 VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3991_ net186 VGND VGND VPWR VPWR rdata[14] sky130_fd_sc_hd__buf_2
XFILLER_0_71_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2942_ _1608_ _1648_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2873_ _0684_ _0704_ _0708_ _0703_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__a31o_1
X_1824_ _1501_ _1507_ _1509_ _1512_ VGND VGND VPWR VPWR _1513_ sky130_fd_sc_hd__or4_1
XFILLER_0_60_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3425_ _1141_ _1258_ _1128_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3356_ _1051_ _1054_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__xnor2_1
X_3287_ _1120_ _1121_ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__nor2_1
X_2307_ _1725_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[4\]
+ sky130_fd_sc_hd__inv_2
X_2238_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[44\] VGND VGND VPWR VPWR
+ _1660_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2169_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] VGND VGND VPWR VPWR _1591_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_67_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2115__S net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2672__A_N myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2359__B1 _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1954__S net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input15_A addr[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2025__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1864__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3011__B2 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3210_ _1043_ _1044_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__or2_1
X_3141_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\] _1648_ VGND VGND VPWR VPWR _0977_
+ sky130_fd_sc_hd__nand2_1
X_3072_ _0605_ _0803_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2023_ net324 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] net94 VGND
+ VGND VPWR VPWR _0169_ sky130_fd_sc_hd__mux2_1
X_3992__187 VGND VGND VPWR VPWR _3992__187/HI net187 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_81_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3974_ net171 VGND VGND VPWR VPWR error sky130_fd_sc_hd__buf_2
XFILLER_0_18_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3250__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3250__B2 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2443__B net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2925_ _0463_ _0469_ _0760_ _0464_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_33_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2856_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[33\]
+ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__and2_1
XANTENNA__3797__RESET_B net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1807_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] _1655_ _1656_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[16\]
+ VGND VGND VPWR VPWR _1496_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2787_ _0622_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__inv_2
XANTENNA__3274__B myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3408_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] _1241_ _1242_ net121 VGND VGND
+ VPWR VPWR _1243_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input7_A addr[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3339_ _1069_ _1173_ _1090_ VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_69_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1949__S net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3449__B myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[46\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1859__S net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2710_ _0545_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__inv_2
XANTENNA__3890__RESET_B net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3690_ clknet_leaf_31_CLK _0050_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2641_ _0466_ _0467_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__nand2_1
X_2572_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\] _0409_ VGND VGND VPWR VPWR
+ _0412_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3124_ _0954_ _0957_ _0959_ _0953_ _0958_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_66_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3055_ _0501_ _0870_ _0503_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__o21ai_1
X_2006_ net301 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\] net96 VGND VGND
+ VPWR VPWR _0152_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout152_A net154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3957_ clknet_leaf_30_CLK _0249_ net143 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3907__RESET_B net154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2908_ _0743_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3888_ clknet_leaf_21_CLK _0214_ net163 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[37\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2839_ _0495_ _0674_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3195__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2539__A _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3811_ clknet_leaf_4_CLK _0137_ net150 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3742_ clknet_leaf_0_CLK _0102_ net136 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3673_ clknet_leaf_1_CLK _0033_ net134 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\]
+ sky130_fd_sc_hd__dfrtp_4
X_2624_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[63\]
+ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2555_ _0399_ _0400_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[24\]
+ sky130_fd_sc_hd__nor2_1
X_2486_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[0\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[1\]
+ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[2\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.count_enable
+ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__and4_1
X_3998__193 VGND VGND VPWR VPWR _3998__193/HI net193 sky130_fd_sc_hd__conb_1
X_3107_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] _1642_ VGND VGND VPWR VPWR
+ _0943_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3038_ _0545_ _0873_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__xnor2_1
XANTENNA__2184__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2123__S net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3829__RESET_B net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput37 wdata[12] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_12_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput26 addr[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput15 addr[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput59 wdata[3] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_2
Xinput48 wdata[22] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_2
XANTENNA__2033__S net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1872__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2340_ net123 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[14\]
+ _1742_ VGND VGND VPWR VPWR _1749_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2271_ _1549_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[0\] _1572_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\]
+ _1692_ VGND VGND VPWR VPWR _1693_ sky130_fd_sc_hd__o221a_1
XANTENNA__1921__A1 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3426__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1988__A1 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1986_ net300 net47 net74 VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3725_ clknet_leaf_29_CLK _0085_ net143 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[38\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_55_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3656_ clknet_leaf_33_CLK _0016_ net139 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_3587_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\] _1411_ _1412_ net126 VGND VGND
+ VPWR VPWR _1422_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2607_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[18\]
+ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2538_ net110 net109 _0385_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__and3_1
XANTENNA__1912__A1 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2469_ _1614_ net111 _1618_ net109 _0330_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2118__S net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1979__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1957__S net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_2_0__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_4005__200 VGND VGND VPWR VPWR _4005__200/HI net200 sky130_fd_sc_hd__conb_1
XANTENNA_input45_A wdata[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1903__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout170 net33 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_4
XANTENNA__3408__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_88_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2028__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1867__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1840_ net4 net7 net6 net9 VGND VGND VPWR VPWR _1528_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_25_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3510_ _1331_ _1333_ _1344_ VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2395__A1 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3441_ _1263_ _1275_ _1264_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3372_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\] _1194_ _1195_ net126 _1206_
+ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__a221oi_1
X_2323_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[9\] _1734_ _1736_ VGND VGND VPWR
+ VPWR _1737_ sky130_fd_sc_hd__o21ai_2
X_2254_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] _1577_ _1592_ net117
+ VGND VGND VPWR VPWR _1676_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2185_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\] VGND VGND VPWR VPWR _1607_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1969_ net220 net60 net75 VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3708_ clknet_leaf_0_CLK _0068_ net134 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_95_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3639_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[7\] _1664_ _1472_ _1473_ VGND VGND
+ VPWR VPWR _1474_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2356__B myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_66_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Left_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input48_X net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold4 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[42\] VGND VGND VPWR VPWR net208
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_58_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3990_ net185 VGND VGND VPWR VPWR rdata[13] sky130_fd_sc_hd__buf_2
XFILLER_0_71_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2941_ _0514_ _0776_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2872_ net116 _0683_ _0698_ _0699_ _0700_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1823_ net118 _1651_ _1652_ net119 _1511_ VGND VGND VPWR VPWR _1512_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3424_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] _1653_ _1122_ _1132_
+ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3355_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[8\] _1189_ VGND VGND VPWR VPWR _1190_
+ sky130_fd_sc_hd__nor2_1
X_3286_ _1094_ _1108_ _1114_ _1018_ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__o211a_1
X_2306_ net71 _1723_ _1724_ VGND VGND VPWR VPWR _1725_ sky130_fd_sc_hd__or3_1
X_2237_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[45\] VGND VGND VPWR VPWR
+ _1659_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2168_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] VGND VGND VPWR VPWR
+ _1590_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2099_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.count_enable net34 _1545_ VGND VGND
+ VPWR VPWR _0241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2359__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout95_A _1541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1970__S net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2367__A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2404__A1_N myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2041__S net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1880__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3140_ _0972_ _0973_ _0974_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__a21bo_1
X_3071_ _0851_ _0905_ _0906_ _0835_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__a211o_1
X_2022_ net237 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] net94 VGND
+ VGND VPWR VPWR _0168_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3973_ clknet_leaf_2_CLK _0265_ net138 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2924_ _0472_ _0588_ _0466_ _0470_ _0471_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__a2111o_1
X_2855_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[2\] _0690_ VGND VGND VPWR VPWR _0691_
+ sky130_fd_sc_hd__or2_1
X_1806_ _1490_ _1492_ _1493_ _1491_ VGND VGND VPWR VPWR _1495_ sky130_fd_sc_hd__or4b_1
XFILLER_0_72_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2786_ _0620_ _0621_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_92_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3407_ _1104_ _1239_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__xnor2_1
XANTENNA__3766__RESET_B net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3338_ _1063_ _1089_ _1172_ _1062_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__o31a_1
XANTENNA__2265__A2_N net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3269_ _1102_ _1103_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_69_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2187__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2277__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1965__S net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout98_X net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2268__B1 _1562_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3480__A2 _1312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2036__S net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2640_ _0466_ _0470_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1875__S net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2571_ _0411_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[29\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3123_ _1626_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[58\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[57\]
+ _1624_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3054_ _0888_ _0889_ _0869_ _0872_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_38_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2005_ net275 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] net97 VGND VGND
+ VPWR VPWR _0151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3956_ clknet_2_1__leaf_CLK _0248_ net143 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout145_A net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2907_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[26\] _0740_ _0742_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\]
+ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_91_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3887_ clknet_leaf_21_CLK _0213_ net164 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_36_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_36_CLK sky130_fd_sc_hd__clkbuf_8
X_2838_ _0489_ _0498_ _0672_ _0567_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2769_ _0603_ _0604_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__nand2_4
XANTENNA_fanout100_X net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_27_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2098__Y _1545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3810_ clknet_leaf_5_CLK _0136_ net152 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3741_ clknet_leaf_0_CLK _0101_ net134 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_18_CLK clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_18_CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__2290__A myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3672_ clknet_leaf_1_CLK _0032_ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2623_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[63\]
+ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2554_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[24\] _0396_ net69 VGND VGND VPWR
+ VPWR _0400_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2485_ _0351_ _0352_ _0353_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[1\]
+ sky130_fd_sc_hd__nor3_1
X_3106_ _1619_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\] _0940_ _0941_
+ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__a211o_1
XFILLER_0_77_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3037_ _0538_ _0774_ _0536_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3296__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3939_ clknet_leaf_38_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[16\]
+ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_61_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3380__B2 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3477__Y _1312_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_30_Left_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput16 addr[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_12_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput27 addr[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
Xinput38 wdata[13] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_2
Xinput49 wdata[23] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3371__B2 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2270_ _1552_ net127 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] _1591_
+ VGND VGND VPWR VPWR _1692_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_7_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_7_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_48_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1985_ net270 net46 net74 VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__mux2_1
XANTENNA__2291__Y _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3724_ clknet_leaf_28_CLK _0084_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[37\]
+ sky130_fd_sc_hd__dfrtp_2
X_3655_ clknet_leaf_30_CLK _0015_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2606_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[22\]
+ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__xor2_1
X_3586_ net126 _1412_ _1413_ net127 _1420_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__o221a_1
XFILLER_0_11_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2537_ net110 _0385_ net109 VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__a21oi_1
X_2468_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] _1613_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[24\]
+ _1622_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__a22o_1
X_2399_ _1711_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable VGND VGND VPWR VPWR
+ _0270_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_78_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3962__RESET_B net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1973__S net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout80_X net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input38_A wdata[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout160 net161 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_17_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2044__S net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3229__A_N myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[46\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1883__S net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3440_ _1270_ _1271_ _1272_ _1267_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__a31o_1
XFILLER_0_69_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3371_ net126 _1195_ _1197_ net127 _1205_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__o221a_1
X_2322_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[9\] _1734_ net71 VGND VGND VPWR
+ VPWR _1736_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2253_ _1570_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] _1586_ net118 _1674_
+ VGND VGND VPWR VPWR _1675_ sky130_fd_sc_hd__a221o_1
X_2184_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] VGND VGND VPWR VPWR
+ _1606_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1968_ net225 net59 net75 VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__mux2_1
X_1899_ net224 net56 net79 VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__mux2_1
X_3707_ clknet_leaf_0_CLK _0067_ net135 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_95_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3638_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[7\] _1664_ _1665_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[6\]
+ VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3569_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[8\] _1403_ VGND VGND VPWR VPWR _1404_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1897__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1968__S net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1888__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold5 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[46\] VGND VGND VPWR VPWR net209
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2039__S net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1878__S net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2940_ _0536_ _0543_ _0542_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2871_ net115 _0706_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1822_ _1589_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[60\] _1510_ VGND
+ VGND VPWR VPWR _1511_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3423_ _1120_ _1121_ _1136_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__or3b_1
X_3354_ _1169_ _1188_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__or2_1
X_3285_ _1003_ _1010_ _1014_ _1119_ _1018_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__o41a_1
X_2305_ net126 _1720_ VGND VGND VPWR VPWR _1724_ sky130_fd_sc_hd__nor2_1
X_2236_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[46\] VGND VGND VPWR VPWR
+ _1658_ sky130_fd_sc_hd__inv_2
X_2167_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[28\] VGND VGND VPWR VPWR _1589_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2098_ _1533_ _1539_ VGND VGND VPWR VPWR _1545_ sky130_fd_sc_hd__nor2_2
XANTENNA__2056__A1 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2047__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input60_X net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3070_ net108 _0837_ _0843_ net109 _0838_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_89_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2021_ net262 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] net94 VGND
+ VGND VPWR VPWR _0167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3972_ clknet_leaf_37_CLK _0264_ net145 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2923_ _0645_ _0738_ _0753_ _0758_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_33_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2854_ _0525_ _0531_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1805_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] _1655_ VGND VGND VPWR VPWR
+ _1494_ sky130_fd_sc_hd__nor2_1
XANTENNA__3538__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_2785_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[61\]
+ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3406_ _1098_ _1240_ VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3337_ _1088_ _1171_ _1061_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__o21ba_1
X_3268_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[51\]
+ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_69_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2277__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3199_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[2\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[34\]
+ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__or2_1
X_2219_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[50\] VGND VGND VPWR VPWR
+ _1641_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_77_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3299__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2029__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_86_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1981__S net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input20_A addr[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_95_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2052__S net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2570_ _0409_ _0410_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_78_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1891__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3122_ _1627_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[59\] VGND VGND VPWR
+ VPWR _0958_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3053_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\] _0859_ _0887_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[6\]
+ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2004_ net221 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] net96 VGND VGND
+ VPWR VPWR _0150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3955_ clknet_leaf_26_CLK myPWM.g_pwm_channel\[0\].CHANNEL.pwm_next net148 VGND VGND
+ VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.pwm_out sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2906_ _0609_ _0741_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__xnor2_1
XANTENNA__2751__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout138_A net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3886_ clknet_leaf_22_CLK _0212_ net162 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[35\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2837_ _0489_ _0498_ _0672_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__nand3_1
XFILLER_0_45_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2768_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[25\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[57\]
+ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__nand2_2
X_2699_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[37\]
+ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2198__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1976__S net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3982__177 VGND VGND VPWR VPWR _3982__177/HI net177 sky130_fd_sc_hd__conb_1
XFILLER_0_47_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2047__S net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1886__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3740_ clknet_leaf_0_CLK _0100_ net134 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2413__B2 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2964__A2 _0798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3671_ clknet_leaf_2_CLK _0031_ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[17\]
+ sky130_fd_sc_hd__dfrtp_2
X_2622_ _0440_ _0458_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.rollover_flag_c
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2553_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[24\]
+ _0395_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2484_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[0\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.count_enable
+ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[1\] VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__a21oi_1
X_3105_ net110 _1641_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__nor2_1
X_3036_ _1611_ _0871_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2101__A0 myPWM.g_pwm_channel\[0\].CHANNEL.alignment VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3938_ clknet_leaf_36_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[15\]
+ net144 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[15\] sky130_fd_sc_hd__dfrtp_1
X_3869_ clknet_leaf_8_CLK _0195_ net157 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2199__Y _1621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput28 addr[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput17 addr[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput39 wdata[14] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3397__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_1984_ net287 net44 net74 VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3723_ clknet_leaf_29_CLK _0083_ net143 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[36\]
+ sky130_fd_sc_hd__dfrtp_4
X_3654_ clknet_leaf_29_CLK _0014_ net143 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_2605_ _1623_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[25\] VGND VGND VPWR
+ VPWR _0442_ sky130_fd_sc_hd__xnor2_1
X_3585_ net127 _1413_ _1414_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\] _1419_
+ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2536_ net110 _0385_ _0387_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[18\]
+ sky130_fd_sc_hd__a21oi_1
X_2467_ _0332_ _0333_ _0334_ _0335_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__nand4_1
XFILLER_0_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2322__B1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2398_ _1578_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[23\] VGND VGND VPWR
+ VPWR _0269_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3019_ _0491_ _0854_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__xnor2_1
XANTENNA__2482__Y _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout161 net169 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_4
Xfanout150 net151 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout73_X net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2616__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3988__183 VGND VGND VPWR VPWR _3988__183/HI net183 sky130_fd_sc_hd__conb_1
XFILLER_0_69_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3672__RESET_B net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3370_ net127 _1197_ _1203_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\] _1204_
+ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__a221o_1
XANTENNA__2060__S net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2321_ _1735_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[8\]
+ sky130_fd_sc_hd__inv_2
X_2252_ _1565_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[15\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\]
+ _1567_ VGND VGND VPWR VPWR _1674_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2183_ net116 VGND VGND VPWR VPWR _1605_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3280__A1 _1094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3032__B2 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3706_ clknet_leaf_1_CLK _0066_ net135 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1967_ net256 net56 net75 VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__mux2_1
X_1898_ net213 net45 net79 VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3637_ _1469_ _1470_ _1471_ VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__a21o_1
X_3568_ _1083_ _1306_ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2543__B1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2519_ net113 _0375_ _0350_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3499_ _0998_ _1323_ _1324_ _1325_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__or4_1
XFILLER_0_39_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2653__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1984__S net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input50_A wdata[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_CLK_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold6 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[35\] VGND VGND VPWR VPWR net210
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_58_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2055__S net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2870_ _0556_ _0705_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__nand2_1
X_1821_ _1593_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[62\] VGND VGND VPWR
+ VPWR _1510_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3422_ _1236_ _1244_ _1254_ _1256_ _1253_ VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__a311o_1
XFILLER_0_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3353_ _1053_ _1057_ _1083_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3284_ _1118_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__inv_2
X_2304_ net127 net126 _1717_ VGND VGND VPWR VPWR _1723_ sky130_fd_sc_hd__and3_1
X_2235_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[47\] VGND VGND VPWR VPWR
+ _1657_ sky130_fd_sc_hd__inv_2
X_2166_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] VGND VGND VPWR VPWR
+ _1588_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout168_A net169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2097_ net281 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[63\] net90 VGND
+ VGND VPWR VPWR _0240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2999_ net107 _0833_ _0834_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[22\] VGND VGND
+ VPWR VPWR _0835_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_71_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3821__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1979__S net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input53_X net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2020_ net288 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] net95 VGND
+ VGND VPWR VPWR _0166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1889__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2574__A _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3971_ clknet_leaf_34_CLK _0263_ net132 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2922_ _0645_ _0750_ _0754_ _0755_ _0757_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__a311o_1
XFILLER_0_18_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2853_ _0532_ _0688_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1804_ net121 _1654_ VGND VGND VPWR VPWR _1493_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2784_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[61\]
+ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3405_ _1104_ _1239_ _1110_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__a21o_1
X_3336_ _1079_ _1080_ _1169_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__and3_1
X_3267_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[51\]
+ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_69_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3198_ _1551_ _1669_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__nor2_1
X_2218_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\] VGND VGND VPWR VPWR
+ _1640_ sky130_fd_sc_hd__inv_2
X_2149_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR _1571_
+ sky130_fd_sc_hd__inv_2
XANTENNA__3775__RESET_B net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3704__RESET_B net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1788__A1 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input13_A addr[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3121_ _0951_ _0956_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3456__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3052_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\] _0874_ _0887_ net116 _0886_
+ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__o221a_1
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2003_ net278 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] net96 VGND VGND
+ VPWR VPWR _0149_ sky130_fd_sc_hd__mux2_1
X_3954_ clknet_leaf_40_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[31\]
+ net131 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[31\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_85_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2905_ _0593_ _0605_ _0616_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__a21o_1
X_3885_ clknet_leaf_23_CLK _0211_ net160 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[34\]
+ sky130_fd_sc_hd__dfrtp_2
X_2836_ _0488_ _0670_ _0566_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2767_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[25\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[57\]
+ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2698_ _0519_ _0533_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__nand2_1
XANTENNA_input5_A addr[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3319_ _1153_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_1_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2661__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1992__S net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2110__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_503 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2063__S net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3670_ clknet_leaf_37_CLK _0030_ net144 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_2621_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] _0414_ _0455_ _0457_
+ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2552_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[23\] VGND VGND VPWR VPWR
+ _0398_ sky130_fd_sc_hd__inv_2
XANTENNA__1924__A1 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2483_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[0\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[1\]
+ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.count_enable VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__and3_1
XANTENNA__3126__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3104_ net109 _1640_ _1641_ net110 VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__a22o_1
X_3035_ _0504_ _0870_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__xor2_2
XANTENNA__2101__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2762__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3937_ clknet_leaf_36_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[14\]
+ net144 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[14\] sky130_fd_sc_hd__dfrtp_1
X_3868_ clknet_leaf_8_CLK _0194_ net157 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3799_ clknet_leaf_15_CLK _0125_ net165 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3593__A _1560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2819_ _0473_ _0654_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1915__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1987__S net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput18 addr[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
Xinput29 addr[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_75_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1906__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2058__S net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1897__S net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1983_ net226 net43 net74 VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3722_ clknet_leaf_31_CLK _0082_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[35\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3653_ clknet_leaf_41_CLK _0013_ net130 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_2604_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[28\]
+ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3584_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\] _1414_ _1416_ _1417_ _1418_
+ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__o221a_1
XFILLER_0_11_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2535_ net110 _0385_ net69 VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__o21ai_1
X_2466_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[3\] _1601_ _1606_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\]
+ _0327_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__o221a_1
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2397_ _1592_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[30\] VGND VGND VPWR
+ VPWR _0268_ sky130_fd_sc_hd__or2_1
X_3018_ _0487_ _0785_ _0486_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1833__B1 myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3824__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3971__RESET_B net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout140 net141 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
Xfanout151 net154 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_4
Xfanout162 net164 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_17_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3734__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2320_ net72 _1733_ _1734_ VGND VGND VPWR VPWR _1735_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2251_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] _1550_ _1555_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[7\]
+ _1672_ VGND VGND VPWR VPWR _1673_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2182_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\] VGND VGND VPWR VPWR
+ _1604_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1966_ net235 net45 net76 VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3705_ clknet_leaf_1_CLK _0065_ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1897_ net231 net34 net79 VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3636_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[6\] _1665_ _1666_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\]
+ VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3567_ _1560_ _1400_ VGND VGND VPWR VPWR _1402_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2518_ _0375_ _0376_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[11\]
+ sky130_fd_sc_hd__nor2_1
X_3498_ net117 _1330_ _1332_ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__o21a_1
X_2449_ _0314_ _0315_ _0316_ _0317_ _0309_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3819__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input43_A wdata[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2397__A _1592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold7 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[50\] VGND VGND VPWR VPWR net211
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2470__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1820_ _1591_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[61\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[60\]
+ _1589_ _1508_ VGND VGND VPWR VPWR _1509_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2071__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3893__RESET_B net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3421_ _1223_ _1227_ _1235_ _1255_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__o211ai_1
X_3352_ _1080_ _1186_ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2303_ _1722_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[3\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_0_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3283_ _1116_ _1117_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__nand2_2
X_2234_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\] VGND VGND VPWR VPWR
+ _1656_ sky130_fd_sc_hd__inv_2
X_2165_ net118 VGND VGND VPWR VPWR _1587_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2096_ net292 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[62\] net90 VGND
+ VGND VPWR VPWR _0239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2770__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2998_ _0470_ _0829_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1949_ net302 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\] net99 VGND
+ VGND VPWR VPWR _0098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3619_ _1360_ _1361_ _1450_ _1354_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__or4b_1
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2680__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1995__S net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input46_X net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2066__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3970_ clknet_leaf_34_CLK _0262_ net139 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2921_ _1632_ _0632_ _0756_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\] VGND VGND
+ VPWR VPWR _0757_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_17_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2852_ _0519_ _0520_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__nand2_2
X_1803_ _1571_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[51\] VGND VGND VPWR
+ VPWR _1492_ sky130_fd_sc_hd__and2_1
X_2783_ _0611_ _0618_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3404_ _1106_ _1238_ _1112_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__a21o_1
X_3335_ _1080_ _1169_ _1086_ VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__a21o_1
X_3266_ _1099_ _1100_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2217_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\] VGND VGND VPWR VPWR
+ _1639_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3197_ _1031_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2148_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] VGND VGND VPWR VPWR
+ _1570_ sky130_fd_sc_hd__inv_2
X_2079_ net274 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[45\] net93 VGND
+ VGND VPWR VPWR _0222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_39_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_39_CLK sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_18_CLK_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3744__RESET_B net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout93_A _1544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3832__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2962__X _0798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3120_ _0950_ _0952_ _0955_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__a21o_1
XFILLER_0_93_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3051_ _0516_ _0780_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__xor2_1
X_2002_ net220 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] net96 VGND VGND
+ VPWR VPWR _0148_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3953_ clknet_leaf_40_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[30\]
+ net131 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3884_ clknet_leaf_21_CLK _0210_ net162 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[33\]
+ sky130_fd_sc_hd__dfrtp_2
X_2904_ _0601_ _0739_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3917__Q myPWM.g_pwm_channel\[0\].CHANNEL.alignment VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2835_ _0488_ _0670_ _0565_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_73_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2766_ _0597_ _0600_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2697_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] _1649_ _0525_ _0531_
+ _0521_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3318_ _1151_ _1152_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__nand2_2
X_3249_ _1083_ _1080_ _1079_ _1071_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__and4b_1
XANTENNA__2495__A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3827__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout96_X net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3666__RESET_B net144 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2620_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] _0411_ _0416_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\]
+ _0456_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2551_ _0396_ _0397_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[23\]
+ sky130_fd_sc_hd__nor2_1
X_2482_ net69 VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_50_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3103_ _0938_ _0934_ _0933_ _0931_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__and4bb_1
X_3034_ _0782_ _0783_ _0765_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1860__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout143_A net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3936_ clknet_leaf_35_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[13\]
+ net141 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3867_ clknet_leaf_8_CLK _0193_ net157 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3798_ clknet_leaf_15_CLK _0124_ net165 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_2818_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] _1638_ _0646_ VGND
+ VGND VPWR VPWR _0654_ sky130_fd_sc_hd__a21oi_1
X_2749_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] _1639_ _0584_ VGND
+ VGND VPWR VPWR _0585_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1851__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput19 addr[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_467 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2074__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1982_ net271 net42 net74 VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3721_ clknet_leaf_33_CLK _0081_ net140 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[34\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_28_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3652_ clknet_leaf_41_CLK _0012_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3583_ _1416_ _1417_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[1\] VGND VGND VPWR
+ VPWR _1418_ sky130_fd_sc_hd__a21o_1
X_2603_ _1628_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[29\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[31\]
+ _1631_ _0439_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2534_ _0385_ _0386_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[17\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2465_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\] _1597_ _1623_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\]
+ _0313_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__o221a_1
X_2396_ net117 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] _1784_ _0267_ net72
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[31\] sky130_fd_sc_hd__a311oi_2
XFILLER_0_78_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3017_ _0498_ _0852_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3586__B2 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3919_ clknet_leaf_21_CLK _0245_ net163 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout130 net131 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_4
XANTENNA__3840__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout152 net154 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_4
Xfanout163 net164 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__buf_2
Xfanout141 net149 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1998__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2001__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2250_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] _1550_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\]
+ _1560_ VGND VGND VPWR VPWR _1672_ sky130_fd_sc_hd__o22ai_1
XANTENNA__2069__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2181_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[4\] VGND VGND VPWR VPWR _1603_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1965_ net245 net34 net75 VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3704_ clknet_leaf_2_CLK _0064_ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1896_ _1548_ net338 net77 VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3635_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\] _1666_ _1667_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[4\]
+ VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__o22a_1
XFILLER_0_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3566_ _1078_ _1399_ VGND VGND VPWR VPWR _1401_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2768__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2517_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[11\] _0374_ _0350_ VGND VGND VPWR
+ VPWR _0376_ sky130_fd_sc_hd__o21ai_1
X_3497_ _1151_ _1328_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] VGND VGND VPWR
+ VPWR _1332_ sky130_fd_sc_hd__a21o_1
X_2448_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] net108 VGND VGND VPWR
+ VPWR _0317_ sky130_fd_sc_hd__or2_1
XANTENNA__3769__RESET_B net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2379_ net120 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[26\] _1772_ VGND VGND VPWR
+ VPWR _1776_ sky130_fd_sc_hd__and3_1
XANTENNA__2059__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2678__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input36_A wdata[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold8 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[36\] VGND VGND VPWR VPWR net212
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2416__A1_N myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3420_ _1227_ _1231_ _1232_ _1224_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__or4b_1
X_3351_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] _1663_ _1169_ VGND
+ VGND VPWR VPWR _1186_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2302_ net71 _1720_ _1721_ VGND VGND VPWR VPWR _1722_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3862__RESET_B net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3282_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[53\]
+ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__or2_1
X_2233_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[49\] VGND VGND VPWR VPWR
+ _1655_ sky130_fd_sc_hd__inv_2
X_2164_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] VGND VGND VPWR VPWR
+ _1586_ sky130_fd_sc_hd__inv_2
X_2095_ net331 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[61\] net90 VGND
+ VGND VPWR VPWR _0238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2997_ _0473_ _0832_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__xnor2_1
X_1948_ net211 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[50\] net99 VGND
+ VGND VPWR VPWR _0097_ sky130_fd_sc_hd__mux2_1
XANTENNA__3655__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1879_ net251 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[17\] net103 VGND
+ VGND VPWR VPWR _0031_ sky130_fd_sc_hd__mux2_1
X_3618_ _1370_ _1448_ _1451_ _1452_ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__o31a_1
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3549_ _1099_ _1381_ _1105_ VGND VGND VPWR VPWR _1384_ sky130_fd_sc_hd__a21o_1
X_3978__173 VGND VGND VPWR VPWR _3978__173/HI net173 sky130_fd_sc_hd__conb_1
XFILLER_0_98_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2201__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input39_X net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkload1_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2920_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[31\] _0628_ _0631_ _0629_ VGND VGND
+ VPWR VPWR _0756_ sky130_fd_sc_hd__o31a_1
XANTENNA__2871__A net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2082__S net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2851_ _0534_ _0538_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__xnor2_1
X_1802_ _1571_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[51\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[50\]
+ _1569_ VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__o22a_1
X_2782_ _0602_ _0617_ _0614_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3403_ _1094_ _1101_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3334_ _1053_ _1057_ _1083_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_0_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3265_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[17\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[49\]
+ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_37_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2216_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[53\] VGND VGND VPWR VPWR
+ _1638_ sky130_fd_sc_hd__inv_2
X_3196_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[35\]
+ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__xor2_2
X_2147_ net121 VGND VGND VPWR VPWR _1569_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2078_ net303 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[44\] net93 VGND
+ VGND VPWR VPWR _0221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout86_A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Left_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2370__B1 _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2425__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3050_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\] _0874_ _0884_ _0885_ _0876_
+ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__a221o_1
X_2001_ net225 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] net96 VGND VGND
+ VPWR VPWR _0147_ sky130_fd_sc_hd__mux2_1
XANTENNA__2077__S net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2416__B2 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3952_ clknet_leaf_40_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[29\]
+ net130 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2903_ _0593_ _0605_ _0609_ _0617_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__a31o_1
X_3883_ clknet_leaf_23_CLK _0209_ net160 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2834_ _0506_ _0509_ _0556_ _0563_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__o31ai_2
X_2765_ _0600_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_91_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2696_ _0525_ _0531_ _0521_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3317_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[63\]
+ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__or2_1
X_3248_ _1081_ _1082_ VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__and2_2
XANTENNA__2104__A0 myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_3179_ _1012_ _1013_ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_1_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3843__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1861__Y _1535_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2550_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] _0395_ net70 VGND VGND VPWR
+ VPWR _0397_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2481_ _1633_ _0349_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3126__A2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_CLK_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3102_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\] _1635_ VGND VGND VPWR VPWR
+ _0938_ sky130_fd_sc_hd__nor2_1
X_3033_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\] _0859_ _0863_ _0866_ _0868_
+ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_73_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3935_ clknet_leaf_35_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[12\]
+ net144 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3866_ clknet_leaf_12_CLK _0192_ net159 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_3797_ clknet_leaf_16_CLK _0123_ net168 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2817_ _0646_ _0652_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__or2_1
X_2748_ _0481_ _0583_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__and2_1
XANTENNA__3663__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2679_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[39\]
+ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__or2_1
XANTENNA__2876__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4003__198 VGND VGND VPWR VPWR _4003__198/HI net198 sky130_fd_sc_hd__conb_1
XFILLER_0_68_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3838__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input66_A wen VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1981_ net284 net41 net74 VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__mux2_1
X_3720_ clknet_leaf_30_CLK _0080_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[33\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_99_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3651_ clknet_leaf_42_CLK _0011_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2090__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3582_ _1035_ _1295_ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2602_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[27\]
+ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_97_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2533_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] _0384_ net69 VGND VGND VPWR
+ VPWR _0386_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2464_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] _1607_ _1612_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[13\]
+ _0328_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__o221a_1
XFILLER_0_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2395_ net117 _1784_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] VGND VGND VPWR
+ VPWR _0267_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3215__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3016_ _0487_ _0492_ _0785_ _0790_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__a31o_1
XFILLER_0_66_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1833__A2 _1521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3658__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3918_ clknet_leaf_2_CLK _0244_ net153 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_mod\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3849_ clknet_leaf_2_CLK _0175_ net153 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_89_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout120 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[25\] VGND VGND VPWR VPWR net120
+ sky130_fd_sc_hd__buf_2
Xfanout131 net132 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_4
Xfanout153 net154 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_4
Xfanout164 net169 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_4
Xfanout142 net143 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2180_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] VGND VGND VPWR VPWR
+ _1602_ sky130_fd_sc_hd__inv_2
XANTENNA__2296__D myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2085__S net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1964_ _1536_ _1539_ VGND VGND VPWR VPWR _1540_ sky130_fd_sc_hd__nor2_4
XFILLER_0_50_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3703_ clknet_leaf_2_CLK _0063_ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[48\]
+ sky130_fd_sc_hd__dfrtp_1
X_3634_ net126 _1667_ _1668_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[3\] _1468_
+ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1895_ _1536_ net26 net66 VGND VGND VPWR VPWR _1537_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_24_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3565_ _1078_ _1399_ VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3496_ net117 _1330_ _1329_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__a21oi_1
X_2516_ net114 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[11\]
+ _0370_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__and4_1
X_2447_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] net108 VGND VGND VPWR
+ VPWR _0316_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2378_ _1774_ _1775_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[25\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__2784__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1990__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout71_X net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold9 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[33\] VGND VGND VPWR VPWR net213
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input29_A addr[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2470__A2 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1981__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3350_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[10\] _1182_ _1184_ net124 VGND VGND
+ VPWR VPWR _1185_ sky130_fd_sc_hd__a22oi_1
X_2301_ net127 _1717_ VGND VGND VPWR VPWR _1721_ sky130_fd_sc_hd__nor2_1
X_3281_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[53\]
+ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__nand2_1
X_2232_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[50\] VGND VGND VPWR VPWR
+ _1654_ sky130_fd_sc_hd__inv_2
X_2163_ net119 VGND VGND VPWR VPWR _1585_ sky130_fd_sc_hd__inv_2
X_2094_ net306 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[60\] net90 VGND
+ VGND VPWR VPWR _0237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2996_ _0588_ _0828_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1947_ net267 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[49\] net99 VGND
+ VGND VPWR VPWR _0096_ sky130_fd_sc_hd__mux2_1
XANTENNA__1972__A1 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1878_ net229 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[16\] net105 VGND
+ VGND VPWR VPWR _0030_ sky130_fd_sc_hd__mux2_1
X_3617_ _1370_ _1449_ _1451_ _1376_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_101_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3548_ _1099_ _1105_ _1381_ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__nand3_1
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3479_ _1101_ _1105_ VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__nand2_1
XANTENNA__3403__A _1094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3468__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2850_ _0545_ _0685_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1801_ _1488_ _1489_ VGND VGND VPWR VPWR _1490_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2781_ _0609_ _0616_ _0615_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3402_ net122 _1175_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3333_ _1162_ _1163_ _1167_ _1160_ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__and4b_1
XFILLER_0_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3264_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[17\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[49\]
+ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2215_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\] VGND VGND VPWR VPWR
+ _1637_ sky130_fd_sc_hd__inv_2
X_3195_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[35\]
+ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2146_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] VGND VGND VPWR VPWR
+ _1568_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout166_A net169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2077_ net259 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[43\] net93 VGND
+ VGND VPWR VPWR _0220_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2979_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\] _0813_ VGND VGND VPWR VPWR
+ _0815_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_32_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1945__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2302__A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout79_A _1537_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2122__A1 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input51_X net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2113__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2000_ net256 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[2\] net96 VGND VGND
+ VPWR VPWR _0146_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3951_ clknet_leaf_40_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[28\]
+ net130 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_58_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2093__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2902_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] _0649_ _0734_ _0737_ VGND VGND
+ VPWR VPWR _0738_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3882_ clknet_leaf_3_CLK _0208_ net151 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2833_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] _0662_ _0668_ net109 VGND VGND
+ VPWR VPWR _0669_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2764_ _0598_ _0599_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__nor2_1
XANTENNA__1927__A1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2695_ _0528_ _0529_ _0530_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3316_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[63\]
+ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__nand2_1
XANTENNA__2776__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3247_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[41\]
+ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__or2_1
XANTENNA__2104__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3178_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[56\]
+ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2129_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[2\] VGND VGND VPWR VPWR
+ _1551_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_37_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout169_X net169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1900__S net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4008__203 VGND VGND VPWR VPWR _4008__203/HI net203 sky130_fd_sc_hd__conb_1
XANTENNA__1918__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3934__RESET_B net144 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input11_A addr[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1909__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2480_ _0336_ _0341_ _0348_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__or3_1
X_3101_ _0930_ _0932_ _0936_ myPWM.g_pwm_channel\[0\].CHANNEL.alignment VGND VGND
+ VPWR VPWR _0937_ sky130_fd_sc_hd__a211o_1
XANTENNA__2088__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3032_ net114 _0860_ _0861_ _0864_ net115 VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__o32a_1
XFILLER_0_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3934_ clknet_leaf_35_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[11\]
+ net144 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2270__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3865_ clknet_leaf_24_CLK _0191_ net159 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_2816_ _0586_ _0589_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__and2_1
X_3796_ clknet_leaf_18_CLK _0122_ net167 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout129_A net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2747_ _0484_ _0582_ _0580_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2678_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[39\]
+ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input3_A addr[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input59_A wdata[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1980_ net332 net40 net73 VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__mux2_1
XANTENNA__2252__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3650_ clknet_leaf_42_CLK _0010_ net128 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_3581_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[32\] _1199_ _1200_ _1415_
+ VGND VGND VPWR VPWR _1416_ sky130_fd_sc_hd__a22o_1
X_2601_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[14\]
+ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_97_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2532_ net111 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[16\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\]
+ _0380_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__and4_1
XFILLER_0_51_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2463_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] _1603_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\]
+ _1629_ _0326_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__o221a_1
X_2394_ net117 _1784_ _0266_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[30\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3015_ _0847_ _0849_ _0850_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_64_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3917_ clknet_leaf_30_CLK _0243_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.alignment
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3848_ clknet_leaf_3_CLK _0174_ net151 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_3779_ clknet_leaf_11_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[26\]
+ net154 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout121 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[18\] VGND VGND VPWR VPWR net121
+ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_20_CLK clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_20_CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__2310__A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout110 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] VGND VGND VPWR VPWR net110
+ sky130_fd_sc_hd__buf_2
Xfanout165 net169 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__buf_4
Xfanout154 net170 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_4
Xfanout132 net33 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__buf_2
Xfanout143 net149 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_4
XANTENNA__3125__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3849__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_2_0__f_CLK_A clknet_0_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_CLK_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3316__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_11_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_11_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_87_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2473__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1963_ net26 net66 VGND VGND VPWR VPWR _1539_ sky130_fd_sc_hd__nand2_1
X_3702_ clknet_leaf_40_CLK _0062_ net130 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1894_ net12 _1532_ net1 net23 VGND VGND VPWR VPWR _1536_ sky130_fd_sc_hd__or4b_4
XFILLER_0_55_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3633_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[3\] _1668_ _1669_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\]
+ _1467_ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__o221a_1
XFILLER_0_70_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3564_ _1306_ _1307_ _1291_ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_11_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2515_ _0351_ _0373_ _0374_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[10\]
+ sky130_fd_sc_hd__nor3_1
X_3495_ _1153_ _1327_ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__xnor2_1
XANTENNA__2130__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2446_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] net110 VGND VGND VPWR
+ VPWR _0315_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2377_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[25\] _1772_ _1713_ VGND VGND VPWR
+ VPWR _1775_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3778__RESET_B net154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_65_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3280_ _1094_ _1108_ _1114_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__o21ai_2
X_2300_ net127 _1717_ VGND VGND VPWR VPWR _1720_ sky130_fd_sc_hd__and2_1
X_2231_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[57\] VGND VGND VPWR VPWR
+ _1653_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2162_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] VGND VGND VPWR VPWR
+ _1584_ sky130_fd_sc_hd__inv_2
X_2093_ net282 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[59\] net90 VGND
+ VGND VPWR VPWR _0236_ sky130_fd_sc_hd__mux2_1
XANTENNA__2096__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2995_ _0466_ _0830_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1946_ net330 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[48\] net99 VGND
+ VGND VPWR VPWR _0095_ sky130_fd_sc_hd__mux2_1
X_1877_ net206 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[15\] net102 VGND
+ VGND VPWR VPWR _0029_ sky130_fd_sc_hd__mux2_1
X_3616_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\] _1368_ _1373_ VGND VGND VPWR
+ VPWR _1451_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3547_ _1101_ _1313_ VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3478_ _1287_ _1312_ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2429_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] _1750_ _1753_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\]
+ _0298_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__a221o_1
XANTENNA__1903__S net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input41_A wdata[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1800_ _1573_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\] _1487_ VGND
+ VGND VPWR VPWR _1489_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2780_ _1623_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[57\] VGND VGND VPWR
+ VPWR _0616_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_1__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_2_1__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3401_ _1227_ _1234_ _1235_ _1224_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__and4b_1
XANTENNA__3772__Q myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_3332_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[28\] _1165_ _1166_ VGND VGND VPWR
+ VPWR _1167_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3263_ _1095_ _1097_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__nand2_2
X_3194_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] _1668_ VGND VGND VPWR
+ VPWR _1029_ sky130_fd_sc_hd__and2_1
X_2214_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\] VGND VGND VPWR VPWR
+ _1636_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2145_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[16\] VGND VGND VPWR VPWR _1567_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_56_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2076_ net261 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[42\] net93 VGND
+ VGND VPWR VPWR _0219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1890__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2978_ _0460_ _0811_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[31\] VGND VGND VPWR
+ VPWR _0814_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_32_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1929_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.rollover_flag myPWM.g_pwm_channel\[0\].CHANNEL.data_mod\[1\]
+ VGND VGND VPWR VPWR _1538_ sky130_fd_sc_hd__nand2_2
XFILLER_0_31_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3682__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1881__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input44_X net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold90 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[47\] VGND VGND VPWR VPWR net294
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_89_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1872__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3950_ clknet_leaf_39_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[27\]
+ net132 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2901_ _0666_ _0669_ _0730_ _0731_ _0736_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__o311a_1
XFILLER_0_58_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3881_ clknet_leaf_3_CLK _0207_ net151 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2832_ _0481_ _0667_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2763_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[59\]
+ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2403__A _1570_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2694_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[34\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\]
+ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3315_ _1145_ _1146_ _0995_ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3246_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[41\]
+ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3177_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[56\]
+ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2128_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[1\] VGND VGND VPWR VPWR _1550_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_65_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1863__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2059_ net286 net52 net85 VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3677__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3409__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__2040__A1 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout91_A _1544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3903__RESET_B net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1854__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3100_ _0931_ _0933_ _0934_ _0935_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__and4_1
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2476__A1_N myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3031_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[9\] _0860_ _0861_ VGND VGND VPWR
+ VPWR _0867_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_62_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3933_ clknet_leaf_35_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[10\]
+ net144 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3864_ clknet_leaf_15_CLK _0190_ net166 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2815_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[22\] _0650_ VGND VGND VPWR VPWR
+ _0651_ sky130_fd_sc_hd__nand2_1
X_3795_ clknet_leaf_18_CLK _0121_ net167 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2133__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2022__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2746_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[17\] _1642_ _0574_ _0581_
+ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__a31o_1
X_2677_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[40\]
+ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__xor2_2
XFILLER_0_68_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3229_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[46\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\]
+ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__nand2b_1
XANTENNA__1911__S net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout94_X net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3580_ _1549_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[32\] VGND VGND VPWR
+ VPWR _1415_ sky130_fd_sc_hd__nand2_1
XANTENNA__2004__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2600_ _0423_ _0424_ _0432_ _0436_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_97_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2531_ _0351_ _0383_ _0384_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[16\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_51_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1792__A _1560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3504__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__2099__S _1545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2462_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[21\] _1620_ _1615_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[15\]
+ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__a2bb2o_1
X_2393_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[30\] _1784_ net72 VGND VGND VPWR
+ VPWR _0266_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3014_ net109 _0843_ _0844_ net110 VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3916_ clknet_leaf_29_CLK _0242_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.polarity
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout141_A net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_88_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3847_ clknet_leaf_4_CLK _0173_ net150 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\]
+ sky130_fd_sc_hd__dfrtp_4
X_3778_ clknet_leaf_11_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[25\]
+ net154 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2729_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[13\] _1644_ VGND VGND VPWR
+ VPWR _0565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1906__S net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout122 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[15\] VGND VGND VPWR VPWR net122
+ sky130_fd_sc_hd__clkbuf_2
Xfanout100 _1538_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__buf_4
Xfanout111 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[15\] VGND VGND VPWR VPWR net111
+ sky130_fd_sc_hd__buf_2
Xfanout155 net156 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_4
Xfanout133 net136 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_4
Xfanout144 net149 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_4
Xfanout166 net169 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1962_ _1548_ net335 net81 VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1893_ net241 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\] net102 VGND
+ VGND VPWR VPWR _0045_ sky130_fd_sc_hd__mux2_1
X_3701_ clknet_leaf_34_CLK _0061_ net139 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_3632_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\] _1669_ _1670_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[1\]
+ _1466_ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3563_ _1559_ _1395_ _1397_ VGND VGND VPWR VPWR _1398_ sky130_fd_sc_hd__nand3_1
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2514_ net114 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\] _0370_ VGND VGND VPWR
+ VPWR _0374_ sky130_fd_sc_hd__and3_1
X_3494_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] _1151_ _1328_ VGND VGND VPWR
+ VPWR _1329_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2445_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] net110 VGND VGND VPWR
+ VPWR _0314_ sky130_fd_sc_hd__or2_1
X_2376_ net120 _1772_ VGND VGND VPWR VPWR _1774_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2464__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout144_X net144 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3101__C1 myPWM.g_pwm_channel\[0\].CHANNEL.alignment VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3327__A _1594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2391__B1 _1713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2230_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[58\] VGND VGND VPWR VPWR
+ _1652_ sky130_fd_sc_hd__inv_2
X_2161_ net120 VGND VGND VPWR VPWR _1583_ sky130_fd_sc_hd__inv_2
X_2092_ net286 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[58\] net90 VGND
+ VGND VPWR VPWR _0235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2994_ _0470_ _0829_ _0469_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__o21a_1
X_1945_ net250 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\] net98 VGND
+ VGND VPWR VPWR _0094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1876_ net246 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] net104 VGND
+ VGND VPWR VPWR _0028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3237__A _1562_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3615_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[24\] _1357_ VGND VGND VPWR VPWR
+ _1450_ sky130_fd_sc_hd__nor2_1
X_3546_ _1101_ _1313_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout104_A _1535_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3477_ _1306_ _1310_ _1311_ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__a21oi_2
X_2428_ _1562_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[12\] VGND VGND VPWR
+ VPWR _0298_ sky130_fd_sc_hd__xnor2_1
X_2359_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] _1760_ _1713_ VGND VGND VPWR
+ VPWR _1762_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_15_CLK_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input34_A wdata[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_476 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3400_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\] _1226_ VGND VGND VPWR VPWR
+ _1235_ sky130_fd_sc_hd__nand2_1
XANTENNA__3156__A2 _0991_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3331_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] _1147_ _1148_ _1165_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[28\]
+ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__a32o_1
X_3262_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\]
+ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__or2_1
X_3193_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[36\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\]
+ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__nand2b_1
X_2213_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[60\] VGND VGND VPWR VPWR
+ _1635_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2144_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] VGND VGND VPWR VPWR
+ _1566_ sky130_fd_sc_hd__inv_2
X_2075_ net243 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[41\] net93 VGND
+ VGND VPWR VPWR _0218_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_2_2__f_CLK_X clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2977_ _0462_ _0810_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_32_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1928_ net230 net58 net77 VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_15_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1859_ net264 net57 net81 VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2355__B1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_3529_ _1355_ _1362_ _1352_ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__o21ba_1
XANTENNA__1914__S net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3762__RESET_B net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Left_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input37_X net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_42_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold80 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[16\] VGND VGND VPWR VPWR net284
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[61\] VGND VGND VPWR VPWR net295
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_89_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2900_ _0651_ _0656_ _0732_ _0735_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__and4_1
XFILLER_0_73_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3880_ clknet_leaf_4_CLK _0206_ net150 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2831_ _0484_ _0661_ _0580_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_51_Left_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2762_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[59\]
+ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2693_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[33\]
+ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__nand2b_1
X_3314_ _0995_ _1145_ _1146_ VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_60_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3245_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[42\]
+ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_67_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3176_ _1007_ _1009_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__or2_2
XFILLER_0_83_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2127_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[0\] VGND VGND VPWR VPWR _1549_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2058_ net322 net51 net85 VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1909__S net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout84_A _1534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3943__RESET_B net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1790__A1 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3030_ net115 _0864_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_62_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3684__RESET_B net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3932_ clknet_leaf_35_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[9\] net141
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[9\] sky130_fd_sc_hd__dfrtp_1
X_3863_ clknet_leaf_15_CLK _0189_ net166 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2270__A2 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2814_ _0470_ _0647_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_42_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3229__B myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3794_ clknet_leaf_20_CLK _0120_ net164 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2745_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] _1641_ VGND VGND VPWR
+ VPWR _0581_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2676_ _1608_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[40\] _0511_ VGND
+ VGND VPWR VPWR _0512_ sky130_fd_sc_hd__o21a_1
XANTENNA__3245__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3228_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] _1658_ VGND VGND VPWR
+ VPWR _1063_ sky130_fd_sc_hd__and2_1
XANTENNA__3286__A1 _1094_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3159_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[62\]
+ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout87_X net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3277__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2530_ net111 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[16\] _0380_ VGND VGND VPWR
+ VPWR _0384_ sky130_fd_sc_hd__and3_1
XANTENNA__1792__B net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2461_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[22\]
+ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__xor2_1
XFILLER_0_51_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2392_ _1784_ _1785_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[29\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3013_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] _0846_ _0848_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[16\]
+ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__a22oi_1
XANTENNA__2409__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3915_ clknet_leaf_29_CLK _0241_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.count_enable
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__2144__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3846_ clknet_leaf_4_CLK _0172_ net150 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3777_ clknet_leaf_11_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[24\]
+ net153 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[24\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2728_ _0499_ _0562_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__and2b_1
XFILLER_0_100_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2659_ _0493_ _0494_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout112 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[13\] VGND VGND VPWR VPWR net112
+ sky130_fd_sc_hd__buf_2
Xfanout101 _1538_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_2
Xfanout156 net170 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_4
Xfanout123 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[12\] VGND VGND VPWR VPWR net123
+ sky130_fd_sc_hd__buf_2
XANTENNA__1922__S net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout134 net136 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_4
Xfanout145 net149 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_2
Xfanout167 net168 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_7_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1993__A1 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input64_A wdata[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3498__A1 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2413__A1_N myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1961_ net230 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[63\] net98 VGND
+ VGND VPWR VPWR _0110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3700_ clknet_leaf_24_CLK _0060_ net144 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1892_ net264 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] net102 VGND
+ VGND VPWR VPWR _0044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1984__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3631_ _1549_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[32\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[1\]
+ _1670_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_24_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3562_ _1083_ _1306_ _1396_ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2513_ net114 _0370_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\] VGND VGND VPWR
+ VPWR _0373_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3493_ _0994_ _0996_ _1326_ _1153_ _0993_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__a311o_1
X_2444_ _1596_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[1\] _1609_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[9\]
+ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__o22a_1
X_2375_ _1773_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[24\]
+ sky130_fd_sc_hd__inv_2
XFILLER_0_75_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2274__A2_N myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout137_X net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3829_ clknet_leaf_16_CLK _0155_ net168 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__1975__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2602__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1917__S net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3716__RESET_B net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1966__A1 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2391__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2160_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] VGND VGND VPWR VPWR
+ _1582_ sky130_fd_sc_hd__inv_2
X_2091_ net322 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[57\] net90 VGND
+ VGND VPWR VPWR _0234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2993_ _0472_ _0588_ _0828_ _0471_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1944_ net209 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\] net100 VGND
+ VGND VPWR VPWR _0093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3614_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\] _1368_ VGND VGND VPWR VPWR
+ _1449_ sky130_fd_sc_hd__or2_1
X_1875_ net227 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[13\] net105 VGND
+ VGND VPWR VPWR _0027_ sky130_fd_sc_hd__mux2_1
X_3545_ _1104_ _1377_ VGND VGND VPWR VPWR _1380_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3476_ _1289_ _1293_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2427_ _1588_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[28\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[30\]
+ _1592_ _0296_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2358_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] _1760_ VGND VGND VPWR VPWR
+ _1761_ sky130_fd_sc_hd__and2_1
X_2289_ _1691_ _1710_ VGND VGND VPWR VPWR _1711_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_27_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input27_A addr[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2507__A net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3330_ _1144_ _1164_ VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__or2_1
X_3261_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\]
+ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__nor2_1
XANTENNA__2116__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3192_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[36\]
+ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__nand2b_2
X_2212_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[62\] VGND VGND VPWR VPWR
+ _1634_ sky130_fd_sc_hd__inv_2
X_2143_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\] VGND VGND VPWR VPWR
+ _1565_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2074_ net248 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[40\] net92 VGND
+ VGND VPWR VPWR _0217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2976_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[31\] _0460_ _0811_ VGND VGND VPWR
+ VPWR _0812_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1927_ net272 net57 net77 VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__mux2_1
XANTENNA__2152__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_1858_ net319 net55 net81 VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1789_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[10\] _1662_ _1476_ _1477_ VGND VGND
+ VPWR VPWR _1478_ sky130_fd_sc_hd__o211a_1
X_3528_ net119 _1353_ VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__xnor2_1
X_3459_ _1553_ _1667_ VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__nor2_1
XANTENNA__2107__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1930__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2327__A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2001__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold70 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[45\] VGND VGND VPWR VPWR net274
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[36\] VGND VGND VPWR VPWR net285
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[52\] VGND VGND VPWR VPWR net296
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_89_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2282__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2830_ _0665_ _0663_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_100_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2761_ _0594_ _0596_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__nor2_2
XFILLER_0_26_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2692_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[34\]
+ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_14_CLK_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1 _1540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2700__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3313_ _1145_ _1146_ _0995_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__a21bo_1
X_3244_ _1072_ _1074_ _1078_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_29_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3175_ _1007_ _1009_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2126_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.rollover_flag VGND VGND VPWR VPWR _1548_
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_1_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout164_A net169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2057_ net222 net50 net85 VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2273__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2959_ _0481_ _0484_ _0794_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1925__S net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2610__A _1621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout77_A _1537_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_41_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_41_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2255__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3931_ clknet_leaf_35_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[8\] net141
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3862_ clknet_leaf_17_CLK _0188_ net168 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2813_ _0465_ _0648_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_42_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3793_ clknet_leaf_18_CLK _0119_ net167 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2744_ _1618_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\] VGND VGND VPWR
+ VPWR _0580_ sky130_fd_sc_hd__nor2_1
X_2675_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\] _1648_ _0510_ VGND
+ VGND VPWR VPWR _0511_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3227_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[46\]
+ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__nand2b_1
XANTENNA__3261__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2148__Y _1570_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3158_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[62\]
+ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__nor2_1
X_2109_ net232 net56 net83 VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__mux2_1
X_3089_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[24\] _0908_ _0912_ _0921_ _0924_
+ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_92_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2605__A _1623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_23_CLK clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_23_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2515__A _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_CLK clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_14_CLK sky130_fd_sc_hd__clkbuf_8
X_2460_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[11\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[11\]
+ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__xor2_1
X_2391_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] _1781_ _1713_ VGND VGND VPWR
+ VPWR _1785_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3012_ _0577_ _0792_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3914_ clknet_leaf_3_CLK _0240_ net151 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[63\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_46_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3845_ clknet_leaf_4_CLK _0171_ net152 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3776_ clknet_leaf_10_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[23\]
+ net158 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_14_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2400__A0 myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_2727_ _0562_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2160__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2658_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[16\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[48\]
+ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__nand2_1
Xfanout102 _1535_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__buf_4
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2589_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\] _0371_ VGND VGND VPWR
+ VPWR _0426_ sky130_fd_sc_hd__nor2_1
Xfanout113 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[12\] VGND VGND VPWR VPWR net113
+ sky130_fd_sc_hd__buf_2
Xfanout124 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] VGND VGND VPWR VPWR net124
+ sky130_fd_sc_hd__buf_2
XFILLER_0_10_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout146 net148 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_4
Xfanout135 net136 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input1_A addr[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout157 net158 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_4
Xfanout168 net169 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3166__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input57_A wdata[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2458__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_3_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_3_CLK sky130_fd_sc_hd__clkbuf_8
X_1960_ net272 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[62\] net98 VGND
+ VGND VPWR VPWR _0109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1891_ net319 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] net102 VGND
+ VGND VPWR VPWR _0043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3630_ _1558_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[40\] VGND VGND VPWR
+ VPWR _1465_ sky130_fd_sc_hd__nand2_1
X_3561_ _1080_ _1081_ VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3076__A myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_2512_ net114 _0370_ _0372_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[9\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3492_ _0994_ _0996_ _1326_ _0993_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__a31o_1
X_2443_ _1608_ net115 VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__nor2_1
X_2374_ net72 _1771_ _1772_ VGND VGND VPWR VPWR _1773_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_22_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3828_ clknet_leaf_19_CLK _0154_ net167 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_50_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3759_ clknet_leaf_12_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[6\] net161
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1933__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2004__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2090_ net222 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[56\] net90 VGND
+ VGND VPWR VPWR _0233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2992_ _0796_ _0798_ _0590_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1943_ net265 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[45\] net101 VGND
+ VGND VPWR VPWR _0092_ sky130_fd_sc_hd__mux2_1
X_3613_ _1390_ _1446_ _1447_ VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1874_ net233 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] net105 VGND
+ VGND VPWR VPWR _0026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3544_ _1098_ _1378_ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__xor2_1
X_3475_ _1289_ _1308_ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__and2b_1
XFILLER_0_12_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2426_ _1584_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[26\] _1783_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\]
+ _0295_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3331__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_2357_ net72 _1759_ _1760_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[19\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2288_ _1700_ _1702_ _1704_ _1709_ VGND VGND VPWR VPWR _1710_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_27_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1928__S net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2412__A1_N myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3937__RESET_B net144 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3322__A1 _1592_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1884__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2061__A1 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2523__A _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3260_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\]
+ VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3191_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] _1666_ VGND VGND VPWR
+ VPWR _1026_ sky130_fd_sc_hd__and2_1
X_2211_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.count_enable VGND VGND VPWR VPWR _1633_
+ sky130_fd_sc_hd__inv_2
X_2142_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[14\] VGND VGND VPWR VPWR _1564_
+ sky130_fd_sc_hd__inv_2
X_2073_ net298 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[39\] net93 VGND
+ VGND VPWR VPWR _0216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2052__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2975_ _0461_ _0810_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1926_ net295 net55 net77 VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1857_ net297 net54 net81 VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1788_ net124 _1661_ _1663_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[9\] VGND VGND
+ VPWR VPWR _1477_ sky130_fd_sc_hd__o22a_1
X_3527_ net119 _1353_ _1359_ net120 _1360_ VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3458_ _1075_ _1077_ _1292_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[44\]
+ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\] VGND VGND VPWR VPWR _1293_
+ sky130_fd_sc_hd__a32o_1
X_3389_ _1222_ _1223_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__and2_1
X_2409_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] _1740_ VGND VGND VPWR
+ VPWR _0279_ sky130_fd_sc_hd__xnor2_1
XANTENNA__1866__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3991__186 VGND VGND VPWR VPWR _3991__186/HI net186 sky130_fd_sc_hd__conb_1
XFILLER_0_82_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2043__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3771__RESET_B net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3700__RESET_B net144 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1857__A1 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold71 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[7\] VGND VGND VPWR VPWR net275
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[58\] VGND VGND VPWR VPWR net286
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[30\] VGND VGND VPWR VPWR net264
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_89_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold93 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[28\] VGND VGND VPWR VPWR net297
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2034__A1 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2760_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[60\]
+ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_584 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2691_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[34\]
+ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3312_ _0995_ _1144_ _1146_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__or3b_1
XFILLER_0_21_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3243_ _1076_ _1077_ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__nand2_2
XANTENNA__1848__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3174_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[55\]
+ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__nor2_1
XANTENNA__2428__A _1562_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2125_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.rollover_flag VGND VGND VPWR VPWR _1547_
+ sky130_fd_sc_hd__inv_2
X_2056_ net266 net49 net86 VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__mux2_1
XANTENNA__2273__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout157_A net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2273__B2 _1594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2025__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2958_ _0573_ _0576_ _0572_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_72_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1909_ net263 net37 net80 VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__mux2_1
X_2889_ _0715_ _0718_ _0724_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_9_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1941__S net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2016__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_3__f_CLK_A clknet_0_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2012__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input42_X net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1851__S net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2255__A1 _1562_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3930_ clknet_leaf_33_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[7\] net141
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3861_ clknet_leaf_18_CLK _0187_ net168 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2007__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2812_ _0470_ _0647_ _0467_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_42_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3792_ clknet_leaf_21_CLK _0118_ net162 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2743_ _0578_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2674_ _1606_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[39\] VGND VGND VPWR
+ VPWR _0510_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3226_ _1059_ _1060_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__nor2_2
XFILLER_0_94_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2158__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3157_ _1650_ _0991_ _0992_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.pwm_next
+ sky130_fd_sc_hd__a21oi_1
X_2108_ net307 net45 net83 VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__mux2_1
X_3088_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] _0831_ _0911_ VGND VGND VPWR
+ VPWR _0924_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_76_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2039_ net242 net62 net87 VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1936__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3997__192 VGND VGND VPWR VPWR _3997__192/HI net192 sky130_fd_sc_hd__conb_1
XFILLER_0_99_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_13_CLK_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2007__S net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_28_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2531__A _0351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2390_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[28\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\]
+ _1779_ VGND VGND VPWR VPWR _1784_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2249__Y _1671_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3011_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] _0844_ _0846_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\]
+ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_19_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Left_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3913_ clknet_leaf_3_CLK _0239_ net151 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[62\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_58_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3844_ clknet_leaf_5_CLK _0170_ net152 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3775_ clknet_leaf_10_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[22\]
+ net158 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[22\] sky130_fd_sc_hd__dfrtp_2
X_2726_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] _1645_ _0505_ _0559_
+ _0561_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__a221o_1
X_2657_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[16\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[48\]
+ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2588_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] _0361_ _0365_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\]
+ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__a22o_1
Xfanout103 _1535_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__buf_2
Xfanout125 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[6\] VGND VGND VPWR VPWR net125
+ sky130_fd_sc_hd__buf_2
Xfanout114 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[9\] VGND VGND VPWR VPWR net114
+ sky130_fd_sc_hd__buf_2
Xfanout147 net148 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_4
Xfanout136 net138 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
Xfanout158 net170 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_4
Xfanout169 net170 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__buf_2
X_3209_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[37\]
+ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout92_X net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2458__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1890_ net297 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] net102 VGND
+ VGND VPWR VPWR _0042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3560_ _1306_ _1307_ _1290_ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2261__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2511_ net114 _0370_ net70 VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3491_ _1323_ _1324_ _1325_ _0998_ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__o31ai_4
X_2442_ _1625_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[26\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\]
+ _1632_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__a22o_1
X_2373_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[24\]
+ _1767_ VGND VGND VPWR VPWR _1772_ sky130_fd_sc_hd__and3_1
XANTENNA__2697__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3827_ clknet_leaf_17_CLK _0153_ net168 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_61_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3758_ clknet_leaf_23_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[5\] net161
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__2171__A net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2709_ _0542_ _0544_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__nand2_2
X_3689_ clknet_leaf_33_CLK _0049_ net140 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2110__S net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2612__B2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3177__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2020__S net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2991_ _0812_ _0826_ _0814_ _0815_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__or4b_1
XFILLER_0_29_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1942_ net263 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[44\] net101 VGND
+ VGND VPWR VPWR _0091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1873_ net218 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[11\] net105 VGND
+ VGND VPWR VPWR _0025_ sky130_fd_sc_hd__mux2_1
X_3612_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] _1375_ _1379_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\]
+ _1376_ VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3543_ _1103_ _1377_ _1102_ VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__a21bo_1
X_3474_ _1306_ _1308_ _1293_ VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2425_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] _1773_ _0292_ _0293_
+ _0294_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__a2111o_1
X_2356_ net121 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] _1756_ VGND VGND VPWR
+ VPWR _1760_ sky130_fd_sc_hd__and3_1
XANTENNA__1819__A1_N _1594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2287_ _1705_ _1706_ _1707_ _1708_ VGND VGND VPWR VPWR _1709_ sky130_fd_sc_hd__and4b_1
XFILLER_0_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2172__Y _1594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1944__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2015__S net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1854__S net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2210_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[31\] VGND VGND VPWR VPWR _1632_
+ sky130_fd_sc_hd__inv_2
X_3190_ _1023_ _1024_ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__or2_2
X_2141_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\] VGND VGND VPWR VPWR _1563_
+ sky130_fd_sc_hd__inv_2
X_2072_ net242 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[38\] net92 VGND
+ VGND VPWR VPWR _0215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2974_ _0621_ _0636_ _0809_ _0635_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1925_ net313 net54 net77 VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1856_ net308 net53 net81 VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1787_ _1465_ _1474_ _1475_ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__a21bo_1
X_3526_ net120 _1359_ VGND VGND VPWR VPWR _1361_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout102_A _1535_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3457_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[11\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[43\]
+ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[42\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\]
+ _1290_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__a221o_1
X_3388_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[22\] _1221_ VGND VGND VPWR VPWR
+ _1223_ sky130_fd_sc_hd__nand2_1
X_2408_ _1566_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[16\] _0271_ _0274_
+ _0275_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__o2111ai_1
X_2339_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[14\] _1746_ VGND VGND VPWR VPWR
+ _1748_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_68_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4009_ net204 VGND VGND VPWR VPWR request_stall sky130_fd_sc_hd__buf_2
XFILLER_0_67_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1939__S net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input32_A addr[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold50 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[3\] VGND VGND VPWR VPWR net254
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[19\] VGND VGND VPWR VPWR net287
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[52\] VGND VGND VPWR VPWR net276
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold61 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[45\] VGND VGND VPWR VPWR net265
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[39\] VGND VGND VPWR VPWR net298
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_11_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1849__S net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2690_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[34\]
+ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3311_ _1590_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[61\] VGND VGND VPWR
+ VPWR _1146_ sky130_fd_sc_hd__or2_1
XANTENNA__3899__RESET_B net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3242_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[11\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[43\]
+ VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__or2_1
X_3173_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[55\]
+ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__nand2_1
X_2124_ net251 net42 net82 VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2411__A1_N myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2055_ net321 net48 net86 VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3470__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2957_ _0574_ _0577_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2888_ _0677_ _0680_ _0720_ _0723_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__or4b_1
X_1908_ net219 net36 net80 VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__mux2_1
X_1839_ net28 net30 net29 net32 VGND VGND VPWR VPWR _1527_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3275__A _1570_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout105_X net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3509_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] _1338_ _1339_ _1343_ VGND VGND
+ VPWR VPWR _1344_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3213__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3185__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input35_X net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3974__171 VGND VGND VPWR VPWR _3974__171/HI net171 sky130_fd_sc_hd__conb_1
XFILLER_0_53_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3452__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3860_ clknet_leaf_19_CLK _0186_ net167 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_2811_ _0473_ _0586_ _0589_ _0475_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_39_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3791_ clknet_leaf_22_CLK _0117_ net162 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_70_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2742_ _0481_ _0484_ _0574_ _0577_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__and4_1
X_2673_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[42\]
+ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__xor2_4
XFILLER_0_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3225_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[45\]
+ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2439__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3156_ _1650_ _0991_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.count_enable VGND VGND
+ VPWR VPWR _0992_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2107_ net205 net34 net83 VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__mux2_1
X_3087_ _0917_ _0922_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2038_ net268 net61 net87 VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2174__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3989_ net184 VGND VGND VPWR VPWR rdata[12] sky130_fd_sc_hd__buf_2
XFILLER_0_17_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2113__S net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1952__S net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout82_A _1534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1996__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2023__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1862__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1920__A1 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2259__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3010_ _0574_ _0845_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_19_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3912_ clknet_leaf_4_CLK _0238_ net150 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[61\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1987__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3843_ clknet_leaf_4_CLK _0169_ net150 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_73_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3774_ clknet_leaf_10_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[21\]
+ net158 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2725_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] _1645_ _0560_ VGND
+ VGND VPWR VPWR _0561_ sky130_fd_sc_hd__o21a_1
X_2656_ _0489_ _0490_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__nand2_1
Xfanout104 _1535_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__buf_4
X_2587_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[11\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[11\]
+ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__xor2_1
Xfanout126 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[4\] VGND VGND VPWR VPWR net126
+ sky130_fd_sc_hd__buf_2
XFILLER_0_10_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1911__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout115 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\] VGND VGND VPWR VPWR net115
+ sky130_fd_sc_hd__buf_2
Xfanout137 net138 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2169__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xfanout159 net161 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_4
Xfanout148 net149 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__buf_2
X_3208_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[37\]
+ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__and2_1
X_3139_ net115 _1648_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[39\] _1607_
+ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__2108__S net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1978__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1947__S net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2632__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout85_X net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2018__S net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1969__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_466 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1857__S net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3490_ _1131_ _1134_ _1322_ _1133_ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__a211oi_2
XANTENNA__2394__A1 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2510_ _0371_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[8\]
+ sky130_fd_sc_hd__inv_2
X_2441_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] net113 VGND VGND VPWR
+ VPWR _0310_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2372_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[24\] _1769_ VGND VGND VPWR VPWR
+ _1771_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_3_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2717__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3826_ clknet_leaf_20_CLK _0152_ net164 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout132_A net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3757_ clknet_leaf_23_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[4\] net161
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2708_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[38\]
+ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_12_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3688_ clknet_leaf_31_CLK _0048_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_2639_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] _1637_ _0474_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\]
+ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__a22oi_2
XANTENNA__1896__B1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2627__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[24\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_67_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3765__RESET_B net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2362__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_80_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input62_A wdata[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_76_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_85_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2990_ _0820_ _0825_ _0818_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__or3b_1
XFILLER_0_83_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1941_ net219 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[43\] net101 VGND
+ VGND VPWR VPWR _0090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1872_ net326 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] net104 VGND
+ VGND VPWR VPWR _0024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3611_ _1440_ _1443_ _1445_ VGND VGND VPWR VPWR _1446_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3542_ _1315_ _1317_ VGND VGND VPWR VPWR _1377_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3473_ _1078_ _1307_ _1075_ VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__and3b_1
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2119__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2424_ _1584_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[26\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[24\]
+ _1580_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2355_ net121 _1756_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR
+ VPWR _1759_ sky130_fd_sc_hd__a21oi_1
X_2286_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\]
+ VGND VGND VPWR VPWR _1708_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3809_ clknet_leaf_6_CLK _0135_ net155 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2121__S net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1960__S net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2357__A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3188__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input65_X net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1870__S net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2140_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\] VGND VGND VPWR VPWR
+ _1562_ sky130_fd_sc_hd__inv_2
X_2071_ net268 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[37\] net92 VGND
+ VGND VPWR VPWR _0214_ sky130_fd_sc_hd__mux2_1
X_2973_ _0805_ _0806_ _0807_ _0622_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__a31o_1
XFILLER_0_56_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2588__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2588__B2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_1924_ net299 net53 net77 VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1855_ net234 net52 net81 VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1786_ _1559_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[41\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[40\]
+ _1558_ VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3525_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[24\] _1357_ _1359_ net120 VGND VGND
+ VPWR VPWR _1360_ sky130_fd_sc_hd__a22o_1
X_3456_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[42\]
+ _1290_ VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__a21o_1
X_2407_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[11\] _1743_ VGND VGND VPWR
+ VPWR _0277_ sky130_fd_sc_hd__xnor2_1
X_3387_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[22\] _1221_ VGND VGND VPWR VPWR
+ _1222_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2338_ _1747_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[13\]
+ sky130_fd_sc_hd__inv_2
X_2269_ _1680_ _1686_ _1688_ _1690_ VGND VGND VPWR VPWR _1691_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_68_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4008_ net203 VGND VGND VPWR VPWR rdata[31] sky130_fd_sc_hd__buf_2
XFILLER_0_67_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2116__S net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1955__S net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold40 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[4\] VGND VGND VPWR VPWR net244
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[49\] VGND VGND VPWR VPWR net277
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A addr[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold62 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[55\] VGND VGND VPWR VPWR net266
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[34\] VGND VGND VPWR VPWR net255
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[22\] VGND VGND VPWR VPWR net288
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[59\] VGND VGND VPWR VPWR net299
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2267__B1 _1570_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3780__RESET_B net154 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2026__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1865__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_44_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_44_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_41_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3310_ _1139_ _1143_ _0998_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3241_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[11\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[43\]
+ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__nand2_1
X_3172_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[55\]
+ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__and2_1
X_2123_ net229 net41 net82 VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2054_ net305 net47 net85 VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2956_ _0786_ _0787_ _0791_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2887_ net112 _0679_ _0717_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[11\] _0719_
+ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__o221a_1
X_1907_ net208 net35 net79 VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1838_ net31 net3 net2 net5 VGND VGND VPWR VPWR _1526_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_35_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_35_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3508_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[28\] _1335_ VGND VGND VPWR VPWR
+ _1343_ sky130_fd_sc_hd__or2_1
X_3439_ _1264_ _1270_ _1273_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__nor3b_1
XANTENNA__3291__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2635__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_531 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_26_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_26_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3790_ clknet_leaf_20_CLK _0116_ net164 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2810_ _0586_ _0589_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_70_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2741_ _0575_ _0576_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__nand2_2
Xclkbuf_leaf_17_CLK clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_17_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2672_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[42\]
+ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3981__176 VGND VGND VPWR VPWR _3981__176/HI net176 sky130_fd_sc_hd__conb_1
X_3224_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[45\]
+ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__and2_1
.ends


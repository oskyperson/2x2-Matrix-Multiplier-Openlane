* NGSPICE file created from calculator_top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

.subckt calculator_top ColOut[0] ColOut[1] ColOut[2] ColOut[3] RowIn[0] RowIn[1] RowIn[2]
+ RowIn[3] VGND VPWR clk complete display_output[0] display_output[10] display_output[11]
+ display_output[12] display_output[13] display_output[14] display_output[15] display_output[1]
+ display_output[2] display_output[3] display_output[4] display_output[5] display_output[6]
+ display_output[7] display_output[8] display_output[9] input_state_FPGA[0] input_state_FPGA[1]
+ input_state_FPGA[2] key_pressed nRST
X_2106_ input_ctrl_inst.debounce_cnt\[11\] input_ctrl_inst.debounce_cnt\[10\] _1155_
+ VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__and3_1
XFILLER_39_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2037_ gencon_inst.mult_calc.compCount.in2\[5\] _1100_ _1103_ gencon_inst.mult_calc.compCount.in2\[6\]
+ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__a22o_1
XFILLER_62_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1270_ gencon_inst.operand1\[7\] net45 _0604_ _0605_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__o22a_1
XFILLER_51_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2724_ clknet_leaf_17_clk _0268_ net153 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[3\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1606_ net109 gencon_inst.add_calc.main.in2\[4\] VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__or2_1
X_2655_ clknet_leaf_33_clk _0204_ net126 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2586_ clknet_leaf_11_clk _0001_ net136 VGND VGND VPWR VPWR gencon_inst.add_calc.state\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1399_ gencon_inst.ALU_in2\[15\] gencon_inst.ALU_in1\[15\] VGND VGND VPWR VPWR _0696_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_47_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout138 net5 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_2
X_1537_ net415 net90 _0759_ net102 VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__a22o_1
Xfanout149 net150 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_4
X_1468_ gencon_inst.mult_calc.main.a0.in2 gencon_inst.mult_calc.main.a0.in1 VGND VGND
+ VPWR VPWR _0701_ sky130_fd_sc_hd__nand2_1
Xfanout127 net130 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_4
Xfanout116 input_ctrl_inst.col_index\[2\] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
Xfanout105 gencon_inst.mult_calc.next_finish VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_4
XFILLER_42_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold170 _0181_ VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold181 _0212_ VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 gencon_inst.mult_calc.compCount.in2\[14\] VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2440_ input_ctrl_inst.col_index\[30\] _0528_ _0551_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__and3_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1253_ net72 _0590_ net43 VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__a21o_1
X_1322_ gencon_inst.operand2\[2\] gencon_inst.latched_keypad_input\[2\] VGND VGND
+ VPWR VPWR _0648_ sky130_fd_sc_hd__or2_1
X_2371_ input_ctrl_inst.col_index\[8\] _0509_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__nor2_1
XFILLER_64_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2707_ clknet_leaf_11_clk _0251_ net136 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2569_ clknet_leaf_5_clk _0122_ net128 VGND VGND VPWR VPWR gencon_inst.operand2\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_2638_ clknet_leaf_36_clk _0187_ net126 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.a0.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1871_ gencon_inst.operand1\[15\] net435 net46 VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__mux2_1
X_1940_ gencon_inst.operand2\[0\] net51 net34 net344 VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__a22o_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2423_ input_ctrl_inst.col_index\[25\] input_ctrl_inst.col_index\[26\] _0540_ VGND
+ VGND VPWR VPWR _0544_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_67_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1305_ gencon_inst.operand1\[14\] net44 _0632_ _0633_ VGND VGND VPWR VPWR _0121_
+ sky130_fd_sc_hd__o22a_1
XFILLER_49_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1236_ _0576_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__inv_2
X_2285_ input_ctrl_inst.scan_timer\[9\] input_ctrl_inst.scan_timer\[11\] input_ctrl_inst.scan_timer\[10\]
+ _0461_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__and4_1
X_2354_ net116 _0411_ _0429_ _0432_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__or4_1
XFILLER_52_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2070_ _1054_ _1055_ _1064_ _1132_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__a22o_1
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1785_ net362 _0956_ net112 VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__mux2_1
X_1854_ gencon_inst.operand2\[14\] net250 net49 VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__mux2_1
X_1923_ gencon_inst.operand1\[10\] _0378_ net61 gencon_inst.mult_calc.out\[10\] VGND
+ VGND VPWR VPWR _1018_ sky130_fd_sc_hd__a22o_1
XFILLER_69_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2406_ _0527_ _0532_ _0529_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__o21ai_1
XFILLER_69_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1219_ net93 _0561_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__nor2_1
X_2268_ input_ctrl_inst.scan_timer\[1\] input_ctrl_inst.scan_timer\[2\] _0439_ input_ctrl_inst.scan_timer\[3\]
+ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__a31o_1
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2337_ net94 net243 net78 gencon_inst.mult_calc.count.GENERATE_ADDER\[4\].thingy.in1
+ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__a22o_1
X_2199_ net117 input_ctrl_inst.col_index\[1\] net116 input_ctrl_inst.col_index\[3\]
+ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__or4_1
XFILLER_71_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold52 gencon_inst.ALU_in2\[13\] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 _0308_ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 gencon_inst.prev_operator_input\[1\] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 input_ctrl_inst.scan_timer\[17\] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold74 _0073_ VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_71_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold96 gencon_inst.ALU_in2\[0\] VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold85 input_ctrl_inst.scan_timer\[16\] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1570_ net107 gencon_inst.add_calc.main.in2\[13\] VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__or2_1
XFILLER_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2122_ _1053_ _1132_ _1169_ _1054_ _1055_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__a32o_1
XFILLER_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2053_ _1087_ _1116_ _1119_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__o21ai_1
X_1768_ gencon_inst.ALU_in2\[5\] gencon_inst.ALU_in1\[5\] net65 VGND VGND VPWR VPWR
+ _0948_ sky130_fd_sc_hd__mux2_1
X_1906_ net52 _0972_ net39 net21 VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__a22o_1
X_1837_ gencon_inst.read_input gencon_inst.operator_input\[2\] VGND VGND VPWR VPWR
+ _0987_ sky130_fd_sc_hd__and2b_1
X_1699_ _0849_ _0904_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__xnor2_1
XFILLER_57_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput20 net20 VGND VGND VPWR VPWR display_output[3] sky130_fd_sc_hd__buf_2
Xoutput7 net7 VGND VGND VPWR VPWR ColOut[1] sky130_fd_sc_hd__buf_2
XFILLER_63_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1622_ _0834_ _0836_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__nor2_1
X_2740_ clknet_leaf_35_clk _0284_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2671_ clknet_leaf_36_clk _0220_ net140 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1484_ gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in1
+ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__nand2_1
X_1553_ _0770_ _0771_ _0772_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__or3_1
X_2105_ input_ctrl_inst.debounce_cnt\[10\] net37 _1158_ _1159_ VGND VGND VPWR VPWR
+ _0009_ sky130_fd_sc_hd__a22o_1
X_2036_ _1077_ _1102_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__or2_1
XFILLER_50_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2723_ clknet_leaf_12_clk _0267_ net137 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[2\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1605_ gencon_inst.add_calc.main.GENERATE_ADDER\[5\].thingy.in1 _0817_ _0818_ VGND
+ VGND VPWR VPWR _0820_ sky130_fd_sc_hd__nand3_1
X_2585_ clknet_leaf_11_clk net110 net136 VGND VGND VPWR VPWR gencon_inst.add_calc.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1536_ _0756_ _0758_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__xnor2_1
X_2654_ clknet_leaf_37_clk _0203_ net126 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout106 net109 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__buf_2
Xfanout128 net130 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_4
Xfanout117 input_ctrl_inst.col_index\[0\] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
Xfanout139 net145 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_4
X_1398_ gencon_inst.mult_calc.state\[2\] _1084_ net89 net216 VGND VGND VPWR VPWR _0152_
+ sky130_fd_sc_hd__a22o_1
X_1467_ net352 net307 net100 VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__mux2_1
X_2019_ _1080_ _1085_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_19_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold171 gencon_inst.add_calc.main.in2\[11\] VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 gencon_inst.mult_calc.INn2\[13\] VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 input_ctrl_inst.scan_timer\[7\] VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in2 VGND VGND VPWR
+ VPWR net320 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_48_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1252_ _0590_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__inv_2
X_1321_ gencon_inst.operand2\[2\] gencon_inst.latched_keypad_input\[2\] VGND VGND
+ VPWR VPWR _0647_ sky130_fd_sc_hd__nand2_1
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2370_ _0507_ _0509_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__nor2_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2706_ clknet_leaf_11_clk _0250_ net136 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2568_ clknet_leaf_24_clk _0121_ net157 VGND VGND VPWR VPWR gencon_inst.operand1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_1519_ gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in1
+ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__nand2_1
X_2499_ clknet_leaf_32_clk net244 net139 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[4\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2637_ clknet_leaf_36_clk _0186_ net127 VGND VGND VPWR VPWR gencon_inst.mult_calc.finish
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1870_ gencon_inst.operand1\[14\] net241 net49 VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2422_ input_ctrl_inst.col_index\[25\] _0540_ input_ctrl_inst.col_index\[26\] VGND
+ VGND VPWR VPWR _0543_ sky130_fd_sc_hd__a21oi_1
X_2353_ net116 _0496_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__nand2_1
X_1304_ gencon_inst.ALU_out\[14\] net69 net56 gencon_inst.mult_calc.out\[14\] _0565_
+ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__a221o_1
X_1235_ gencon_inst.operand1\[2\] gencon_inst.latched_keypad_input\[2\] VGND VGND
+ VPWR VPWR _0576_ sky130_fd_sc_hd__nand2_1
XFILLER_37_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2284_ net398 _0463_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_50_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1999_ input_ctrl_inst.input_control_state\[2\] _1056_ net83 gencon_inst.key_read
+ _1054_ VGND VGND VPWR VPWR input_ctrl_inst.next_state\[2\] sky130_fd_sc_hd__a221o_1
XFILLER_75_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1922_ _1016_ _1017_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__or2_1
XFILLER_34_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1784_ gencon_inst.ALU_in2\[13\] gencon_inst.ALU_in1\[13\] net63 VGND VGND VPWR VPWR
+ _0956_ sky130_fd_sc_hd__mux2_1
X_1853_ gencon_inst.operand2\[13\] net212 net48 VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__mux2_1
XFILLER_69_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2336_ net94 net247 net78 gencon_inst.mult_calc.count.GENERATE_ADDER\[3\].thingy.in1
+ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__a22o_1
X_2405_ _0530_ _0531_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__or2_1
XFILLER_55_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1218_ gencon_inst.gencon_state\[3\] _1214_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__nand2_1
X_2267_ input_ctrl_inst.scan_timer\[1\] input_ctrl_inst.scan_timer\[3\] input_ctrl_inst.scan_timer\[2\]
+ _0439_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__and4_1
X_2198_ net117 input_ctrl_inst.col_index\[1\] net116 input_ctrl_inst.col_index\[3\]
+ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__nor4_1
XFILLER_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold64 gencon_inst.ALU_in1\[3\] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 gencon_inst.add_calc.start VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 gencon_inst.ALU_in1\[5\] VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 gencon_inst.mult_calc.INn1\[6\] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in1 VGND VGND VPWR VPWR
+ net191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 _0474_ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold20 gencon_inst.mult_calc.INn1\[0\] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold75 gencon_inst.mult_calc.countSave\[6\] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2121_ _1171_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__inv_2
XFILLER_34_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2052_ gencon_inst.mult_calc.compCount.in2\[11\] _1086_ _1118_ gencon_inst.mult_calc.compCount.in2\[12\]
+ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__o22a_1
X_1905_ gencon_inst.ALU_out\[4\] net71 net60 gencon_inst.mult_calc.out\[4\] VGND VGND
+ VPWR VPWR _1006_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1698_ _0799_ _0800_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__nand2b_1
X_1767_ net404 _0947_ net111 VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__mux2_1
X_1836_ net190 _0986_ _0962_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2319_ input_ctrl_inst.decoded_key\[0\] input_ctrl_inst.decoded_key\[2\] net83 VGND
+ VGND VPWR VPWR _0485_ sky130_fd_sc_hd__o21ai_1
XFILLER_45_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput10 net10 VGND VGND VPWR VPWR complete sky130_fd_sc_hd__buf_2
Xoutput21 net21 VGND VGND VPWR VPWR display_output[4] sky130_fd_sc_hd__buf_2
XFILLER_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput8 net8 VGND VGND VPWR VPWR ColOut[2] sky130_fd_sc_hd__buf_2
XFILLER_56_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1621_ gencon_inst.add_calc.main.GENERATE_ADDER\[1\].thingy.in1 _0833_ _0835_ VGND
+ VGND VPWR VPWR _0836_ sky130_fd_sc_hd__a21oi_1
X_2670_ clknet_leaf_35_clk _0219_ net129 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1552_ _0765_ _0767_ _0766_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__a21boi_1
XFILLER_8_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2104_ input_ctrl_inst.debounce_cnt\[10\] _1155_ _1156_ VGND VGND VPWR VPWR _1159_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_39_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1483_ gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in1
+ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__nor2_1
X_2035_ gencon_inst.mult_calc.count.GENERATE_ADDER\[6\].thingy.in1 _1076_ VGND VGND
+ VPWR VPWR _1102_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_20_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2799_ clknet_leaf_6_clk _0343_ net135 VGND VGND VPWR VPWR gencon_inst.operand1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1819_ gencon_inst.operand2\[10\] gencon_inst.operand1\[10\] net76 VGND VGND VPWR
+ VPWR _0978_ sky130_fd_sc_hd__mux2_1
XFILLER_42_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2722_ clknet_leaf_12_clk _0266_ net137 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[1\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1604_ _0817_ _0818_ gencon_inst.add_calc.main.GENERATE_ADDER\[5\].thingy.in1 VGND
+ VGND VPWR VPWR _0819_ sky130_fd_sc_hd__a21oi_1
Xfanout107 net109 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_2
X_2584_ clknet_leaf_10_clk _0000_ net136 VGND VGND VPWR VPWR gencon_inst.add_calc.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout118 net119 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_4
Xfanout129 net130 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
X_1535_ gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in1
+ _0757_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__o21bai_1
X_2653_ clknet_leaf_37_clk net268 net126 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1397_ net87 _1122_ net89 net233 VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__a2bb2o_1
X_1466_ net381 net342 net101 VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__mux2_1
XFILLER_23_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2018_ gencon_inst.mult_calc.count.GENERATE_ADDER\[10\].thingy.in1 _1079_ gencon_inst.mult_calc.count.GENERATE_ADDER\[11\].thingy.in1
+ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold194 gencon_inst.add_calc.main.GENERATE_ADDER\[6\].thingy.in1 VGND VGND VPWR VPWR
+ net354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 _0153_ VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 gencon_inst.add_calc.state\[0\] VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 gencon_inst.mult_calc.compCount.in2\[7\] VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 gencon_inst.mult_calc.state\[0\] VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1320_ _0638_ _0642_ _0641_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__o21bai_1
X_1251_ _0583_ _0586_ gencon_inst.operand1\[4\] VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__o21ai_1
XFILLER_49_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_20_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2705_ clknet_leaf_13_clk _0249_ net137 VGND VGND VPWR VPWR gencon_inst.ALU_out\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_2636_ clknet_leaf_29_clk net296 net147 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[14\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2567_ clknet_leaf_23_clk _0120_ net157 VGND VGND VPWR VPWR gencon_inst.operand1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1449_ net189 net177 net101 VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__mux2_1
X_1518_ gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in1
+ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__nor2_1
X_2498_ clknet_leaf_37_clk net248 net139 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[3\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1303_ _0630_ _0631_ _0558_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__and3b_1
X_2283_ net119 net59 _0461_ input_ctrl_inst.scan_timer\[9\] _0463_ VGND VGND VPWR
+ VPWR _0041_ sky130_fd_sc_hd__o221a_1
X_2421_ input_ctrl_inst.col_index\[25\] net58 _0528_ _0542_ VGND VGND VPWR VPWR _0100_
+ sky130_fd_sc_hd__a22o_1
X_2352_ net116 _0496_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__or2_1
XFILLER_64_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1234_ gencon_inst.operand1\[1\] _0575_ net44 VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__mux2_1
XFILLER_60_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1998_ net92 net196 _1067_ VGND VGND VPWR VPWR input_ctrl_inst.next_state\[1\] sky130_fd_sc_hd__a21oi_1
X_2619_ clknet_leaf_29_clk _0168_ net146 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1852_ gencon_inst.operand2\[12\] net225 net48 VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__mux2_1
X_1921_ net53 _0977_ net39 net26 VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__a22o_1
XFILLER_42_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1783_ net379 _0955_ net113 VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2266_ net375 _0452_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__xnor2_1
X_2404_ input_ctrl_inst.col_index\[20\] _0525_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__nor2_1
X_2335_ net94 net232 net78 net293 VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__a22o_1
X_1217_ gencon_inst.gencon_state\[3\] _1214_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__and2_1
X_2197_ net93 _1208_ _0394_ VGND VGND VPWR VPWR gencon_inst.next_state\[3\] sky130_fd_sc_hd__and3_1
XFILLER_37_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_33_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold43 gencon_inst.ALU_in1\[11\] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 gencon_inst.ALU_in2\[12\] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 gencon_inst.ALU_in2\[4\] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 gencon_inst.ALU_in1\[4\] VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 gencon_inst.keypad_input\[3\] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in1 VGND VGND VPWR
+ VPWR net181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold10 gencon_inst.mult_calc.main.GENERATE_ADDER\[14\].thingy.in1 VGND VGND VPWR
+ VPWR net170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 gencon_inst.mult_calc.countSave\[3\] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 _0066_ VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_51_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_60_Left_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2120_ input_ctrl_inst.debounce_cnt\[13\] input_ctrl_inst.debounce_cnt\[14\] _1163_
+ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__and3_1
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2051_ _1081_ _1117_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_60_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1904_ _1004_ _1005_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__or2_1
X_1835_ gencon_inst.read_input gencon_inst.operator_input\[1\] VGND VGND VPWR VPWR
+ _0986_ sky130_fd_sc_hd__and2b_1
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1697_ _0858_ _0902_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__nand2_1
X_1766_ gencon_inst.ALU_in2\[4\] gencon_inst.ALU_in1\[4\] net62 VGND VGND VPWR VPWR
+ _0947_ sky130_fd_sc_hd__mux2_1
X_2318_ input_ctrl_inst.decoded_key\[1\] input_ctrl_inst.decoded_key\[3\] _0483_ VGND
+ VGND VPWR VPWR _0484_ sky130_fd_sc_hd__nor3_1
X_2249_ input_ctrl_inst.scan_timer\[0\] net123 _1055_ net84 VGND VGND VPWR VPWR _0439_
+ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_23_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput11 net11 VGND VGND VPWR VPWR display_output[0] sky130_fd_sc_hd__buf_2
XFILLER_48_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput22 net22 VGND VGND VPWR VPWR display_output[5] sky130_fd_sc_hd__buf_2
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput9 net9 VGND VGND VPWR VPWR ColOut[3] sky130_fd_sc_hd__buf_2
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1620_ net106 gencon_inst.add_calc.main.a0.in1 gencon_inst.add_calc.main.in2\[0\]
+ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__mux2_1
X_1482_ net390 net91 _0712_ net103 VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__a22o_1
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1551_ gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in1
+ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__and2_1
X_2103_ net35 _1155_ input_ctrl_inst.debounce_cnt\[10\] VGND VGND VPWR VPWR _1158_
+ sky130_fd_sc_hd__a21o_1
XFILLER_54_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2034_ gencon_inst.mult_calc.compCount.in2\[4\] _1097_ _1100_ gencon_inst.mult_calc.compCount.in2\[5\]
+ _1098_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__o221a_1
X_2798_ clknet_leaf_5_clk _0342_ net128 VGND VGND VPWR VPWR gencon_inst.key_read sky130_fd_sc_hd__dfrtp_2
X_1818_ net179 _0977_ net42 VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1749_ net334 _0938_ net113 VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__mux2_1
XFILLER_45_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2721_ clknet_leaf_11_clk _0265_ net136 VGND VGND VPWR VPWR gencon_inst.add_calc.main.a0.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2652_ clknet_leaf_26_clk _0201_ net147 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[14\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1603_ net106 gencon_inst.add_calc.main.in2\[5\] VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__nand2_1
Xfanout108 net109 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_2
X_2583_ clknet_leaf_25_clk _0136_ net143 VGND VGND VPWR VPWR gencon_inst.operand2\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_1534_ _0738_ _0743_ _0746_ _0750_ _0744_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__o311a_1
Xfanout119 _1038_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__buf_2
X_1465_ net388 net374 net101 VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__mux2_1
XFILLER_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1396_ net87 _1118_ net89 net221 VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__a2bb2o_1
X_2017_ _1083_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__inv_2
XFILLER_23_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold151 gencon_inst.add_calc.main.in2\[1\] VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 gencon_inst.add_calc.main.in2\[14\] VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 gencon_inst.mult_calc.adderSave\[9\] VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold195 gencon_inst.mult_calc.INn2\[4\] VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 gencon_inst.mult_calc.INn2\[0\] VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _0209_ VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1250_ gencon_inst.operand1\[3\] net44 _0588_ _0589_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__o22a_1
XFILLER_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2704_ clknet_leaf_19_clk _0248_ net158 VGND VGND VPWR VPWR gencon_inst.ALU_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_2635_ clknet_leaf_29_clk net274 net148 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2566_ clknet_leaf_21_clk _0119_ net157 VGND VGND VPWR VPWR gencon_inst.operand1\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_1448_ net181 net169 net100 VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__mux2_1
X_1517_ net103 _0741_ _0742_ net279 net88 VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__a32o_1
X_2497_ clknet_leaf_32_clk _0062_ net139 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[2\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1379_ gencon_inst.operand2\[14\] _0689_ net74 VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_2_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2420_ input_ctrl_inst.col_index\[25\] _0540_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__xor2_1
Xfanout90 net91 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_2
X_1233_ gencon_inst.ALU_out\[1\] net68 net56 gencon_inst.mult_calc.out\[1\] _0574_
+ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__a221o_1
X_1302_ gencon_inst.operand1\[12\] gencon_inst.operand1\[13\] _0618_ gencon_inst.operand1\[14\]
+ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__a31o_1
XFILLER_49_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2282_ input_ctrl_inst.scan_timer\[9\] _0461_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__nand2_1
X_2351_ _0495_ _0496_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__nor2_1
XFILLER_52_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1997_ gencon_inst.key_read _1061_ _1063_ _1066_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__o211a_1
X_2549_ clknet_leaf_3_clk _0031_ net125 VGND VGND VPWR VPWR input_ctrl_inst.read_input_flag
+ sky130_fd_sc_hd__dfrtp_1
X_2618_ clknet_leaf_28_clk _0167_ net150 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_7_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1851_ gencon_inst.operand2\[11\] net211 net49 VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__mux2_1
X_1920_ gencon_inst.ALU_out\[9\] net69 net61 gencon_inst.mult_calc.out\[9\] VGND VGND
+ VPWR VPWR _1016_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_12_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1782_ gencon_inst.ALU_in2\[12\] gencon_inst.ALU_in1\[12\] net63 VGND VGND VPWR VPWR
+ _0955_ sky130_fd_sc_hd__mux2_1
X_2403_ input_ctrl_inst.col_index\[20\] _0525_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__and2_1
XFILLER_69_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1216_ net93 gencon_inst.gencon_state\[3\] gencon_inst.gencon_state\[2\] gencon_inst.gencon_state\[1\]
+ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__or4b_4
X_2196_ _0387_ _0389_ _0395_ _1212_ VGND VGND VPWR VPWR gencon_inst.next_state\[2\]
+ sky130_fd_sc_hd__a211o_1
X_2265_ _0452_ _0453_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__and2_1
XFILLER_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2334_ net94 net251 net78 gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.in1
+ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__a22o_1
XFILLER_40_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold11 gencon_inst.mult_calc.INn1\[2\] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in1 VGND VGND VPWR VPWR
+ net182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_20_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold55 gencon_inst.latched_operator_input\[2\] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 net16 VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold33 gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in1 VGND VGND VPWR VPWR
+ net193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in1 VGND VGND VPWR VPWR
+ net259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 input_ctrl_inst.col_index\[18\] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 _0063_ VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 gencon_inst.mult_calc.countSave\[5\] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_61_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2050_ gencon_inst.mult_calc.count.GENERATE_ADDER\[12\].thingy.in1 _1080_ VGND VGND
+ VPWR VPWR _1117_ sky130_fd_sc_hd__nor2_1
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1765_ net364 _0946_ net111 VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__mux2_1
X_1903_ net52 _0971_ net40 net20 VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__a22o_1
X_1834_ net175 _0985_ _0962_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__mux2_1
XFILLER_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1696_ _0892_ _0895_ _0899_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__or3_1
XFILLER_72_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2179_ gencon_inst.mult_calc.finish _0380_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__nor2_1
X_2317_ input_ctrl_inst.decoded_key\[0\] input_ctrl_inst.decoded_key\[2\] VGND VGND
+ VPWR VPWR _0483_ sky130_fd_sc_hd__nand2_1
X_2248_ input_ctrl_inst.scan_timer\[1\] input_ctrl_inst.scan_timer\[0\] input_ctrl_inst.scan_timer\[3\]
+ input_ctrl_inst.scan_timer\[2\] VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_23_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput12 net12 VGND VGND VPWR VPWR display_output[10] sky130_fd_sc_hd__buf_2
Xoutput23 net23 VGND VGND VPWR VPWR display_output[6] sky130_fd_sc_hd__buf_2
XFILLER_31_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1481_ _0709_ _0711_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__xnor2_1
X_1550_ gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in1
+ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__nor2_1
X_2102_ net413 net37 _1154_ _1157_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__a22o_1
XFILLER_54_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2033_ _1076_ _1099_ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__or2_1
X_1748_ gencon_inst.ALU_in1\[10\] gencon_inst.ALU_in2\[10\] net64 VGND VGND VPWR VPWR
+ _0938_ sky130_fd_sc_hd__mux2_1
X_2797_ clknet_leaf_6_clk _0341_ net132 VGND VGND VPWR VPWR gencon_inst.latched_keypad_input\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_1817_ gencon_inst.operand2\[9\] gencon_inst.operand1\[9\] net77 VGND VGND VPWR VPWR
+ _0977_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1679_ _0879_ _0881_ _0886_ net31 VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__o31ai_1
XFILLER_13_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1602_ net106 gencon_inst.add_calc.main.in2\[5\] VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__or2_1
X_2720_ clknet_leaf_16_clk _0264_ net154 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2582_ clknet_leaf_27_clk _0135_ net150 VGND VGND VPWR VPWR gencon_inst.operand2\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2651_ clknet_leaf_29_clk _0200_ net148 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
Xfanout109 gencon_inst.add_calc.diffSign VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_2
X_1533_ _0754_ _0755_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__and2b_1
X_1395_ net87 _1086_ net89 net276 VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__a2bb2o_1
X_1464_ net312 gencon_inst.mult_calc.INn2\[11\] net100 VGND VGND VPWR VPWR _0213_
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2016_ gencon_inst.mult_calc.count.GENERATE_ADDER\[14\].thingy.in1 _1082_ VGND VGND
+ VPWR VPWR _1083_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_30_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
Xhold130 gencon_inst.add_calc.main.in2\[7\] VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 gencon_inst.add_calc.main.in2\[10\] VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _0361_ VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 gencon_inst.mult_calc.adderSave\[12\] VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 gencon_inst.mult_calc.compCount.in2\[11\] VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in2 VGND VGND VPWR
+ VPWR net323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 gencon_inst.add_calc.main.GENERATE_ADDER\[10\].thingy.in1 VGND VGND VPWR
+ VPWR net356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_21_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_12_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_32_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2703_ clknet_leaf_21_clk _0247_ net158 VGND VGND VPWR VPWR gencon_inst.ALU_out\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_2565_ clknet_leaf_23_clk _0118_ net156 VGND VGND VPWR VPWR gencon_inst.operand1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1516_ _0737_ _0739_ _0740_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__a21o_1
X_2634_ clknet_leaf_28_clk net288 net149 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
X_1378_ gencon_inst.operand2\[14\] _0689_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__and2_1
X_1447_ net193 net179 net101 VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__mux2_1
X_2496_ clknet_leaf_37_clk _0061_ net126 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout80 _1068_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_4
Xfanout91 _0695_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_2
X_1232_ _0572_ _0573_ net72 VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__and3b_1
X_1301_ gencon_inst.operand1\[13\] gencon_inst.operand1\[14\] _0622_ VGND VGND VPWR
+ VPWR _0630_ sky130_fd_sc_hd__and3_1
XFILLER_49_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2281_ _0445_ _0460_ _0462_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
X_2350_ net117 input_ctrl_inst.col_index\[1\] _0444_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__and3_1
XFILLER_64_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1996_ net30 _1058_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__nand2_1
X_2548_ clknet_leaf_2_clk net92 net124 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dfrtp_1
X_2617_ clknet_leaf_26_clk _0166_ net150 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_7_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2479_ clknet_leaf_10_clk _0010_ net133 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload0 clknet_2_0__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_66_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1781_ net361 _0954_ net113 VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__mux2_1
X_1850_ gencon_inst.operand2\[10\] net292 net48 VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2333_ net94 net228 net78 gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.cIn
+ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__a22o_1
X_2402_ net428 net59 VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__nand2_1
X_2195_ net73 _0386_ _0396_ VGND VGND VPWR VPWR gencon_inst.next_state\[1\] sky130_fd_sc_hd__or3_1
X_2264_ input_ctrl_inst.scan_timer\[1\] _0439_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__or2_1
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1979_ input_ctrl_inst.debounce_cnt\[14\] _1050_ _1046_ VGND VGND VPWR VPWR _1051_
+ sky130_fd_sc_hd__o21a_2
XFILLER_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold45 net14 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in1 VGND VGND VPWR VPWR
+ net183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 gencon_inst.mult_calc.INn1\[5\] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 gencon_inst.mult_calc.countSave\[14\] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 gencon_inst.mult_calc.main.a0.in1 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold89 gencon_inst.ALU_in1\[0\] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold67 gencon_inst.mult_calc.count.GENERATE_ADDER\[12\].thingy.in1 VGND VGND VPWR
+ VPWR net227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 _0065_ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1902_ gencon_inst.ALU_out\[3\] net68 net60 gencon_inst.mult_calc.out\[3\] VGND VGND
+ VPWR VPWR _1004_ sky130_fd_sc_hd__a22o_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1764_ gencon_inst.ALU_in2\[3\] gencon_inst.ALU_in1\[3\] net62 VGND VGND VPWR VPWR
+ _0946_ sky130_fd_sc_hd__mux2_1
X_1833_ gencon_inst.read_input _1031_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__nor2_1
XFILLER_30_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1695_ _0901_ _0900_ gencon_inst.ALU_out\[9\] net85 VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__a2bb2o_1
X_2316_ input_ctrl_inst.input_control_state\[2\] _1055_ _1056_ _1187_ net118 VGND
+ VGND VPWR VPWR _0482_ sky130_fd_sc_hd__a311oi_4
XFILLER_65_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2178_ _0380_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__inv_2
X_2247_ input_ctrl_inst.scan_timer\[5\] input_ctrl_inst.scan_timer\[7\] input_ctrl_inst.scan_timer\[6\]
+ input_ctrl_inst.scan_timer\[4\] VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__or4bb_1
XFILLER_25_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput24 net24 VGND VGND VPWR VPWR display_output[7] sky130_fd_sc_hd__buf_2
Xoutput13 net13 VGND VGND VPWR VPWR display_output[11] sky130_fd_sc_hd__buf_2
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1480_ _0704_ _0710_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__or2_1
X_2101_ _1155_ _1156_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2032_ gencon_inst.mult_calc.count.GENERATE_ADDER\[4\].thingy.in1 _1075_ gencon_inst.mult_calc.count.GENERATE_ADDER\[5\].thingy.in1
+ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__a21oi_1
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1747_ net318 _0937_ net113 VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__mux2_1
X_1678_ net445 _0887_ net114 VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2796_ clknet_leaf_6_clk _0340_ net132 VGND VGND VPWR VPWR gencon_inst.latched_keypad_input\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1816_ net178 _0976_ net42 VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_39_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1601_ gencon_inst.add_calc.main.GENERATE_ADDER\[6\].thingy.in1 _0813_ _0814_ VGND
+ VGND VPWR VPWR _0816_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_57_Left_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2581_ clknet_leaf_27_clk _0134_ net149 VGND VGND VPWR VPWR gencon_inst.operand2\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_1532_ gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in1
+ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__nand2_1
X_2650_ clknet_leaf_28_clk _0199_ net149 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1394_ net87 _1114_ net89 net269 VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__a2bb2o_1
X_1463_ net340 gencon_inst.mult_calc.INn2\[10\] net100 VGND VGND VPWR VPWR _0212_
+ sky130_fd_sc_hd__mux2_1
X_2015_ gencon_inst.mult_calc.count.GENERATE_ADDER\[13\].thingy.in1 _1081_ VGND VGND
+ VPWR VPWR _1082_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_75_Left_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold197 gencon_inst.add_calc.main.GENERATE_ADDER\[8\].thingy.in1 VGND VGND VPWR VPWR
+ net357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold186 gencon_inst.ALU_in1\[8\] VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 gencon_inst.ALU_in2\[7\] VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__dlygate4sd3_1
X_2779_ clknet_leaf_16_clk _0323_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[5\] sky130_fd_sc_hd__dfxtp_1
Xhold142 gencon_inst.latched_operator_input\[0\] VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 gencon_inst.mult_calc.adderSave\[1\] VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 gencon_inst.mult_calc.count.GENERATE_ADDER\[9\].thingy.in1 VGND VGND VPWR
+ VPWR net280 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold153 _0213_ VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _0174_ VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2702_ clknet_leaf_21_clk _0246_ net158 VGND VGND VPWR VPWR gencon_inst.ALU_out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_2564_ clknet_leaf_22_clk _0117_ net156 VGND VGND VPWR VPWR gencon_inst.operand1\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_2633_ clknet_leaf_28_clk net337 net149 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
X_1515_ _0737_ _0739_ _0740_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__nand3_1
X_2495_ clknet_leaf_37_clk _0060_ net126 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.cIn
+ sky130_fd_sc_hd__dfrtp_2
X_1377_ gencon_inst.operand2\[13\] _0691_ net55 VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__mux2_1
X_1446_ net187 net178 net100 VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__mux2_1
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout70 net71 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_2
Xfanout92 input_ctrl_inst.input_control_state\[2\] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_2
XFILLER_6_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout81 _1068_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1231_ gencon_inst.operand1\[0\] gencon_inst.latched_keypad_input\[0\] _0569_ _0571_
+ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__a22o_1
X_1300_ gencon_inst.operand1\[13\] net45 _0629_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__o21a_1
X_2280_ _0461_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__inv_2
XFILLER_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1995_ _1051_ _1064_ _1062_ _1054_ VGND VGND VPWR VPWR input_ctrl_inst.next_state\[0\]
+ sky130_fd_sc_hd__a211o_1
X_2616_ clknet_leaf_26_clk _0165_ net150 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2478_ clknet_leaf_10_clk _0009_ net133 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_2547_ clknet_leaf_2_clk net196 net124 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dfrtp_1
X_1429_ net96 gencon_inst.mult_calc.adderSave\[8\] net305 net80 VGND VGND VPWR VPWR
+ _0179_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_7_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload1 clknet_2_1__leaf_clk VGND VGND VPWR VPWR clkload1/X sky130_fd_sc_hd__clkbuf_8
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1780_ gencon_inst.ALU_in2\[11\] gencon_inst.ALU_in1\[11\] net64 VGND VGND VPWR VPWR
+ _0954_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2332_ _0482_ _0493_ _0494_ net192 net118 VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__a32o_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2401_ net446 net58 _0526_ _0528_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__a22o_1
XFILLER_65_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2194_ gencon_inst.mult_calc.finish _0381_ _0387_ _0393_ _0395_ VGND VGND VPWR VPWR
+ _0396_ sky130_fd_sc_hd__a221o_1
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2263_ input_ctrl_inst.scan_timer\[1\] _0439_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_63_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1978_ _1048_ _1049_ input_ctrl_inst.debounce_cnt\[13\] VGND VGND VPWR VPWR _1050_
+ sky130_fd_sc_hd__o21a_1
XFILLER_20_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold46 gencon_inst.ALU_in2\[2\] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 net12 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 gencon_inst.prev_operator_input\[2\] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 gencon_inst.mult_calc.INn2\[1\] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 input_ctrl_inst.scan_timer\[19\] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold68 gencon_inst.mult_calc.countSave\[0\] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 _0152_ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1901_ _1002_ _1003_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__or2_1
X_1832_ gencon_inst.latched_operator_input\[0\] net262 net46 VGND VGND VPWR VPWR _0297_
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1763_ net338 _0945_ net110 VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__mux2_1
X_1694_ net31 _0897_ _0899_ net85 VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__a31o_1
XFILLER_57_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2315_ net401 net118 _0480_ _0481_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__a22o_1
X_2246_ input_ctrl_inst.scan_timer\[13\] input_ctrl_inst.scan_timer\[12\] input_ctrl_inst.scan_timer\[15\]
+ input_ctrl_inst.scan_timer\[14\] VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__or4bb_1
X_2177_ gencon_inst.gencon_state\[3\] _0379_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_11_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput14 net14 VGND VGND VPWR VPWR display_output[12] sky130_fd_sc_hd__buf_2
Xoutput25 net25 VGND VGND VPWR VPWR display_output[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_74_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2100_ _1053_ _1132_ net35 VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__a21oi_2
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2031_ gencon_inst.mult_calc.compCount.in2\[3\] _1088_ _1097_ gencon_inst.mult_calc.compCount.in2\[4\]
+ _1096_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__a221o_1
XFILLER_22_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2795_ clknet_leaf_6_clk _0339_ net134 VGND VGND VPWR VPWR gencon_inst.latched_keypad_input\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1815_ gencon_inst.operand2\[8\] gencon_inst.operand1\[8\] net77 VGND VGND VPWR VPWR
+ _0976_ sky130_fd_sc_hd__mux2_1
XFILLER_30_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1746_ gencon_inst.ALU_in1\[9\] gencon_inst.ALU_in2\[9\] net64 VGND VGND VPWR VPWR
+ _0937_ sky130_fd_sc_hd__mux2_1
X_1677_ _0884_ _0886_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2229_ input_ctrl_inst.col_index\[29\] input_ctrl_inst.col_index\[28\] input_ctrl_inst.col_index\[31\]
+ input_ctrl_inst.col_index\[30\] VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__and4_1
XFILLER_53_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1600_ _0813_ _0814_ gencon_inst.add_calc.main.GENERATE_ADDER\[6\].thingy.in1 VGND
+ VGND VPWR VPWR _0815_ sky130_fd_sc_hd__a21oi_1
X_2580_ clknet_leaf_23_clk _0133_ net149 VGND VGND VPWR VPWR gencon_inst.operand2\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_1531_ gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in1
+ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__nor2_1
XFILLER_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1462_ net409 net298 net100 VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__mux2_1
X_1393_ net86 _1111_ net89 net264 VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2014_ gencon_inst.mult_calc.count.GENERATE_ADDER\[12\].thingy.in1 _1080_ VGND VGND
+ VPWR VPWR _1081_ sky130_fd_sc_hd__and2_1
X_2778_ clknet_leaf_16_clk _0322_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold110 gencon_inst.latched_operator_input\[1\] VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 gencon_inst.add_calc.main.in2\[5\] VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__dlygate4sd3_1
X_1729_ net442 _0928_ net110 VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__mux2_1
Xhold187 gencon_inst.ALU_out\[15\] VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 gencon_inst.ALU_in2\[1\] VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 gencon_inst.ALU_in2\[10\] VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 gencon_inst.ALU_in1\[7\] VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 equal_input VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in2 VGND VGND VPWR
+ VPWR net336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in2 VGND VGND VPWR
+ VPWR net303 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2701_ clknet_leaf_19_clk _0245_ net158 VGND VGND VPWR VPWR gencon_inst.ALU_out\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2632_ clknet_leaf_28_clk net330 net149 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
X_2563_ clknet_leaf_24_clk _0116_ net157 VGND VGND VPWR VPWR gencon_inst.operand1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2494_ clknet_leaf_6_clk _0059_ VGND VGND VPWR VPWR gencon_inst.keypad_input\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1445_ net183 net167 net100 VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__mux2_1
X_1514_ _0731_ _0735_ _0732_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__o21ai_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1376_ _0689_ _0690_ gencon_inst.mult_calc.out\[13\] net67 VGND VGND VPWR VPWR _0691_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout60 _0997_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_4
Xfanout71 _0562_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout93 gencon_inst.gencon_state\[0\] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_2
Xfanout82 _1061_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_2
XFILLER_6_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1230_ gencon_inst.operand1\[0\] gencon_inst.latched_keypad_input\[0\] _0569_ _0571_
+ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__and4_1
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1994_ net92 _1063_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_15_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload30 clknet_leaf_15_clk VGND VGND VPWR VPWR clkload30/Y sky130_fd_sc_hd__inv_12
X_2615_ clknet_leaf_26_clk _0164_ net150 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2477_ clknet_leaf_9_clk _0026_ net133 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2546_ clknet_leaf_7_clk net252 net131 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfrtp_1
X_1428_ net94 net279 net294 net78 VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__a22o_1
X_1359_ gencon_inst.operand2\[9\] _0674_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__xor2_1
Xclkload2 clknet_2_3__leaf_clk VGND VGND VPWR VPWR clkload2/X sky130_fd_sc_hd__clkbuf_8
XFILLER_7_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2400_ _0451_ _0500_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__nor2_2
X_2331_ gencon_inst.keypad_input\[3\] _1060_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__or2_1
X_2262_ _0439_ _0440_ _0445_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_63_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2193_ net93 _0394_ _1207_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1977_ input_ctrl_inst.debounce_cnt\[9\] input_ctrl_inst.debounce_cnt\[11\] input_ctrl_inst.debounce_cnt\[10\]
+ input_ctrl_inst.debounce_cnt\[12\] VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__or4_1
X_2529_ clknet_leaf_39_clk _0090_ net120 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold47 gencon_inst.ALU_in1\[2\] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold69 gencon_inst.ALU_in1\[13\] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 gencon_inst.ALU_in2\[15\] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 input_ctrl_inst.input_control_state\[1\] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 _0051_ VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in1 VGND VGND VPWR VPWR
+ net185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1900_ net52 _0970_ net40 net19 VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__a22o_1
X_1831_ net119 gencon_inst.latched_operator_input\[2\] gencon_inst.latched_operator_input\[1\]
+ _0392_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__or4bb_2
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1693_ net31 _0897_ _0899_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__a21oi_1
X_1762_ gencon_inst.ALU_in2\[2\] gencon_inst.ALU_in1\[2\] net62 VGND VGND VPWR VPWR
+ _0945_ sky130_fd_sc_hd__mux2_1
XFILLER_65_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2176_ net93 _1214_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__nand2_1
X_2314_ _1042_ input_ctrl_inst.decoded_key\[2\] VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__nor2_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2245_ input_ctrl_inst.scan_timer\[17\] input_ctrl_inst.scan_timer\[16\] input_ctrl_inst.scan_timer\[19\]
+ input_ctrl_inst.scan_timer\[18\] VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__or4_1
XFILLER_53_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput26 net26 VGND VGND VPWR VPWR display_output[9] sky130_fd_sc_hd__buf_2
Xoutput15 net15 VGND VGND VPWR VPWR display_output[13] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2030_ gencon_inst.mult_calc.count.GENERATE_ADDER\[4\].thingy.in1 _1075_ VGND VGND
+ VPWR VPWR _1097_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1745_ net328 _0936_ net112 VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__mux2_1
X_2794_ clknet_leaf_6_clk _0338_ net132 VGND VGND VPWR VPWR gencon_inst.latched_keypad_input\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_1814_ net167 _0975_ net42 VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__mux2_1
XFILLER_30_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1676_ _0843_ _0885_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2159_ input_ctrl_inst.RowSync\[2\] _1199_ _1200_ _1201_ VGND VGND VPWR VPWR _1202_
+ sky130_fd_sc_hd__a31o_1
XFILLER_26_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2228_ _0424_ _0426_ _0421_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__a21bo_1
XFILLER_53_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_33_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_42_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1530_ net102 _0752_ _0753_ net300 net89 VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__a32o_1
X_1392_ net86 _1108_ net89 net254 VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__a2bb2o_1
X_1461_ net396 net366 net100 VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__mux2_1
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2013_ gencon_inst.mult_calc.count.GENERATE_ADDER\[11\].thingy.in1 gencon_inst.mult_calc.count.GENERATE_ADDER\[10\].thingy.in1
+ _1079_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__and3_1
XFILLER_50_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_15_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_33_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1728_ gencon_inst.ALU_in1\[0\] gencon_inst.ALU_in2\[0\] net62 VGND VGND VPWR VPWR
+ _0928_ sky130_fd_sc_hd__mux2_1
X_2777_ clknet_leaf_16_clk _0321_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[3\] sky130_fd_sc_hd__dfxtp_1
Xhold100 gencon_inst.ALU_in2\[3\] VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 gencon_inst.keypad_input\[2\] VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 gencon_inst.keypad_input\[1\] VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 _0175_ VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold133 gencon_inst.mult_calc.count.GENERATE_ADDER\[2\].thingy.in1 VGND VGND VPWR
+ VPWR net293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 gencon_inst.add_calc.main.in2\[3\] VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__dlygate4sd3_1
X_1659_ net32 _0869_ _0871_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__a21oi_1
Xhold188 gencon_inst.ALU_in1\[10\] VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 gencon_inst.mult_calc.INn2\[11\] VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 _0182_ VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in2 VGND VGND VPWR
+ VPWR net326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2700_ clknet_leaf_19_clk _0244_ net158 VGND VGND VPWR VPWR gencon_inst.ALU_out\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2562_ clknet_leaf_24_clk _0115_ net152 VGND VGND VPWR VPWR gencon_inst.operand1\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_2631_ clknet_leaf_28_clk _0180_ net150 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
X_2493_ clknet_leaf_6_clk _0058_ VGND VGND VPWR VPWR gencon_inst.keypad_input\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1375_ gencon_inst.operand2\[13\] _0686_ net74 VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_4_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
X_1513_ gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in1
+ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__nand2_1
X_1444_ net259 net213 net99 VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__mux2_1
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2829_ clknet_leaf_25_clk _0369_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout72 _0558_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_2
Xfanout61 _0997_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout83 _1060_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_2
Xfanout50 net51 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_2
XFILLER_13_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout94 gencon_inst.mult_calc.state\[4\] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_4
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1993_ net92 _1063_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_15_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload31 clknet_leaf_17_clk VGND VGND VPWR VPWR clkload31/Y sky130_fd_sc_hd__inv_12
Xclkload20 clknet_leaf_25_clk VGND VGND VPWR VPWR clkload20/Y sky130_fd_sc_hd__bufinv_16
X_2614_ clknet_leaf_26_clk _0163_ net144 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2545_ clknet_leaf_1_clk _0106_ net122 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_2476_ clknet_leaf_10_clk _0025_ net133 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1358_ gencon_inst.operand2\[8\] net54 _0676_ _0677_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__o22a_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1427_ net95 gencon_inst.mult_calc.adderSave\[6\] net371 net79 VGND VGND VPWR VPWR
+ _0177_ sky130_fd_sc_hd__a22o_1
X_1289_ gencon_inst.ALU_out\[11\] net69 net57 gencon_inst.mult_calc.out\[11\] _0565_
+ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__a221o_1
XFILLER_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload3 clknet_leaf_0_clk VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__inv_8
XFILLER_74_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2192_ gencon_inst.mult_calc.finish gencon_inst.ALU_finish VGND VGND VPWR VPWR _0394_
+ sky130_fd_sc_hd__or2_1
X_2330_ _1205_ _0477_ _0481_ net82 VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__a31o_1
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2261_ _1059_ _0448_ _0449_ _0450_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__or4_1
XFILLER_65_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1976_ input_ctrl_inst.debounce_cnt\[5\] input_ctrl_inst.debounce_cnt\[6\] input_ctrl_inst.debounce_cnt\[7\]
+ input_ctrl_inst.debounce_cnt\[8\] VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__o31a_1
X_2528_ clknet_leaf_39_clk _0089_ net120 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold15 gencon_inst.prev_operator_input\[0\] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 gencon_inst.mult_calc.INn1\[13\] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 gencon_inst.mult_calc.INn1\[15\] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 gencon_inst.mult_calc.diffSign VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ clknet_leaf_1_clk _0047_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[15\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold26 gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in1 VGND VGND VPWR VPWR
+ net186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_51_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1761_ gencon_inst.add_calc.main.GENERATE_ADDER\[1\].thingy.in1 _0944_ net110 VGND
+ VGND VPWR VPWR _0266_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1830_ net197 _0983_ net41 VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__mux2_1
XFILLER_30_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1692_ _0847_ _0898_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__xnor2_1
X_2313_ net419 net119 _1042_ _0480_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__a22o_1
XFILLER_65_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2175_ gencon_inst.gencon_state\[3\] _1215_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__nor2_2
X_2244_ net104 net343 net286 VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__o21ba_1
XFILLER_15_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1959_ gencon_inst.operator_input\[0\] VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput16 net16 VGND VGND VPWR VPWR display_output[14] sky130_fd_sc_hd__buf_2
Xoutput27 net27 VGND VGND VPWR VPWR input_state_FPGA[0] sky130_fd_sc_hd__buf_2
XFILLER_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_15_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1744_ gencon_inst.ALU_in1\[8\] gencon_inst.ALU_in2\[8\] net63 VGND VGND VPWR VPWR
+ _0936_ sky130_fd_sc_hd__mux2_1
X_2793_ clknet_leaf_6_clk _0337_ net134 VGND VGND VPWR VPWR gencon_inst.latched_operator_input\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1813_ gencon_inst.operand2\[7\] gencon_inst.operand1\[7\] net77 VGND VGND VPWR VPWR
+ _0975_ sky130_fd_sc_hd__mux2_1
XFILLER_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1675_ _0815_ _0816_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2089_ input_ctrl_inst.debounce_cnt\[6\] _1144_ net36 VGND VGND VPWR VPWR _1148_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_38_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2158_ input_ctrl_inst.RowSync\[2\] input_ctrl_inst.col_index\[3\] input_ctrl_inst.RowSync\[3\]
+ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2227_ _0402_ _0409_ _0411_ _0425_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1391_ net86 _1105_ net89 net242 VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__a2bb2o_1
X_1460_ net332 gencon_inst.mult_calc.INn2\[7\] net98 VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2012_ gencon_inst.mult_calc.count.GENERATE_ADDER\[9\].thingy.in1 gencon_inst.mult_calc.count.GENERATE_ADDER\[8\].thingy.in1
+ gencon_inst.mult_calc.count.GENERATE_ADDER\[7\].thingy.in1 _1077_ VGND VGND VPWR
+ VPWR _1079_ sky130_fd_sc_hd__and4_1
XFILLER_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold156 gencon_inst.add_calc.main.in2\[2\] VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__dlygate4sd3_1
X_1658_ _0838_ _0870_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__xor2_1
Xhold112 gencon_inst.ALU_in1\[1\] VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__dlygate4sd3_1
X_2776_ clknet_leaf_13_clk _0320_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[2\] sky130_fd_sc_hd__dfxtp_1
X_1727_ gencon_inst.ALU_in1\[15\] _0697_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__nand2_1
Xhold101 _0305_ VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold167 _0173_ VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in2 VGND VGND VPWR
+ VPWR net305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in2 VGND VGND VPWR
+ VPWR net294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 gencon_inst.mult_calc.count.GENERATE_ADDER\[14\].thingy.in1 VGND VGND VPWR
+ VPWR net283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 gencon_inst.add_calc.main.GENERATE_ADDER\[2\].thingy.in1 VGND VGND VPWR VPWR
+ net338 sky130_fd_sc_hd__dlygate4sd3_1
X_1589_ gencon_inst.add_calc.main.GENERATE_ADDER\[9\].thingy.in1 _0801_ _0802_ VGND
+ VGND VPWR VPWR _0804_ sky130_fd_sc_hd__nand3_1
Xhold189 gencon_inst.add_calc.main.in2\[12\] VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2561_ clknet_leaf_24_clk _0114_ net152 VGND VGND VPWR VPWR gencon_inst.operand1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2492_ clknet_leaf_6_clk _0057_ VGND VGND VPWR VPWR gencon_inst.keypad_input\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2630_ clknet_leaf_26_clk net306 net150 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
X_1512_ _0737_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__inv_2
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1374_ gencon_inst.operand2\[13\] gencon_inst.operand2\[12\] _0683_ VGND VGND VPWR
+ VPWR _0689_ sky130_fd_sc_hd__and3_1
X_1443_ net185 net172 net98 VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__mux2_1
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2828_ clknet_leaf_25_clk _0368_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2759_ clknet_leaf_13_clk _0303_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_73_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout62 net65 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_4
Xfanout40 _0998_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_52_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout73 _1210_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_2
Xfanout51 _0964_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_1_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout95 gencon_inst.mult_calc.state\[4\] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1992_ input_ctrl_inst.input_control_state\[0\] input_ctrl_inst.input_control_state\[1\]
+ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__nand2b_1
Xclkload10 clknet_leaf_39_clk VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_15_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload32 clknet_leaf_18_clk VGND VGND VPWR VPWR clkload32/Y sky130_fd_sc_hd__inv_12
X_2475_ clknet_leaf_9_clk _0024_ net133 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2613_ clknet_leaf_26_clk _0162_ net144 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload21 clknet_leaf_26_clk VGND VGND VPWR VPWR clkload21/Y sky130_fd_sc_hd__clkinv_2
X_2544_ clknet_leaf_1_clk _0105_ net121 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1288_ _0618_ _0619_ net72 VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__and3b_1
X_1357_ gencon_inst.mult_calc.out\[8\] net67 _0635_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__a21o_1
X_1426_ net94 net289 net320 net78 VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__a22o_1
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload4 clknet_leaf_1_clk VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__inv_6
XFILLER_59_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2191_ equal_input gencon_inst.read_input VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__nand2b_1
X_2260_ input_ctrl_inst.scan_timer\[1\] input_ctrl_inst.scan_timer\[0\] input_ctrl_inst.scan_timer\[15\]
+ input_ctrl_inst.scan_timer\[14\] VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_63_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1975_ _1046_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__inv_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold16 gencon_inst.mult_calc.INn1\[4\] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in1 VGND VGND VPWR VPWR
+ net187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in1 VGND VGND VPWR VPWR
+ net198 sky130_fd_sc_hd__dlygate4sd3_1
X_1409_ gencon_inst.mult_calc.out\[4\] net397 net104 VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__mux2_1
X_2458_ clknet_leaf_1_clk _0046_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_2527_ clknet_leaf_39_clk _0088_ net120 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold49 gencon_inst.mult_calc.INn1\[12\] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__dlygate4sd3_1
X_2389_ net403 _0519_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_26_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1760_ gencon_inst.ALU_in2\[1\] gencon_inst.ALU_in1\[1\] net62 VGND VGND VPWR VPWR
+ _0944_ sky130_fd_sc_hd__mux2_1
X_1691_ _0803_ _0804_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__and2b_1
X_2312_ gencon_inst.operator_input\[0\] net118 input_ctrl_inst.decoded_key\[2\] _0480_
+ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__a22o_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2174_ _1035_ _1214_ VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__nand2_1
X_2243_ net286 net343 VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__and2_1
Xoutput17 net17 VGND VGND VPWR VPWR display_output[15] sky130_fd_sc_hd__buf_2
X_1889_ net43 _0993_ _0994_ _0995_ net438 VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__o32a_1
X_1958_ gencon_inst.operand2\[8\] VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__inv_2
Xoutput28 net28 VGND VGND VPWR VPWR input_state_FPGA[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1743_ net290 _0935_ net112 VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__mux2_1
X_1674_ _0879_ _0881_ net31 VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__o21ai_1
X_2792_ clknet_leaf_6_clk _0336_ net134 VGND VGND VPWR VPWR gencon_inst.latched_operator_input\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1812_ net213 _0974_ net41 VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__mux2_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2226_ input_ctrl_inst.col_index\[4\] _0400_ _0401_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__or3_1
X_2088_ input_ctrl_inst.debounce_cnt\[6\] _1144_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__and2_1
XFILLER_53_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2157_ input_ctrl_inst.RowSync\[0\] input_ctrl_inst.col_index\[3\] input_ctrl_inst.RowSync\[1\]
+ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__or3b_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1390_ net86 _1103_ net88 net235 VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2011_ gencon_inst.mult_calc.count.GENERATE_ADDER\[7\].thingy.in1 _1077_ VGND VGND
+ VPWR VPWR _1078_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_33_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold168 gencon_inst.add_calc.main.in2\[8\] VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__dlygate4sd3_1
X_1588_ _0801_ _0802_ gencon_inst.add_calc.main.GENERATE_ADDER\[9\].thingy.in1 VGND
+ VGND VPWR VPWR _0803_ sky130_fd_sc_hd__a21oi_1
X_1657_ _0827_ _0828_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__nand2b_1
Xhold179 gencon_inst.add_calc.main.in2\[4\] VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__dlygate4sd3_1
X_1726_ net114 net347 net32 _0926_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__o22a_1
X_2775_ clknet_leaf_13_clk _0319_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[1\] sky130_fd_sc_hd__dfxtp_1
Xhold102 gencon_inst.addOrSub VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 _0179_ VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 input_ctrl_inst.col_index\[17\] VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 input_ctrl_inst.col_index\[6\] VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 gencon_inst.mult_calc.main.GENERATE_ADDER\[14\].thingy.in2 VGND VGND VPWR
+ VPWR net295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in2 VGND VGND VPWR
+ VPWR net273 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2209_ _0403_ _0404_ _0407_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__or3b_1
XFILLER_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_13_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2560_ clknet_leaf_24_clk _0113_ net152 VGND VGND VPWR VPWR gencon_inst.operand1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2491_ clknet_leaf_6_clk _0056_ VGND VGND VPWR VPWR gencon_inst.keypad_input\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1442_ net191 net176 net98 VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__mux2_1
X_1511_ gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in1
+ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__or2_1
XFILLER_67_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1373_ gencon_inst.operand2\[12\] _0688_ net55 VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__mux2_1
XFILLER_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2758_ clknet_leaf_13_clk _0302_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[0\] sky130_fd_sc_hd__dfxtp_1
X_2827_ clknet_leaf_25_clk _0367_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_1709_ net31 _0912_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__nand2_1
XFILLER_48_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2689_ clknet_leaf_5_clk _0233_ net128 VGND VGND VPWR VPWR gencon_inst.operand2\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_18_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout85 _1041_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_2
Xfanout63 net65 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_52_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout52 _0959_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_4
Xfanout74 _1210_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_2
Xfanout41 net42 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_4
Xfanout96 gencon_inst.mult_calc.state\[4\] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_63_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_72_Left_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload33 clknet_leaf_19_clk VGND VGND VPWR VPWR clkload33/Y sky130_fd_sc_hd__inv_12
XFILLER_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1991_ gencon_inst.key_read net82 _1059_ _1057_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__o211ai_1
Xclkload11 clknet_leaf_5_clk VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__clkinv_4
Xclkload22 clknet_leaf_27_clk VGND VGND VPWR VPWR clkload22/Y sky130_fd_sc_hd__bufinv_16
X_2612_ clknet_leaf_25_clk _0161_ net144 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2474_ clknet_leaf_9_clk _0023_ net133 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1425_ net95 gencon_inst.mult_calc.adderSave\[4\] net303 net78 VGND VGND VPWR VPWR
+ _0175_ sky130_fd_sc_hd__a22o_1
X_2543_ clknet_leaf_38_clk _0104_ net127 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1287_ gencon_inst.operand1\[10\] _0611_ gencon_inst.operand1\[11\] VGND VGND VPWR
+ VPWR _0619_ sky130_fd_sc_hd__a21o_1
X_1356_ _1030_ _0672_ _0675_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__a21oi_1
Xclkload5 clknet_leaf_2_clk VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__clkinv_4
XFILLER_11_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2190_ _1209_ net73 _0386_ _0391_ VGND VGND VPWR VPWR gencon_inst.next_state\[0\]
+ sky130_fd_sc_hd__or4_1
XFILLER_27_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1974_ input_ctrl_inst.debounce_cnt\[15\] input_ctrl_inst.debounce_cnt\[17\] input_ctrl_inst.debounce_cnt\[16\]
+ input_ctrl_inst.debounce_cnt\[18\] VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__and4_1
Xhold17 gencon_inst.mult_calc.INn1\[11\] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 gencon_inst.mult_calc.INn1\[3\] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 gencon_inst.mult_calc.INn2\[15\] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__dlygate4sd3_1
X_2457_ clknet_leaf_1_clk _0045_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_2526_ clknet_leaf_39_clk _0087_ net120 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_2388_ _0427_ _0508_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__nor2_1
X_1408_ gencon_inst.mult_calc.out\[3\] net387 net104 VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__mux2_1
XFILLER_56_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1339_ gencon_inst.operand2\[4\] net54 _0662_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__o21a_1
XFILLER_24_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1690_ _0892_ _0895_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__or2_1
XFILLER_51_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2311_ net118 _1187_ _1205_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__nor3_1
X_2242_ net102 _1126_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__and2_1
XFILLER_53_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2173_ gencon_inst.gencon_state\[1\] gencon_inst.gencon_state\[2\] VGND VGND VPWR
+ VPWR _1214_ sky130_fd_sc_hd__nor2_1
X_1957_ gencon_inst.operand2\[11\] VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__inv_2
XFILLER_21_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput18 net18 VGND VGND VPWR VPWR display_output[1] sky130_fd_sc_hd__buf_2
X_1888_ gencon_inst.operator_input\[0\] gencon_inst.key_read _0378_ _0383_ net44 VGND
+ VGND VPWR VPWR _0995_ sky130_fd_sc_hd__a41o_1
Xoutput29 net29 VGND VGND VPWR VPWR input_state_FPGA[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2509_ clknet_leaf_30_clk _0074_ net148 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[14\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_36_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_6_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2791_ clknet_leaf_6_clk _0335_ net134 VGND VGND VPWR VPWR gencon_inst.latched_operator_input\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1811_ gencon_inst.operand2\[6\] gencon_inst.operand1\[6\] net77 VGND VGND VPWR VPWR
+ _0974_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1742_ gencon_inst.ALU_in1\[7\] gencon_inst.ALU_in2\[7\] net63 VGND VGND VPWR VPWR
+ _0935_ sky130_fd_sc_hd__mux2_1
X_1673_ _0883_ _0882_ gencon_inst.ALU_out\[5\] _1041_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_7_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2225_ _0410_ _0419_ _0422_ _0423_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__or4b_1
Xclkbuf_leaf_18_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
X_2087_ net432 net38 net36 _1146_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__a22o_1
XFILLER_53_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2156_ _1197_ _1198_ input_ctrl_inst.RowSync\[1\] VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__o21bai_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2010_ gencon_inst.mult_calc.count.GENERATE_ADDER\[6\].thingy.in1 _1076_ VGND VGND
+ VPWR VPWR _1077_ sky130_fd_sc_hd__and2_1
XFILLER_75_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1725_ _1045_ gencon_inst.add_calc.sameSignVal net85 VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__a21o_1
X_2774_ clknet_leaf_13_clk _0318_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold158 gencon_inst.add_calc.main.in2\[9\] VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__dlygate4sd3_1
X_1587_ net108 gencon_inst.add_calc.main.in2\[9\] VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__nand2_1
X_1656_ _0864_ _0866_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__or2_1
Xhold103 _0297_ VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
Xhold147 gencon_inst.mult_calc.INn2\[14\] VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in2 VGND VGND VPWR
+ VPWR net329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 gencon_inst.mult_calc.adderSave\[13\] VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 _0184_ VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 _0185_ VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__dlygate4sd3_1
X_2139_ input_ctrl_inst.debounce_cnt\[18\] _1184_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__xnor2_1
XFILLER_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2208_ _0405_ _0406_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__nor2_1
XFILLER_41_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2490_ clknet_leaf_7_clk _0055_ VGND VGND VPWR VPWR gencon_inst.operator_input\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1441_ net198 net188 net98 VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__mux2_1
X_1510_ net440 net90 _0736_ net102 VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__a22o_1
XFILLER_67_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1372_ _0686_ _0687_ gencon_inst.mult_calc.out\[12\] net67 VGND VGND VPWR VPWR _0688_
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_18_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1708_ _0902_ _0905_ _0909_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__or3_1
X_2757_ clknet_leaf_9_clk _0301_ VGND VGND VPWR VPWR gencon_inst.add_calc.start sky130_fd_sc_hd__dfxtp_1
X_2826_ clknet_leaf_25_clk _0366_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2688_ clknet_leaf_31_clk _0004_ net142 VGND VGND VPWR VPWR gencon_inst.mult_calc.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1639_ _0791_ _0795_ _0851_ _0792_ _0788_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__o311a_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout31 net32 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
Xfanout64 net65 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_52_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout53 _0959_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_2
Xfanout42 _0967_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
Xfanout97 gencon_inst.mult_calc.state\[4\] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout86 _1040_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1990_ net92 input_ctrl_inst.input_control_state\[1\] input_ctrl_inst.input_control_state\[0\]
+ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__nand3b_1
XTAP_TAPCELL_ROW_15_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload34 clknet_leaf_20_clk VGND VGND VPWR VPWR clkload34/Y sky130_fd_sc_hd__inv_12
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload12 clknet_leaf_7_clk VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__inv_8
Xclkload23 clknet_leaf_28_clk VGND VGND VPWR VPWR clkload23/Y sky130_fd_sc_hd__inv_8
X_2542_ clknet_leaf_36_clk _0103_ net127 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_2611_ clknet_leaf_33_clk _0160_ net139 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_2473_ clknet_leaf_9_clk _0022_ net133 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1355_ _1211_ _0674_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__or2_1
X_1424_ net95 gencon_inst.mult_calc.adderSave\[3\] net323 net79 VGND VGND VPWR VPWR
+ _0174_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1286_ gencon_inst.operand1\[10\] gencon_inst.operand1\[11\] _0611_ VGND VGND VPWR
+ VPWR _0618_ sky130_fd_sc_hd__and3_1
Xclkload6 clknet_leaf_3_clk VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__inv_6
XFILLER_59_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2809_ clknet_leaf_23_clk _0353_ net156 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dfrtp_1
XFILLER_3_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1973_ net106 VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__inv_2
X_2525_ clknet_leaf_39_clk _0086_ net120 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1338_ gencon_inst.mult_calc.out\[4\] net66 _0660_ _0661_ VGND VGND VPWR VPWR _0662_
+ sky130_fd_sc_hd__a22o_1
Xhold18 gencon_inst.mult_calc.INn1\[8\] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in1 VGND VGND VPWR
+ VPWR net189 sky130_fd_sc_hd__dlygate4sd3_1
X_1407_ gencon_inst.mult_calc.out\[2\] net390 net104 VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__mux2_1
XFILLER_29_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2387_ _0518_ _0519_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__nor2_1
X_2456_ clknet_leaf_1_clk _0044_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1269_ gencon_inst.ALU_out\[7\] net70 net57 gencon_inst.mult_calc.out\[7\] net43
+ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__a221o_1
XFILLER_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2241_ net277 net321 net246 VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__o21ba_1
X_2172_ gencon_inst.mult_calc.finish _1212_ VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__and2_1
X_2310_ net125 _1187_ _0478_ _0479_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__a211oi_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1887_ net93 gencon_inst.mult_calc.out\[15\] _1214_ net68 gencon_inst.ALU_out\[15\]
+ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_31_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1956_ net119 net286 net41 VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__a21o_1
Xoutput19 net19 VGND VGND VPWR VPWR display_output[2] sky130_fd_sc_hd__buf_2
X_2508_ clknet_leaf_30_clk net234 net148 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[13\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2439_ _0554_ _0555_ _0553_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__o21ai_1
XFILLER_72_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1741_ net420 _0934_ net112 VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__mux2_1
X_2790_ clknet_leaf_4_clk _0334_ VGND VGND VPWR VPWR gencon_inst.prev_read_input sky130_fd_sc_hd__dfxtp_1
X_1810_ net172 _0973_ net41 VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__mux2_1
X_1672_ net31 _0879_ _0881_ net85 VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__a31o_1
X_2155_ input_ctrl_inst.col_index\[2\] input_ctrl_inst.col_index\[3\] VGND VGND VPWR
+ VPWR _1198_ sky130_fd_sc_hd__and2_1
X_2224_ input_ctrl_inst.col_index\[13\] input_ctrl_inst.col_index\[12\] input_ctrl_inst.col_index\[15\]
+ input_ctrl_inst.col_index\[14\] VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__and4_1
X_2086_ _1144_ _1145_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__nor2_1
XFILLER_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1939_ net52 _0983_ net40 net408 _1028_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__a221o_1
XFILLER_67_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1724_ net439 _0925_ net115 VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__mux2_1
X_2773_ clknet_leaf_14_clk _0317_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[15\] sky130_fd_sc_hd__dfxtp_1
Xhold115 input_ctrl_inst.debounce_cnt\[3\] VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_41_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold126 gencon_inst.mult_calc.start VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold104 gencon_inst.mult_calc.countSave\[9\] VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__dlygate4sd3_1
X_1586_ net108 gencon_inst.add_calc.main.in2\[9\] VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__or2_1
X_1655_ _0868_ _0867_ net436 net85 VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__a2bb2o_1
Xhold148 gencon_inst.mult_calc.INn2\[2\] VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 gencon_inst.mult_calc.INn2\[6\] VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 gencon_inst.mult_calc.count.GENERATE_ADDER\[11\].thingy.in1 VGND VGND VPWR
+ VPWR net297 sky130_fd_sc_hd__dlygate4sd3_1
X_2138_ _1183_ _1184_ _1185_ net37 net431 VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__a32o_1
X_2069_ _1054_ net30 _1131_ _1053_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__a22o_1
XFILLER_26_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2207_ input_ctrl_inst.col_index\[21\] input_ctrl_inst.col_index\[20\] input_ctrl_inst.col_index\[23\]
+ input_ctrl_inst.col_index\[22\] VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__or4_1
XFILLER_64_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1371_ gencon_inst.operand2\[12\] _0683_ net74 VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__o21ai_1
X_1440_ net182 net171 net99 VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__mux2_1
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2825_ clknet_leaf_25_clk _0365_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1707_ _0911_ _0910_ gencon_inst.ALU_out\[11\] net85 VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__a2bb2o_1
X_1638_ _0791_ _0795_ _0851_ _0792_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__o31a_1
X_2756_ clknet_leaf_5_clk _0300_ VGND VGND VPWR VPWR gencon_inst.prev_operator_input\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2687_ clknet_leaf_36_clk _0003_ net127 VGND VGND VPWR VPWR gencon_inst.mult_calc.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1569_ _0782_ _0783_ gencon_inst.add_calc.main.GENERATE_ADDER\[14\].thingy.in1 VGND
+ VGND VPWR VPWR _0784_ sky130_fd_sc_hd__a21oi_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout32 _0858_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
Xfanout65 _0927_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_52_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout43 _0565_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_4
Xfanout76 _0388_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_4
Xfanout54 _0636_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout98 net99 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_4
Xfanout87 _1040_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_9_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload35 clknet_leaf_21_clk VGND VGND VPWR VPWR clkload35/Y sky130_fd_sc_hd__clkinv_8
X_2472_ clknet_leaf_9_clk _0021_ net133 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload13 clknet_leaf_8_clk VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__inv_6
X_2610_ clknet_leaf_35_clk _0159_ net143 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2541_ clknet_leaf_38_clk _0102_ net121 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload24 clknet_leaf_29_clk VGND VGND VPWR VPWR clkload24/Y sky130_fd_sc_hd__inv_8
X_1285_ gencon_inst.operand1\[10\] net45 _0616_ _0617_ VGND VGND VPWR VPWR _0117_
+ sky130_fd_sc_hd__o22a_1
X_1354_ gencon_inst.operand2\[8\] gencon_inst.operand2\[7\] _0667_ VGND VGND VPWR
+ VPWR _0674_ sky130_fd_sc_hd__and3_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1423_ net95 gencon_inst.mult_calc.adderSave\[2\] net326 net79 VGND VGND VPWR VPWR
+ _0173_ sky130_fd_sc_hd__a22o_1
XFILLER_70_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2808_ clknet_leaf_22_clk _0352_ net156 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dfrtp_1
Xclkload7 clknet_leaf_4_clk VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__inv_6
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2739_ clknet_leaf_35_clk _0283_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1972_ input_ctrl_inst.col_index\[24\] VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2455_ clknet_leaf_4_clk _0043_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_2524_ clknet_leaf_39_clk _0085_ net120 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1268_ _0602_ _0603_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__nor2_1
X_1337_ gencon_inst.operand2\[4\] _0658_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__or2_1
Xhold19 gencon_inst.mult_calc.INn1\[9\] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__dlygate4sd3_1
X_1406_ gencon_inst.mult_calc.out\[1\] net291 net104 VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__mux2_1
XFILLER_28_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2386_ input_ctrl_inst.col_index\[13\] input_ctrl_inst.col_index\[12\] input_ctrl_inst.col_index\[14\]
+ _0515_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__and4_1
XFILLER_24_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_69_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2240_ net246 net321 VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__and2_1
X_2171_ gencon_inst.gencon_state\[1\] _1035_ _1036_ gencon_inst.gencon_state\[2\]
+ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__and4b_1
XFILLER_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1886_ gencon_inst.operand1\[15\] _0630_ _0992_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__o21a_1
X_1955_ gencon_inst.operand2\[15\] net51 net34 net199 VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_31_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2507_ clknet_leaf_30_clk _0072_ net148 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[12\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2438_ input_ctrl_inst.col_index\[30\] _0551_ _0528_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_39_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2369_ net58 _0508_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__nor2_1
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_75 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1671_ net31 _0879_ _0881_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__a21oi_1
X_1740_ gencon_inst.ALU_in1\[6\] gencon_inst.ALU_in2\[6\] net65 VGND VGND VPWR VPWR
+ _0934_ sky130_fd_sc_hd__mux2_1
XFILLER_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2085_ input_ctrl_inst.debounce_cnt\[4\] _1139_ input_ctrl_inst.debounce_cnt\[5\]
+ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_36_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2154_ input_ctrl_inst.col_index\[2\] input_ctrl_inst.col_index\[3\] VGND VGND VPWR
+ VPWR _1197_ sky130_fd_sc_hd__nor2_1
X_2223_ input_ctrl_inst.col_index\[9\] input_ctrl_inst.col_index\[8\] input_ctrl_inst.col_index\[11\]
+ input_ctrl_inst.col_index\[10\] VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_44_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1869_ gencon_inst.operand1\[13\] net229 net48 VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__mux2_1
X_1938_ _0387_ _0560_ _0994_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__o21a_1
XFILLER_67_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1654_ net32 _0864_ _0866_ net85 VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__a31o_1
X_1723_ _0922_ _0924_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__xnor2_1
Xhold149 gencon_inst.add_calc.sameSignVal VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__dlygate4sd3_1
X_2772_ clknet_leaf_16_clk _0316_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold105 gencon_inst.mult_calc.INn2\[3\] VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 gencon_inst.mult_calc.INn2\[9\] VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in2 VGND VGND VPWR
+ VPWR net287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 gencon_inst.mult_calc.countSave\[11\] VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__dlygate4sd3_1
X_1585_ gencon_inst.add_calc.main.GENERATE_ADDER\[10\].thingy.in1 _0797_ _0798_ VGND
+ VGND VPWR VPWR _0800_ sky130_fd_sc_hd__nand3_1
X_2206_ input_ctrl_inst.col_index\[17\] input_ctrl_inst.col_index\[16\] input_ctrl_inst.col_index\[19\]
+ input_ctrl_inst.col_index\[18\] VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__or4_1
X_2137_ input_ctrl_inst.debounce_cnt\[17\] _1053_ _1132_ net36 VGND VGND VPWR VPWR
+ _1185_ sky130_fd_sc_hd__a31o_1
X_2068_ _1051_ _1055_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__nor2_2
XFILLER_34_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1370_ gencon_inst.operand2\[12\] _0683_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__and2_1
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2824_ clknet_leaf_35_clk _0364_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1706_ net31 _0907_ _0909_ _1041_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__a31o_1
X_1637_ _0795_ _0851_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__nor2_1
X_2755_ clknet_leaf_4_clk _0299_ VGND VGND VPWR VPWR gencon_inst.prev_operator_input\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2686_ clknet_leaf_33_clk _0007_ net142 VGND VGND VPWR VPWR gencon_inst.mult_calc.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1568_ net107 gencon_inst.add_calc.main.in2\[14\] VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__nand2_1
X_1499_ _0724_ _0726_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__nand2_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout44 _0564_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_4
Xfanout55 _0636_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
Xfanout33 net34 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_2
Xfanout77 _0388_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_2
Xfanout66 _0634_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_2
XFILLER_13_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout88 net91 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_2
Xfanout99 gencon_inst.mult_calc.state\[3\] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_4
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_41_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload14 clknet_leaf_9_clk VGND VGND VPWR VPWR clkload14/Y sky130_fd_sc_hd__inv_6
X_2471_ clknet_leaf_9_clk _0020_ net132 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload36 clknet_leaf_22_clk VGND VGND VPWR VPWR clkload36/Y sky130_fd_sc_hd__clkinv_4
X_1422_ net95 net291 net412 net79 VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__a22o_1
Xclkload25 clknet_leaf_30_clk VGND VGND VPWR VPWR clkload25/Y sky130_fd_sc_hd__clkinv_8
X_2540_ clknet_leaf_36_clk _0101_ net127 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_1284_ gencon_inst.ALU_out\[10\] net69 net57 gencon_inst.mult_calc.out\[10\] net43
+ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_50_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1353_ gencon_inst.operand2\[7\] _0673_ net54 VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2807_ clknet_leaf_23_clk _0351_ net151 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dfrtp_1
X_2738_ clknet_leaf_36_clk _0282_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload8 clknet_leaf_37_clk VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__inv_6
X_2669_ clknet_leaf_36_clk _0218_ net129 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1971_ net450 VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__inv_2
XFILLER_68_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1405_ gencon_inst.mult_calc.out\[0\] net395 net104 VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__mux2_1
X_2454_ clknet_leaf_36_clk _0042_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_2385_ input_ctrl_inst.col_index\[13\] _0517_ net425 VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__a21oi_1
X_2523_ clknet_leaf_0_clk _0084_ net120 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1267_ gencon_inst.operand1\[7\] _0598_ net72 VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__o21ai_1
X_1336_ _1211_ _0659_ net54 VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__o21ai_1
Xinput1 RowIn[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_24_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_39_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2170_ gencon_inst.gencon_state\[1\] _1035_ gencon_inst.gencon_state\[3\] _1037_
+ VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__or4_2
XFILLER_25_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1954_ gencon_inst.operand2\[14\] net51 net33 net307 VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__a22o_1
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1885_ gencon_inst.operand1\[15\] _0630_ _0559_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__a21oi_1
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2506_ clknet_leaf_30_clk _0071_ net146 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[11\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2368_ _0421_ _0502_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__nand2_1
X_2437_ input_ctrl_inst.col_index\[30\] _0551_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__nor2_1
XFILLER_56_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1319_ gencon_inst.operand2\[1\] _0645_ net54 VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__mux2_1
X_2299_ net245 _0471_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__xor2_1
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1670_ _0841_ _0880_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__xnor2_2
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2222_ input_ctrl_inst.col_index\[4\] _0398_ _0420_ _0419_ VGND VGND VPWR VPWR _0421_
+ sky130_fd_sc_hd__a31o_1
X_2084_ input_ctrl_inst.debounce_cnt\[4\] input_ctrl_inst.debounce_cnt\[5\] _1139_
+ VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_36_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2153_ input_ctrl_inst.decoded_key\[2\] net82 _1187_ _1196_ VGND VGND VPWR VPWR _0029_
+ sky130_fd_sc_hd__a211o_1
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1937_ _1027_ net226 net39 VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1868_ gencon_inst.operand1\[12\] net230 net48 VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__mux2_1
X_1799_ gencon_inst.operand2\[0\] gencon_inst.operand1\[0\] net76 VGND VGND VPWR VPWR
+ _0968_ sky130_fd_sc_hd__mux2_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2771_ clknet_leaf_24_clk _0315_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2840_ clknet_leaf_36_clk _0377_ VGND VGND VPWR VPWR gencon_inst.mult_calc.start
+ sky130_fd_sc_hd__dfxtp_1
X_1584_ _0797_ _0798_ gencon_inst.add_calc.main.GENERATE_ADDER\[10\].thingy.in1 VGND
+ VGND VPWR VPWR _0799_ sky130_fd_sc_hd__a21oi_1
X_1653_ net32 _0864_ _0866_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__a21oi_1
X_1722_ _0855_ _0923_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__xnor2_1
Xhold117 gencon_inst.add_calc.next_finish VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 gencon_inst.keypad_input\[0\] VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold106 net25 VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 _0183_ VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2205_ net117 input_ctrl_inst.col_index\[1\] net116 input_ctrl_inst.col_index\[3\]
+ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__o31a_1
X_2136_ input_ctrl_inst.debounce_cnt\[17\] _1180_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__nand2_1
X_2067_ _1051_ net30 _1064_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__o21ai_1
XFILLER_22_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1705_ net32 _0907_ _0909_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__a21oi_1
X_2754_ clknet_leaf_5_clk _0298_ VGND VGND VPWR VPWR gencon_inst.prev_operator_input\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2823_ clknet_leaf_5_clk _0363_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1636_ _0799_ _0803_ _0848_ _0800_ _0796_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__o311a_1
X_1567_ net107 gencon_inst.add_calc.main.in2\[14\] VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__or2_1
X_2685_ clknet_leaf_33_clk _0006_ net142 VGND VGND VPWR VPWR gencon_inst.mult_calc.next_finish
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2119_ input_ctrl_inst.debounce_cnt\[12\] input_ctrl_inst.debounce_cnt\[13\] _1160_
+ input_ctrl_inst.debounce_cnt\[14\] VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__a31o_1
X_1498_ gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in1
+ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout45 _0564_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
Xfanout56 _0563_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
Xfanout67 _0634_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_2
Xfanout34 _0966_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
Xfanout78 _1068_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_4
Xfanout89 net91 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
XFILLER_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload15 clknet_leaf_10_clk VGND VGND VPWR VPWR clkload15/Y sky130_fd_sc_hd__clkinv_8
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload26 clknet_leaf_31_clk VGND VGND VPWR VPWR clkload26/Y sky130_fd_sc_hd__clkinv_2
X_2470_ clknet_leaf_8_clk _0019_ net132 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload37 clknet_leaf_23_clk VGND VGND VPWR VPWR clkload37/Y sky130_fd_sc_hd__clkinv_8
X_1421_ net95 net395 net407 net79 VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1283_ gencon_inst.operand1\[10\] _0611_ _0615_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__a21oi_1
X_1352_ net74 _0671_ _0672_ net67 gencon_inst.mult_calc.out\[7\] VGND VGND VPWR VPWR
+ _0673_ sky130_fd_sc_hd__a32o_1
XFILLER_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2806_ clknet_leaf_22_clk _0350_ net156 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dfrtp_1
X_2737_ clknet_leaf_36_clk _0281_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload9 clknet_leaf_38_clk VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__clkinv_8
X_2668_ clknet_leaf_36_clk _0217_ net130 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1619_ gencon_inst.add_calc.main.GENERATE_ADDER\[1\].thingy.in1 _0833_ VGND VGND
+ VPWR VPWR _0834_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_6_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2599_ clknet_leaf_31_clk _0148_ net146 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1970_ input_ctrl_inst.decoded_key\[3\] VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_23_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2522_ clknet_leaf_0_clk _0083_ net120 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1335_ gencon_inst.operand2\[4\] _0658_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__and2_1
X_1404_ net208 _0699_ net99 VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__mux2_1
X_2453_ clknet_leaf_36_clk _0041_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_2384_ net383 _0517_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__xor2_1
XFILLER_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1266_ gencon_inst.operand1\[7\] _0598_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__and2_1
XFILLER_28_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput2 RowIn[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1884_ net165 _0961_ _0991_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__o21ai_1
X_1953_ gencon_inst.operand2\[13\] net50 net34 net342 VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__a22o_1
XFILLER_33_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2505_ clknet_leaf_31_clk _0070_ net146 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[10\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1318_ net73 _0643_ _0644_ net66 gencon_inst.mult_calc.out\[1\] VGND VGND VPWR VPWR
+ _0645_ sky130_fd_sc_hd__a32o_1
X_2298_ _0471_ _0472_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__nor2_1
X_2367_ input_ctrl_inst.col_index\[6\] _0506_ net402 VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__a21oi_1
X_2436_ input_ctrl_inst.col_index\[30\] net58 VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__nand2_1
XFILLER_72_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1249_ gencon_inst.ALU_out\[3\] net71 net56 gencon_inst.mult_calc.out\[3\] net43
+ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_39_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap75 _0397_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_1
X_2152_ net82 _1195_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__nor2_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2221_ input_ctrl_inst.col_index\[5\] input_ctrl_inst.col_index\[7\] input_ctrl_inst.col_index\[6\]
+ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__and3_1
X_2083_ net35 _1142_ _1143_ net38 net410 VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__a32o_1
X_1867_ gencon_inst.operand1\[11\] net203 net48 VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__mux2_1
X_1936_ gencon_inst.ALU_out\[14\] net69 net60 gencon_inst.mult_calc.out\[14\] _1026_
+ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_44_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1798_ gencon_inst.read_input net128 net52 net51 VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_10_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2419_ net418 net58 _0528_ _0541_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__a22o_1
XFILLER_8_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1721_ _0784_ _0856_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__nor2_1
X_2770_ clknet_leaf_22_clk _0314_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1652_ _0837_ _0865_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__xnor2_1
X_1583_ net108 gencon_inst.add_calc.main.in2\[10\] VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__nand2_1
Xhold129 gencon_inst.mult_calc.adderSave\[5\] VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold107 gencon_inst.mult_calc.compCount.in2\[0\] VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in1 VGND VGND VPWR
+ VPWR net278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2135_ input_ctrl_inst.debounce_cnt\[17\] _1180_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__or2_1
X_2204_ _0399_ _0400_ _0401_ net75 VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__o31a_1
X_2066_ _1054_ _1128_ _1130_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__a21bo_1
X_1919_ net266 net39 _1014_ _1015_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__a211o_1
XFILLER_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1704_ _0850_ _0908_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__xnor2_1
X_2753_ clknet_leaf_14_clk net263 VGND VGND VPWR VPWR gencon_inst.addOrSub sky130_fd_sc_hd__dfxtp_1
X_2822_ clknet_leaf_5_clk net240 VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2684_ clknet_leaf_36_clk _0002_ net127 VGND VGND VPWR VPWR gencon_inst.mult_calc.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_1635_ _0799_ _0803_ _0848_ _0800_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__o31a_1
X_1566_ net430 _0781_ net114 VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__mux2_1
X_1497_ _0724_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2118_ input_ctrl_inst.debounce_cnt\[14\] _1064_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_1_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2049_ _1115_ _1113_ gencon_inst.mult_calc.compCount.in2\[10\] _1114_ VGND VGND VPWR
+ VPWR _1116_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout35 net36 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_2
Xfanout46 _0984_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_4
Xfanout57 _0563_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_2
Xfanout68 net71 VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_2
Xfanout79 _1068_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload16 clknet_leaf_11_clk VGND VGND VPWR VPWR clkload16/Y sky130_fd_sc_hd__inv_8
Xclkload38 clknet_leaf_24_clk VGND VGND VPWR VPWR clkload38/Y sky130_fd_sc_hd__clkinv_8
Xclkload27 clknet_leaf_32_clk VGND VGND VPWR VPWR clkload27/Y sky130_fd_sc_hd__inv_6
X_1351_ gencon_inst.operand2\[7\] _0667_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__nand2_1
X_1420_ net253 net208 net104 VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__mux2_1
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1282_ gencon_inst.operand1\[10\] _0611_ net72 VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__o21ai_1
XFILLER_51_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2805_ clknet_leaf_23_clk _0349_ net156 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1618_ gencon_inst.add_calc.main.in2\[1\] net106 VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__xor2_1
X_2736_ clknet_leaf_11_clk _0280_ net136 VGND VGND VPWR VPWR gencon_inst.ALU_finish
+ sky130_fd_sc_hd__dfrtp_1
X_2667_ clknet_leaf_31_clk _0216_ net147 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1549_ net102 _0768_ _0769_ net301 net90 VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_6_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2598_ clknet_leaf_31_clk _0147_ net146 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold290 input_ctrl_inst.read_input_flag VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2521_ clknet_leaf_0_clk _0082_ net122 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1265_ gencon_inst.operand1\[6\] net44 _0600_ _0601_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__o22a_1
XFILLER_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1334_ _0652_ _0654_ _0653_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__o21bai_1
X_1403_ gencon_inst.mult_calc.INn2\[15\] gencon_inst.mult_calc.INn1\[15\] VGND VGND
+ VPWR VPWR _0699_ sky130_fd_sc_hd__xor2_1
X_2452_ clknet_leaf_4_clk _0040_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2383_ _0516_ _0517_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 RowIn[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
X_2719_ clknet_leaf_19_clk _0263_ net158 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1883_ net93 _1207_ _0960_ _0990_ _0989_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__o221a_1
X_1952_ gencon_inst.operand2\[12\] net50 net33 net374 VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__a22o_1
XFILLER_33_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2504_ clknet_leaf_31_clk _0069_ net146 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[9\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2435_ _0527_ _0552_ net441 net58 VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__a2bb2o_1
X_1248_ _0586_ _0587_ net72 VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_39_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1317_ _0638_ _0641_ _0642_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__or3_1
X_2297_ net389 _0469_ _0445_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__o21ai_1
X_2366_ net317 _0506_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__xor2_1
XFILLER_64_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Left_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_65_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_74_Left_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2082_ input_ctrl_inst.debounce_cnt\[4\] _1139_ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__or2_1
X_2151_ net116 _1194_ _1193_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__mux2_1
X_2220_ _0399_ _0404_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__nor2_1
XFILLER_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1866_ gencon_inst.operand1\[10\] net348 net48 VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__mux2_1
X_1935_ _0561_ _0982_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_44_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1797_ net119 _0961_ _0965_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__o21a_1
X_2418_ _0539_ _0540_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__nor2_1
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2349_ net117 _0444_ input_ctrl_inst.col_index\[1\] VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__a21oi_1
XFILLER_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1651_ _0831_ _0832_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__nand2b_1
X_1720_ _0912_ _0915_ _0919_ net31 VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__o31a_1
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold108 _0202_ VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__dlygate4sd3_1
X_1582_ net108 gencon_inst.add_calc.main.in2\[10\] VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__or2_1
Xhold119 gencon_inst.mult_calc.adderSave\[7\] VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2134_ _1179_ _1181_ _1182_ net37 net426 VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__a32o_1
X_2065_ _1051_ _1065_ _1128_ _1129_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_49_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2203_ _0400_ _0401_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__nor2_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1849_ gencon_inst.operand2\[9\] net421 net48 VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__mux2_1
X_1918_ gencon_inst.operand1\[8\] _0378_ net77 VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__and3_1
XFILLER_57_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_20_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2821_ clknet_leaf_35_clk net345 VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1634_ _0803_ _0848_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__nor2_1
X_1703_ _0795_ _0796_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_11_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
X_2683_ clknet_leaf_13_clk _0232_ net136 VGND VGND VPWR VPWR gencon_inst.add_calc.diffSign
+ sky130_fd_sc_hd__dfrtp_1
X_2752_ clknet_leaf_4_clk _0296_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_1565_ gencon_inst.add_calc.main.a0.in1 gencon_inst.add_calc.main.in2\[0\] VGND VGND
+ VPWR VPWR _0781_ sky130_fd_sc_hd__xor2_1
X_1496_ gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in1
+ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__or2_1
X_2117_ input_ctrl_inst.debounce_cnt\[13\] net37 _1166_ _1168_ VGND VGND VPWR VPWR
+ _0012_ sky130_fd_sc_hd__a22o_1
XFILLER_39_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2048_ gencon_inst.mult_calc.compCount.in2\[9\] _1111_ _1114_ gencon_inst.mult_calc.compCount.in2\[10\]
+ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__a22oi_1
Xfanout47 _0984_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
Xfanout36 _1134_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_2
Xfanout69 net70 VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_2
XFILLER_13_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout58 net59 VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_2
XFILLER_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload17 clknet_leaf_12_clk VGND VGND VPWR VPWR clkload17/Y sky130_fd_sc_hd__inv_8
Xclkload28 clknet_leaf_33_clk VGND VGND VPWR VPWR clkload28/Y sky130_fd_sc_hd__inv_6
XFILLER_68_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1281_ gencon_inst.operand1\[9\] net45 _0613_ _0614_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__o22a_1
X_1350_ gencon_inst.operand2\[7\] _0667_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__or2_1
XFILLER_63_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
X_2804_ clknet_leaf_16_clk _0348_ net152 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1617_ gencon_inst.add_calc.main.GENERATE_ADDER\[2\].thingy.in1 _0829_ _0830_ VGND
+ VGND VPWR VPWR _0832_ sky130_fd_sc_hd__nand3_1
X_2735_ clknet_leaf_16_clk _0279_ net154 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[14\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2597_ clknet_leaf_31_clk _0146_ net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2666_ clknet_leaf_31_clk _0215_ net147 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1479_ gencon_inst.mult_calc.main.a0.in2 gencon_inst.mult_calc.main.a0.in1 gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in2
+ gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in1 VGND VGND VPWR VPWR _0710_
+ sky130_fd_sc_hd__a22oi_1
X_1548_ _0765_ _0766_ _0767_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_65_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold280 gencon_inst.mult_calc.adderSave\[6\] VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1402_ gencon_inst.ALU_in1\[15\] net309 _0698_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__mux2_1
X_2451_ clknet_leaf_36_clk _0039_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2520_ clknet_leaf_0_clk _0081_ net122 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1264_ gencon_inst.ALU_out\[6\] net70 net56 gencon_inst.mult_calc.out\[6\] net43
+ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__a221o_1
X_1333_ gencon_inst.operand2\[3\] _0657_ net54 VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__mux2_1
XFILLER_36_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 RowIn[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_2382_ input_ctrl_inst.col_index\[11\] input_ctrl_inst.col_index\[12\] _0513_ VGND
+ VGND VPWR VPWR _0517_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_62_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2718_ clknet_leaf_21_clk _0262_ net159 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_2649_ clknet_leaf_27_clk _0198_ net151 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1882_ _1031_ _0383_ gencon_inst.prev_operator_input\[2\] gencon_inst.prev_operator_input\[0\]
+ gencon_inst.prev_operator_input\[1\] VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__a2111o_1
X_1951_ gencon_inst.operand2\[11\] net50 net33 net359 VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__a22o_1
X_2503_ clknet_leaf_31_clk net255 net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[8\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2365_ _0505_ _0506_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__nor2_1
X_2434_ _0550_ _0551_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__or2_1
X_1247_ _0584_ _0585_ _0577_ _0580_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_39_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1316_ _0641_ _0642_ _0638_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__o21ai_1
X_2296_ input_ctrl_inst.scan_timer\[15\] _0469_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__and2_1
XFILLER_64_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2081_ input_ctrl_inst.debounce_cnt\[4\] _1139_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__nand2_1
XFILLER_38_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2150_ input_ctrl_inst.RowSync\[2\] input_ctrl_inst.RowSync\[0\] net116 VGND VGND
+ VPWR VPWR _1194_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1934_ _1024_ _1025_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__or2_1
X_1865_ gencon_inst.operand1\[9\] net386 net48 VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__mux2_1
X_1796_ net51 VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__inv_2
XFILLER_69_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2348_ net117 net59 VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__xnor2_1
X_2417_ _1044_ _0429_ _0508_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__nor3_2
X_2279_ input_ctrl_inst.scan_timer\[7\] input_ctrl_inst.scan_timer\[8\] _0458_ VGND
+ VGND VPWR VPWR _0461_ sky130_fd_sc_hd__and3_1
XFILLER_16_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1650_ _0781_ _0860_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__nand2b_1
X_1581_ gencon_inst.add_calc.main.GENERATE_ADDER\[11\].thingy.in1 _0793_ _0794_ VGND
+ VGND VPWR VPWR _0796_ sky130_fd_sc_hd__nand3_1
Xhold109 gencon_inst.mult_calc.countSave\[10\] VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__dlygate4sd3_1
X_2202_ input_ctrl_inst.col_index\[9\] input_ctrl_inst.col_index\[8\] input_ctrl_inst.col_index\[11\]
+ input_ctrl_inst.col_index\[10\] VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__or4_1
XFILLER_66_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2133_ input_ctrl_inst.debounce_cnt\[16\] _1053_ _1132_ net36 VGND VGND VPWR VPWR
+ _1182_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_49_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2064_ _1032_ _1052_ _1064_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__or3_1
X_1917_ gencon_inst.operand2\[8\] _0387_ net61 gencon_inst.mult_calc.out\[8\] _0609_
+ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__a221o_1
X_1779_ net356 _0953_ net113 VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__mux2_1
X_1848_ gencon_inst.operand2\[8\] net416 net49 VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__mux2_1
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2820_ clknet_leaf_6_clk gencon_inst.next_state\[3\] net134 VGND VGND VPWR VPWR gencon_inst.gencon_state\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_31_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2751_ clknet_leaf_34_clk _0295_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_1633_ _0807_ _0811_ _0845_ _0808_ _0804_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__o311a_1
XFILLER_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1702_ _0902_ _0905_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__or2_1
X_1564_ gencon_inst.operand2\[15\] _0780_ _0779_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__o21a_1
X_2682_ clknet_leaf_29_clk _0231_ net147 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1495_ net397 net88 _0723_ net103 VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__a22o_1
X_2116_ input_ctrl_inst.debounce_cnt\[13\] _1163_ _1167_ net35 VGND VGND VPWR VPWR
+ _1168_ sky130_fd_sc_hd__o2bb2a_1
Xfanout37 _1133_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
XFILLER_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2047_ gencon_inst.mult_calc.count.GENERATE_ADDER\[10\].thingy.in1 _1079_ VGND VGND
+ VPWR VPWR _1114_ sky130_fd_sc_hd__xnor2_1
Xfanout48 net49 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_4
Xfanout59 _0443_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_17_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload18 clknet_leaf_13_clk VGND VGND VPWR VPWR clkload18/Y sky130_fd_sc_hd__inv_4
Xclkload29 clknet_leaf_34_clk VGND VGND VPWR VPWR clkload29/Y sky130_fd_sc_hd__clkinv_8
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1280_ gencon_inst.ALU_out\[9\] net69 net57 gencon_inst.mult_calc.out\[9\] net43
+ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__a221o_1
XFILLER_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2734_ clknet_leaf_19_clk _0278_ net158 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[13\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2803_ clknet_leaf_14_clk _0347_ net152 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfrtp_1
X_1616_ _0829_ _0830_ gencon_inst.add_calc.main.GENERATE_ADDER\[2\].thingy.in1 VGND
+ VGND VPWR VPWR _0831_ sky130_fd_sc_hd__a21oi_1
X_1547_ _0765_ _0766_ _0767_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__nand3_1
X_2596_ clknet_leaf_32_clk _0145_ net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2665_ clknet_leaf_29_clk _0214_ net148 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1478_ _0707_ _0708_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_65_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold270 gencon_inst.ALU_out\[0\] VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 input_ctrl_inst.col_index\[29\] VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1401_ _0697_ net110 VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__nand2b_1
X_2450_ clknet_leaf_4_clk _0038_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_2381_ input_ctrl_inst.col_index\[12\] _0515_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__nor2_1
X_1263_ _0559_ _0598_ _0599_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__nor3_1
X_1332_ net73 _0655_ _0656_ net66 gencon_inst.mult_calc.out\[3\] VGND VGND VPWR VPWR
+ _0657_ sky130_fd_sc_hd__a32o_1
XFILLER_36_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput5 nRST VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2717_ clknet_leaf_21_clk _0261_ net159 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2579_ clknet_leaf_23_clk _0132_ net156 VGND VGND VPWR VPWR gencon_inst.operand2\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_2648_ clknet_leaf_27_clk _0197_ net151 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1950_ gencon_inst.operand2\[10\] net50 net33 net370 VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__a22o_1
X_1881_ _1212_ net52 _0988_ gencon_inst.key_read VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__or4b_1
X_2502_ clknet_leaf_32_clk _0067_ net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[7\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1315_ gencon_inst.operand2\[1\] gencon_inst.latched_keypad_input\[1\] VGND VGND
+ VPWR VPWR _0642_ sky130_fd_sc_hd__nor2_1
X_2364_ input_ctrl_inst.col_index\[5\] _0504_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__and2_1
X_2433_ input_ctrl_inst.col_index\[29\] input_ctrl_inst.col_index\[28\] _0547_ VGND
+ VGND VPWR VPWR _0551_ sky130_fd_sc_hd__and3_1
X_1246_ _0577_ _0580_ _0584_ _0585_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__o211a_1
X_2295_ _0445_ _0468_ _0470_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_22_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2080_ net36 _1140_ _1141_ net38 net275 VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__a32o_1
XFILLER_38_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1933_ net53 _0981_ net39 net15 VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__a22o_1
X_1864_ gencon_inst.operand1\[8\] net346 net48 VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__mux2_1
X_1795_ gencon_inst.latched_operator_input\[2\] net134 _0392_ _0963_ VGND VGND VPWR
+ VPWR _0964_ sky130_fd_sc_hd__and4_1
XFILLER_69_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2278_ input_ctrl_inst.scan_timer\[7\] _0458_ input_ctrl_inst.scan_timer\[8\] VGND
+ VGND VPWR VPWR _0460_ sky130_fd_sc_hd__a21o_1
X_2347_ net96 net216 net80 net283 VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__a22o_1
X_2416_ _0429_ _0508_ _1044_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__o21a_1
XFILLER_52_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1229_ gencon_inst.operand1\[1\] gencon_inst.latched_keypad_input\[1\] VGND VGND
+ VPWR VPWR _0571_ sky130_fd_sc_hd__or2_1
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1580_ _0793_ _0794_ gencon_inst.add_calc.main.GENERATE_ADDER\[11\].thingy.in1 VGND
+ VGND VPWR VPWR _0795_ sky130_fd_sc_hd__a21oi_1
XFILLER_7_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2132_ _1180_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2201_ input_ctrl_inst.col_index\[13\] input_ctrl_inst.col_index\[12\] input_ctrl_inst.col_index\[15\]
+ input_ctrl_inst.col_index\[14\] VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__or4_1
XFILLER_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2063_ _1032_ _1055_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1847_ gencon_inst.operand2\[7\] net335 net49 VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__mux2_1
X_1916_ _1012_ _1013_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__or2_1
XFILLER_22_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1778_ gencon_inst.ALU_in2\[10\] gencon_inst.ALU_in1\[10\] net64 VGND VGND VPWR VPWR
+ _0953_ sky130_fd_sc_hd__mux2_1
XFILLER_69_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1701_ net444 _0906_ net115 VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__mux2_1
X_2750_ clknet_leaf_27_clk _0294_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2681_ clknet_leaf_29_clk _0230_ net148 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1632_ _0807_ _0811_ _0845_ _0808_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__o31a_1
X_1563_ gencon_inst.operator_input\[0\] gencon_inst.key_read _0383_ _0387_ net54 VGND
+ VGND VPWR VPWR _0780_ sky130_fd_sc_hd__a41o_1
X_1494_ _0720_ _0722_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__xnor2_1
X_2115_ input_ctrl_inst.debounce_cnt\[13\] _1053_ _1132_ VGND VGND VPWR VPWR _1167_
+ sky130_fd_sc_hd__and3_1
XFILLER_39_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout38 _1133_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_2
Xfanout49 _0984_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_52_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2046_ _1107_ _1109_ _1112_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_17_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload19 clknet_leaf_14_clk VGND VGND VPWR VPWR clkload19/Y sky130_fd_sc_hd__inv_6
XFILLER_63_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2733_ clknet_leaf_21_clk _0277_ net159 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[12\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2802_ clknet_leaf_14_clk _0346_ net135 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfrtp_1
XFILLER_8_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2664_ clknet_leaf_31_clk net313 net146 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1615_ net106 gencon_inst.add_calc.main.in2\[2\] VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__nand2_1
X_1546_ _0760_ _0763_ _0761_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__o21ai_1
X_1477_ gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in1
+ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__nand2_1
XFILLER_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2595_ clknet_leaf_32_clk _0144_ net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2029_ gencon_inst.mult_calc.compCount.in2\[3\] _1088_ _1091_ _1094_ _1095_ VGND
+ VGND VPWR VPWR _1096_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_17_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold260 gencon_inst.add_calc.main.in2\[6\] VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 input_ctrl_inst.debounce_cnt\[17\] VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 gencon_inst.add_calc.main.in2\[0\] VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1400_ gencon_inst.addOrSub _0696_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__xnor2_1
X_1331_ _0653_ _0654_ _0652_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__o21ai_1
X_2380_ _0514_ _0515_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__nor2_1
XFILLER_64_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1262_ gencon_inst.operand1\[5\] _0591_ gencon_inst.operand1\[6\] VGND VGND VPWR
+ VPWR _0599_ sky130_fd_sc_hd__a21oi_1
XFILLER_36_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2716_ clknet_leaf_20_clk _0260_ net159 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_2647_ clknet_leaf_27_clk _0196_ net149 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2578_ clknet_leaf_23_clk _0131_ net157 VGND VGND VPWR VPWR gencon_inst.operand2\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_1529_ _0749_ _0750_ _0751_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__a21o_1
XFILLER_19_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1880_ _1035_ _1207_ _0380_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__o21ai_1
XFILLER_41_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2501_ clknet_leaf_32_clk net236 net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[6\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1314_ gencon_inst.operand2\[1\] gencon_inst.latched_keypad_input\[1\] VGND VGND
+ VPWR VPWR _0641_ sky130_fd_sc_hd__and2_1
X_2294_ _0469_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__inv_2
X_2432_ input_ctrl_inst.col_index\[28\] _0547_ input_ctrl_inst.col_index\[29\] VGND
+ VGND VPWR VPWR _0550_ sky130_fd_sc_hd__a21oi_1
X_2363_ input_ctrl_inst.col_index\[5\] _0504_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__nor2_1
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1245_ gencon_inst.operand1\[3\] gencon_inst.latched_keypad_input\[3\] VGND VGND
+ VPWR VPWR _0585_ sky130_fd_sc_hd__or2_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_25_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1863_ gencon_inst.operand1\[7\] net358 net49 VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1932_ gencon_inst.ALU_out\[13\] net69 net61 gencon_inst.mult_calc.out\[13\] VGND
+ VGND VPWR VPWR _1024_ sky130_fd_sc_hd__a22o_1
XFILLER_21_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1794_ gencon_inst.latched_operator_input\[0\] gencon_inst.latched_operator_input\[1\]
+ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__nor2_1
X_2415_ _0536_ _0538_ _0537_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__a21boi_1
XFILLER_69_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1228_ _0569_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__inv_2
X_2277_ net353 _0458_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__xor2_1
X_2346_ net96 net233 net80 gencon_inst.mult_calc.count.GENERATE_ADDER\[13\].thingy.in1
+ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__a22o_1
XFILLER_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_32_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2062_ net246 net277 net114 VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__a21o_1
X_2131_ input_ctrl_inst.debounce_cnt\[15\] input_ctrl_inst.debounce_cnt\[16\] _1171_
+ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_49_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ input_ctrl_inst.col_index\[5\] input_ctrl_inst.col_index\[4\] input_ctrl_inst.col_index\[7\]
+ input_ctrl_inst.col_index\[6\] VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__or4_1
XFILLER_34_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1777_ net360 _0952_ net113 VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_14_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
X_1846_ gencon_inst.operand2\[6\] net222 net49 VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__mux2_1
X_1915_ net53 _0975_ net39 net24 VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2329_ net118 net282 _0482_ _0492_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__a22o_1
XFILLER_27_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1631_ _0811_ _0845_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__nor2_1
X_1700_ _0903_ _0905_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2680_ clknet_leaf_28_clk _0229_ net149 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1562_ gencon_inst.mult_calc.out\[15\] _1212_ _0778_ net73 _0635_ VGND VGND VPWR
+ VPWR _0779_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_3_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
X_1493_ _0713_ _0721_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__or2_1
XFILLER_66_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2114_ input_ctrl_inst.debounce_cnt\[13\] _1163_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__or2_1
X_2045_ gencon_inst.mult_calc.compCount.in2\[8\] _1108_ _1111_ gencon_inst.mult_calc.compCount.in2\[9\]
+ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__o22a_1
Xfanout39 net40 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1829_ gencon_inst.operand2\[15\] gencon_inst.operand1\[15\] net76 VGND VGND VPWR
+ VPWR _0983_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2801_ clknet_leaf_13_clk _0345_ net137 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfrtp_1
XFILLER_44_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1614_ net106 gencon_inst.add_calc.main.in2\[2\] VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__or2_1
X_2732_ clknet_leaf_21_clk _0276_ net159 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[11\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2594_ clknet_leaf_32_clk _0143_ net139 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2663_ clknet_leaf_31_clk net341 net147 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_1476_ gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in1
+ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__nor2_1
X_1545_ gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in1
+ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_6_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2028_ gencon_inst.mult_calc.compCount.in2\[2\] _1074_ _1089_ VGND VGND VPWR VPWR
+ _1095_ sky130_fd_sc_hd__or3_1
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold283 gencon_inst.ALU_out\[7\] VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 input_ctrl_inst.debounce_cnt\[5\] VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold250 input_ctrl_inst.debounce_cnt\[4\] VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 gencon_inst.ALU_in2\[9\] VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1261_ _0583_ _0586_ gencon_inst.operand1\[4\] gencon_inst.operand1\[5\] gencon_inst.operand1\[6\]
+ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__o2111a_1
X_1330_ _0652_ _0653_ _0654_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__or3_1
XFILLER_30_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2715_ clknet_leaf_20_clk _0259_ net159 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2577_ clknet_leaf_25_clk _0130_ net155 VGND VGND VPWR VPWR gencon_inst.operand2\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_2646_ clknet_leaf_26_clk _0195_ net150 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1528_ _0749_ _0750_ _0751_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__nand3_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1459_ net365 net319 net98 VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__mux2_1
XFILLER_70_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2500_ clknet_leaf_32_clk net238 net139 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[5\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2431_ _0527_ _0549_ input_ctrl_inst.col_index\[28\] net58 VGND VGND VPWR VPWR _0103_
+ sky130_fd_sc_hd__a2bb2o_1
X_1244_ gencon_inst.operand1\[3\] gencon_inst.latched_keypad_input\[3\] VGND VGND
+ VPWR VPWR _0584_ sky130_fd_sc_hd__nand2_1
X_1313_ gencon_inst.operand2\[0\] net54 _0640_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__o21a_1
X_2293_ input_ctrl_inst.scan_timer\[13\] input_ctrl_inst.scan_timer\[14\] _0466_ VGND
+ VGND VPWR VPWR _0469_ sky130_fd_sc_hd__and3_1
X_2362_ _0503_ _0504_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__nor2_1
XFILLER_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2629_ clknet_leaf_26_clk _0178_ net144 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_73_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1862_ gencon_inst.operand1\[6\] net210 net49 VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__mux2_1
X_1931_ net205 net40 _1023_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__a21o_1
X_1793_ net118 _0960_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__nor2_1
XFILLER_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2414_ input_ctrl_inst.col_index\[23\] _0444_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__and2_1
XFILLER_69_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1227_ gencon_inst.operand1\[1\] gencon_inst.latched_keypad_input\[1\] VGND VGND
+ VPWR VPWR _0569_ sky130_fd_sc_hd__nand2_1
X_2276_ _0458_ _0459_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__nor2_1
X_2345_ net96 net221 net80 net227 VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__a22o_1
XFILLER_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2130_ input_ctrl_inst.debounce_cnt\[15\] _1171_ input_ctrl_inst.debounce_cnt\[16\]
+ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__a21o_1
XFILLER_19_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2061_ _1034_ _1073_ _1126_ net87 _1127_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__o221ai_1
X_1914_ gencon_inst.ALU_out\[7\] net70 net60 gencon_inst.mult_calc.out\[7\] VGND VGND
+ VPWR VPWR _1012_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1776_ gencon_inst.ALU_in2\[9\] gencon_inst.ALU_in1\[9\] net64 VGND VGND VPWR VPWR
+ _0952_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_62_Left_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1845_ gencon_inst.operand2\[5\] net231 net47 VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_71_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2328_ gencon_inst.keypad_input\[2\] net82 _0489_ _0491_ VGND VGND VPWR VPWR _0492_
+ sky130_fd_sc_hd__a22o_1
X_2259_ input_ctrl_inst.scan_timer\[3\] input_ctrl_inst.scan_timer\[2\] input_ctrl_inst.scan_timer\[5\]
+ input_ctrl_inst.scan_timer\[4\] VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__or4b_1
XFILLER_13_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1630_ _0815_ _0819_ _0842_ _0816_ _0812_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__o311a_1
XFILLER_8_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1561_ gencon_inst.operand2\[15\] _0692_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__xor2_1
X_1492_ _0704_ _0707_ _0710_ _0714_ _0708_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__o311a_1
XFILLER_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2113_ _1163_ _1165_ input_ctrl_inst.debounce_cnt\[12\] net37 VGND VGND VPWR VPWR
+ _0011_ sky130_fd_sc_hd__a2bb2o_1
X_2044_ _1079_ _1110_ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__nand2b_1
XFILLER_30_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1759_ net414 _0943_ net110 VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__mux2_1
X_1828_ net166 _0982_ net42 VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2731_ clknet_leaf_20_clk _0275_ net159 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[10\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2800_ clknet_leaf_6_clk _0344_ net134 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1613_ gencon_inst.add_calc.main.GENERATE_ADDER\[3\].thingy.in1 _0825_ _0826_ VGND
+ VGND VPWR VPWR _0828_ sky130_fd_sc_hd__nand3_1
XFILLER_67_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2593_ clknet_leaf_32_clk _0142_ net139 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2662_ clknet_leaf_31_clk _0211_ net147 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1544_ gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in1
+ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__or2_1
X_1475_ net103 _0705_ _0706_ net291 net91 VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__a32o_1
XFILLER_50_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2027_ gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.cIn gencon_inst.mult_calc.compCount.in2\[0\]
+ _1092_ _1093_ gencon_inst.mult_calc.compCount.in2\[1\] VGND VGND VPWR VPWR _1094_
+ sky130_fd_sc_hd__a32o_1
XFILLER_10_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold284 gencon_inst.ALU_out\[10\] VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 input_ctrl_inst.debounce_cnt\[6\] VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 gencon_inst.ALU_out\[12\] VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 input_ctrl_inst.scan_timer\[12\] VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 gencon_inst.mult_calc.compCount.in2\[4\] VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1260_ gencon_inst.operand1\[5\] net44 _0595_ _0597_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__o22a_1
XFILLER_49_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2714_ clknet_leaf_19_clk _0258_ net158 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_70_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2576_ clknet_leaf_25_clk _0129_ net155 VGND VGND VPWR VPWR gencon_inst.operand2\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_2645_ clknet_leaf_25_clk _0194_ net144 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1527_ _0743_ _0747_ _0744_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__o21ai_1
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1389_ net86 _1100_ net88 net237 VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__a2bb2o_1
X_1458_ net392 net384 net98 VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__mux2_1
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2361_ input_ctrl_inst.col_index\[4\] _0444_ _0502_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__and3_1
X_2430_ input_ctrl_inst.col_index\[28\] _0547_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__xnor2_1
X_1243_ gencon_inst.operand1\[3\] gencon_inst.latched_keypad_input\[3\] VGND VGND
+ VPWR VPWR _0583_ sky130_fd_sc_hd__and2_1
X_1312_ gencon_inst.mult_calc.out\[0\] net66 _0637_ _0639_ VGND VGND VPWR VPWR _0640_
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2292_ input_ctrl_inst.scan_timer\[13\] input_ctrl_inst.scan_timer\[12\] _0464_ input_ctrl_inst.scan_timer\[14\]
+ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__a31o_1
XFILLER_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2559_ clknet_leaf_16_clk _0112_ net152 VGND VGND VPWR VPWR gencon_inst.operand1\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_2628_ clknet_leaf_34_clk net372 net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_73_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1930_ gencon_inst.operand2\[12\] _0387_ net70 gencon_inst.ALU_out\[12\] _1022_ VGND
+ VGND VPWR VPWR _1023_ sky130_fd_sc_hd__a221o_1
XFILLER_14_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1861_ gencon_inst.operand1\[5\] net257 net47 VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__mux2_1
X_1792_ gencon_inst.read_input net52 VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__nand2_2
XFILLER_69_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2344_ net96 net276 net80 net297 VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__a22o_1
X_2413_ input_ctrl_inst.col_index\[21\] input_ctrl_inst.col_index\[22\] _0528_ _0530_
+ input_ctrl_inst.col_index\[23\] VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__a41o_1
X_1226_ gencon_inst.operand1\[0\] net44 _0567_ _0568_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__o22a_1
X_2275_ _0445_ _0457_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__nand2_1
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2060_ net286 net104 VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__nand2_1
XFILLER_19_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1913_ _1010_ _1011_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_32_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1775_ net357 _0951_ net113 VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__mux2_1
X_1844_ gencon_inst.operand2\[4\] net214 net47 VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__mux2_1
X_2327_ input_ctrl_inst.decoded_key\[2\] _1205_ input_ctrl_inst.decoded_key\[3\] VGND
+ VGND VPWR VPWR _0491_ sky130_fd_sc_hd__a21o_1
X_2258_ _0435_ _0446_ _0447_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__or3b_1
XFILLER_65_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2189_ net93 _1207_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__nor2_1
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1560_ net110 net106 _0698_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__o21a_1
XFILLER_8_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2112_ input_ctrl_inst.debounce_cnt\[12\] _1160_ _1164_ VGND VGND VPWR VPWR _1165_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_39_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1491_ _0718_ _0719_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__and2b_1
XFILLER_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2043_ gencon_inst.mult_calc.count.GENERATE_ADDER\[8\].thingy.in1 gencon_inst.mult_calc.count.GENERATE_ADDER\[7\].thingy.in1
+ _1077_ gencon_inst.mult_calc.count.GENERATE_ADDER\[9\].thingy.in1 VGND VGND VPWR
+ VPWR _1110_ sky130_fd_sc_hd__a31o_1
X_1827_ gencon_inst.operand2\[14\] gencon_inst.operand1\[14\] net76 VGND VGND VPWR
+ VPWR _0982_ sky130_fd_sc_hd__mux2_1
XFILLER_13_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1689_ net385 _0896_ net114 VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__mux2_1
X_1758_ gencon_inst.ALU_in2\[0\] gencon_inst.ALU_in1\[0\] net62 VGND VGND VPWR VPWR
+ _0943_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2730_ clknet_leaf_20_clk _0274_ net159 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[9\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2661_ clknet_leaf_31_clk _0210_ net142 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1612_ _0825_ _0826_ gencon_inst.add_calc.main.GENERATE_ADDER\[3\].thingy.in1 VGND
+ VGND VPWR VPWR _0827_ sky130_fd_sc_hd__a21oi_1
X_1543_ net405 net90 _0764_ net102 VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__a22o_1
X_1474_ _0703_ _0704_ _0701_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__o21ai_1
X_2592_ clknet_leaf_32_clk _0141_ net139 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2026_ gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.in1 gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.cIn
+ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__xnor2_1
Xhold285 gencon_inst.ALU_out\[6\] VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold241 gencon_inst.operator_input\[2\] VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 gencon_inst.mult_calc.adderSave\[2\] VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in2 VGND VGND VPWR
+ VPWR net412 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold263 input_ctrl_inst.col_index\[27\] VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 input_ctrl_inst.col_index\[26\] VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2713_ clknet_leaf_18_clk _0257_ net154 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_70_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2644_ clknet_leaf_34_clk _0193_ net144 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2575_ clknet_leaf_25_clk _0128_ net155 VGND VGND VPWR VPWR gencon_inst.operand2\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_1526_ gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in1
+ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__nand2_1
X_1457_ net400 net355 net98 VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__mux2_1
X_1388_ net86 _1097_ net88 net243 VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2009_ gencon_inst.mult_calc.count.GENERATE_ADDER\[5\].thingy.in1 gencon_inst.mult_calc.count.GENERATE_ADDER\[4\].thingy.in1
+ _1075_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__and3_1
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1311_ net73 _0638_ _0635_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__a21o_1
X_2291_ net363 _0466_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__xor2_1
X_2360_ _0444_ _0502_ input_ctrl_inst.col_index\[4\] VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__a21oi_1
XFILLER_64_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1242_ gencon_inst.operand1\[2\] net44 _0581_ _0582_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__o22a_1
XFILLER_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2627_ clknet_leaf_34_clk _0176_ net140 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
X_2558_ clknet_leaf_15_clk _0111_ net152 VGND VGND VPWR VPWR gencon_inst.operand1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2489_ clknet_leaf_3_clk _0054_ VGND VGND VPWR VPWR gencon_inst.operator_input\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1509_ _0733_ _0735_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_73_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_35_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_23_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1860_ gencon_inst.operand1\[4\] net258 net46 VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__mux2_1
XFILLER_36_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_26_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_14_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1791_ net52 VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__inv_2
X_2274_ input_ctrl_inst.scan_timer\[5\] input_ctrl_inst.scan_timer\[4\] input_ctrl_inst.scan_timer\[6\]
+ _0454_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__and4_1
X_2412_ _0535_ _0536_ _0534_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__o21ai_1
X_2343_ net96 net269 net80 gencon_inst.mult_calc.count.GENERATE_ADDER\[10\].thingy.in1
+ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_17_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_52_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1225_ gencon_inst.ALU_out\[0\] net68 net56 gencon_inst.mult_calc.out\[0\] VGND VGND
+ VPWR VPWR _0568_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_35_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1989_ net92 input_ctrl_inst.input_control_state\[1\] input_ctrl_inst.input_control_state\[0\]
+ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__and3b_1
XFILLER_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1843_ gencon_inst.operand2\[3\] net260 net47 VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__mux2_1
X_1912_ net53 _0974_ net39 net23 VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1774_ gencon_inst.ALU_in2\[8\] gencon_inst.ALU_in1\[8\] net63 VGND VGND VPWR VPWR
+ _0951_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_6_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_57_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2326_ net118 net271 _0482_ _0490_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__a22o_1
X_2257_ input_ctrl_inst.scan_timer\[7\] input_ctrl_inst.scan_timer\[6\] input_ctrl_inst.scan_timer\[9\]
+ input_ctrl_inst.scan_timer\[8\] VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__and4b_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2188_ gencon_inst.read_input _0378_ _0382_ _0390_ _1213_ VGND VGND VPWR VPWR _0391_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_9_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1490_ gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in1
+ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__nand2_1
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2111_ input_ctrl_inst.debounce_cnt\[12\] _1053_ _1132_ net35 VGND VGND VPWR VPWR
+ _1164_ sky130_fd_sc_hd__a31o_1
XFILLER_39_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1 input_ctrl_inst.RowMid\[3\] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dlygate4sd3_1
X_2042_ gencon_inst.mult_calc.compCount.in2\[7\] _1105_ _1108_ gencon_inst.mult_calc.compCount.in2\[8\]
+ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__a22o_1
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1826_ net219 _0981_ net42 VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__mux2_1
XFILLER_15_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1688_ _0893_ _0895_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__xnor2_1
X_1757_ net322 _0942_ net112 VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2309_ net125 net83 net314 VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_0_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1611_ net106 gencon_inst.add_calc.main.in2\[3\] VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_14_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2660_ clknet_leaf_31_clk net333 net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1542_ _0762_ _0763_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__xor2_1
X_1473_ _0701_ _0703_ _0704_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__or3_1
X_2591_ clknet_leaf_37_clk _0140_ net126 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2025_ gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.in1 gencon_inst.mult_calc.compCount.in2\[1\]
+ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_59_Left_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold253 input_ctrl_inst.debounce_cnt\[9\] VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__dlygate4sd3_1
X_2789_ clknet_leaf_14_clk _0333_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[15\] sky130_fd_sc_hd__dfxtp_1
X_1809_ gencon_inst.operand2\[5\] gencon_inst.operand1\[5\] net76 VGND VGND VPWR VPWR
+ _0973_ sky130_fd_sc_hd__mux2_1
Xhold220 input_ctrl_inst.scan_timer\[5\] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 gencon_inst.mult_calc.adderSave\[8\] VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 input_ctrl_inst.col_index\[7\] VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 input_ctrl_inst.debounce_cnt\[8\] VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 gencon_inst.ALU_in1\[15\] VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold286 input_ctrl_inst.col_index\[19\] VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2712_ clknet_leaf_16_clk _0256_ net154 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2574_ clknet_leaf_25_clk _0127_ net143 VGND VGND VPWR VPWR gencon_inst.operand2\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2643_ clknet_leaf_35_clk _0192_ net143 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1525_ gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in1
+ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__or2_1
X_1387_ net86 _1088_ net88 net247 VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__a2bb2o_1
X_1456_ net382 net265 net98 VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__mux2_1
XFILLER_70_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2008_ gencon_inst.mult_calc.count.GENERATE_ADDER\[3\].thingy.in1 gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.in1
+ gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.cIn gencon_inst.mult_calc.count.GENERATE_ADDER\[2\].thingy.in1
+ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__and4_1
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1241_ gencon_inst.ALU_out\[2\] net68 net56 gencon_inst.mult_calc.out\[2\] net43
+ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__a221o_1
X_1310_ gencon_inst.operand2\[0\] gencon_inst.latched_keypad_input\[0\] VGND VGND
+ VPWR VPWR _0638_ sky130_fd_sc_hd__nand2_1
X_2290_ _0466_ _0467_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__nor2_1
XFILLER_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2557_ clknet_leaf_15_clk _0110_ net152 VGND VGND VPWR VPWR gencon_inst.operand1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2626_ clknet_leaf_35_clk net304 net143 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2488_ clknet_leaf_7_clk _0053_ VGND VGND VPWR VPWR gencon_inst.operator_input\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1439_ net186 net168 net99 VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__mux2_1
X_1508_ _0725_ _0734_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__or2_1
XFILLER_62_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1790_ _0378_ _0387_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_44_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2411_ input_ctrl_inst.col_index\[21\] input_ctrl_inst.col_index\[22\] _0530_ _0527_
+ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__a31o_1
X_1224_ gencon_inst.operand1\[0\] gencon_inst.latched_keypad_input\[0\] net43 _0566_
+ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__o22a_1
XFILLER_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2273_ input_ctrl_inst.scan_timer\[5\] input_ctrl_inst.scan_timer\[4\] _0454_ input_ctrl_inst.scan_timer\[6\]
+ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__a31o_1
X_2342_ net96 net264 net80 net280 VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__a22o_1
XFILLER_52_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1988_ _1055_ net84 VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__nand2_1
X_2609_ clknet_leaf_33_clk _0158_ net139 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_73_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1773_ net367 _0950_ net112 VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__mux2_1
X_1842_ gencon_inst.operand2\[2\] net206 net47 VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__mux2_1
X_1911_ gencon_inst.ALU_out\[6\] net70 net60 gencon_inst.mult_calc.out\[6\] VGND VGND
+ VPWR VPWR _1010_ sky130_fd_sc_hd__a22o_1
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_31_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2187_ net76 _0389_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__nor2_1
X_2325_ gencon_inst.keypad_input\[1\] net82 _0487_ _0489_ VGND VGND VPWR VPWR _0490_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_40_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2256_ input_ctrl_inst.scan_timer\[11\] input_ctrl_inst.scan_timer\[10\] input_ctrl_inst.scan_timer\[13\]
+ input_ctrl_inst.scan_timer\[12\] VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__or4_1
XFILLER_21_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2110_ input_ctrl_inst.debounce_cnt\[12\] _1160_ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__and2_1
Xhold2 input_ctrl_inst.RowMid\[2\] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dlygate4sd3_1
X_2041_ gencon_inst.mult_calc.count.GENERATE_ADDER\[8\].thingy.in1 _1078_ VGND VGND
+ VPWR VPWR _1108_ sky130_fd_sc_hd__xor2_1
XFILLER_62_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1756_ gencon_inst.ALU_in1\[14\] gencon_inst.ALU_in2\[14\] net63 VGND VGND VPWR VPWR
+ _0942_ sky130_fd_sc_hd__mux2_1
X_1825_ gencon_inst.operand2\[13\] gencon_inst.operand1\[13\] net77 VGND VGND VPWR
+ VPWR _0981_ sky130_fd_sc_hd__mux2_1
X_1687_ _0846_ _0894_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__xnor2_1
X_2308_ input_ctrl_inst.decoded_key\[0\] input_ctrl_inst.decoded_key\[1\] _1204_ net83
+ net125 VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__o311a_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2239_ _0433_ _0434_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__or2_1
XFILLER_70_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1610_ net106 gencon_inst.add_calc.main.in2\[3\] VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__or2_1
XFILLER_60_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2590_ clknet_leaf_37_clk _0139_ net126 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1472_ gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in1
+ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__nor2_1
X_1541_ _0754_ _0758_ _0755_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__o21a_1
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2024_ _1074_ _1089_ gencon_inst.mult_calc.compCount.in2\[2\] VGND VGND VPWR VPWR
+ _1091_ sky130_fd_sc_hd__o21a_1
XFILLER_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1739_ net325 _0933_ net111 VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__mux2_1
Xhold287 gencon_inst.ALU_out\[3\] VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 gencon_inst.ALU_out\[2\] VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 gencon_inst.add_calc.main.a0.in1 VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__dlygate4sd3_1
X_2788_ clknet_leaf_24_clk _0332_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[14\] sky130_fd_sc_hd__dfxtp_1
Xhold210 gencon_inst.mult_calc.INn2\[10\] VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__dlygate4sd3_1
X_1808_ net176 _0972_ net41 VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__mux2_1
Xhold243 input_ctrl_inst.col_index\[15\] VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold265 input_ctrl_inst.col_index\[14\] VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 gencon_inst.mult_calc.compCount.in2\[5\] VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 gencon_inst.mult_calc.compCount.in2\[13\] VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2711_ clknet_leaf_17_clk _0255_ net153 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2573_ clknet_leaf_15_clk _0126_ net152 VGND VGND VPWR VPWR gencon_inst.operand2\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_2642_ clknet_leaf_35_clk _0191_ net143 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1524_ net391 net89 _0748_ net102 VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__a22o_1
X_1386_ net103 _1090_ net88 net232 VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__a22o_1
X_1455_ net378 net308 net99 VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__mux2_1
XFILLER_42_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2007_ gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.in1 gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.cIn
+ gencon_inst.mult_calc.count.GENERATE_ADDER\[2\].thingy.in1 VGND VGND VPWR VPWR _1074_
+ sky130_fd_sc_hd__and3_1
XFILLER_50_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1240_ _0580_ net72 _0579_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__and3b_1
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2556_ clknet_leaf_15_clk _0109_ net152 VGND VGND VPWR VPWR gencon_inst.operand1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2487_ clknet_leaf_3_clk _0052_ VGND VGND VPWR VPWR equal_input sky130_fd_sc_hd__dfxtp_1
X_1507_ _0713_ _0718_ _0721_ _0726_ _0719_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__o311a_1
X_2625_ clknet_leaf_34_clk net324 net139 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
X_1369_ gencon_inst.operand2\[11\] _0685_ net55 VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__mux2_1
X_1438_ net194 net180 net99 VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__mux2_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2410_ input_ctrl_inst.col_index\[21\] _0530_ input_ctrl_inst.col_index\[22\] VGND
+ VGND VPWR VPWR _0535_ sky130_fd_sc_hd__a21oi_1
X_2341_ net96 net254 net80 gencon_inst.mult_calc.count.GENERATE_ADDER\[8\].thingy.in1
+ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__a22o_1
X_1223_ gencon_inst.operand1\[0\] gencon_inst.latched_keypad_input\[0\] _0559_ VGND
+ VGND VPWR VPWR _0566_ sky130_fd_sc_hd__a21oi_1
X_2272_ net380 _0456_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1987_ net92 input_ctrl_inst.input_control_state\[1\] input_ctrl_inst.input_control_state\[0\]
+ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__nor3b_1
X_2608_ clknet_leaf_35_clk _0157_ net129 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2539_ clknet_leaf_37_clk _0100_ net127 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1910_ _1008_ _1009_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_32_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1772_ gencon_inst.ALU_in2\[7\] gencon_inst.ALU_in1\[7\] net63 VGND VGND VPWR VPWR
+ _0950_ sky130_fd_sc_hd__mux2_1
X_1841_ gencon_inst.operand2\[1\] net281 net46 VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__mux2_1
XFILLER_42_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2324_ net83 _1204_ _0488_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__and3_1
XFILLER_65_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2186_ gencon_inst.read_input equal_input VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__or2_1
X_2255_ net119 net59 VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__or2_1
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2040_ gencon_inst.mult_calc.compCount.in2\[6\] _1103_ _1104_ _1101_ _1106_ VGND
+ VGND VPWR VPWR _1107_ sky130_fd_sc_hd__o221a_1
Xhold3 input_ctrl_inst.RowMid\[1\] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_30_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1686_ _0807_ _0808_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__nand2b_1
X_1755_ net368 _0941_ net112 VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__mux2_1
X_1824_ net209 _0980_ net42 VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__mux2_1
XFILLER_57_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2307_ input_ctrl_inst.decoded_key\[0\] input_ctrl_inst.decoded_key\[1\] VGND VGND
+ VPWR VPWR _0477_ sky130_fd_sc_hd__or2_1
XFILLER_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2238_ _0433_ net117 input_ctrl_inst.col_index\[1\] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__or3b_1
X_2169_ gencon_inst.gencon_state\[1\] gencon_inst.gencon_state\[0\] _1036_ gencon_inst.gencon_state\[2\]
+ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_0_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1540_ _0760_ _0761_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__nand2b_1
XFILLER_12_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1471_ gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in1
+ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_65_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2023_ _1074_ _1089_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__nor2_1
X_1807_ gencon_inst.operand2\[4\] gencon_inst.operand1\[4\] net76 VGND VGND VPWR VPWR
+ _0972_ sky130_fd_sc_hd__mux2_1
Xhold200 gencon_inst.add_calc.main.GENERATE_ADDER\[9\].thingy.in1 VGND VGND VPWR VPWR
+ net360 sky130_fd_sc_hd__dlygate4sd3_1
X_1669_ _0819_ _0820_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__and2b_1
Xhold244 gencon_inst.add_calc.main.GENERATE_ADDER\[4\].thingy.in1 VGND VGND VPWR VPWR
+ net404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 gencon_inst.ALU_out\[13\] VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__dlygate4sd3_1
X_1738_ gencon_inst.ALU_in1\[5\] gencon_inst.ALU_in2\[5\] net65 VGND VGND VPWR VPWR
+ _0933_ sky130_fd_sc_hd__mux2_1
X_2787_ clknet_leaf_24_clk _0331_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[13\] sky130_fd_sc_hd__dfxtp_1
Xhold266 input_ctrl_inst.debounce_cnt\[16\] VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 input_ctrl_inst.debounce_cnt\[2\] VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold233 gencon_inst.mult_calc.INn2\[7\] VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 gencon_inst.mult_calc.adderSave\[10\] VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold222 gencon_inst.mult_calc.compCount.in2\[3\] VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in2 VGND VGND VPWR
+ VPWR net371 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2710_ clknet_leaf_17_clk _0254_ net153 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2572_ clknet_leaf_15_clk _0125_ net143 VGND VGND VPWR VPWR gencon_inst.operand2\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_2641_ clknet_leaf_35_clk _0190_ net143 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1523_ _0745_ _0747_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__xnor2_1
X_1454_ net350 net239 net99 VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__mux2_1
XFILLER_67_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1385_ net86 _1093_ net88 net251 VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2006_ net98 _1073_ net94 VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__a21o_1
X_2839_ clknet_leaf_8_clk input_ctrl_inst.next_state\[2\] net131 VGND VGND VPWR VPWR
+ input_ctrl_inst.input_control_state\[2\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_38_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_41_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_30_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2624_ clknet_leaf_35_clk net327 net143 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
X_2555_ clknet_leaf_14_clk _0108_ net135 VGND VGND VPWR VPWR gencon_inst.operand1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2486_ clknet_leaf_8_clk _0017_ net131 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_1506_ _0731_ _0732_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__and2b_1
X_1437_ net104 gencon_inst.mult_calc.finish _0700_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__mux2_1
XFILLER_55_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1299_ net72 _0626_ _0627_ _0628_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__a31o_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1368_ _0683_ _0684_ gencon_inst.mult_calc.out\[11\] net67 VGND VGND VPWR VPWR _0685_
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_38_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2271_ net119 net59 _0454_ input_ctrl_inst.scan_timer\[4\] _0456_ VGND VGND VPWR
+ VPWR _0036_ sky130_fd_sc_hd__o221a_1
X_2340_ net96 net242 net80 gencon_inst.mult_calc.count.GENERATE_ADDER\[7\].thingy.in1
+ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__a22o_1
X_1222_ _0379_ net56 _0382_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__a21o_2
XFILLER_25_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1986_ net92 net30 _1056_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_35_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_9_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
X_2607_ clknet_leaf_35_clk _0156_ net128 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2469_ clknet_leaf_8_clk _0018_ net132 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2538_ clknet_leaf_38_clk _0099_ net121 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1840_ gencon_inst.operand2\[0\] net256 net46 VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__mux2_1
XFILLER_42_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1771_ net354 _0949_ net112 VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2323_ input_ctrl_inst.decoded_key\[3\] _0477_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__nand2_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2254_ net58 VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__inv_2
XFILLER_65_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2185_ gencon_inst.gencon_state\[3\] gencon_inst.gencon_state\[2\] gencon_inst.gencon_state\[1\]
+ net93 VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__or4bb_1
X_1969_ net114 VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__inv_2
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold4 input_ctrl_inst.RowMid\[0\] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_62_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1823_ gencon_inst.operand2\[12\] gencon_inst.operand1\[12\] net77 VGND VGND VPWR
+ VPWR _0980_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1685_ net31 _0892_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__nand2_1
X_1754_ gencon_inst.ALU_in1\[13\] gencon_inst.ALU_in2\[13\] net63 VGND VGND VPWR VPWR
+ _0941_ sky130_fd_sc_hd__mux2_1
XFILLER_57_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2306_ net173 _0475_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__xnor2_1
X_2237_ input_ctrl_inst.col_index\[1\] _0433_ net117 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__or3b_1
X_2099_ input_ctrl_inst.debounce_cnt\[9\] _1151_ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__and2_1
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2168_ net93 gencon_inst.ALU_finish _1207_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_0_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1470_ net103 _0701_ _0702_ net395 net91 VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__a32o_1
XFILLER_69_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2022_ gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.in1 gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.cIn
+ gencon_inst.mult_calc.count.GENERATE_ADDER\[2\].thingy.in1 VGND VGND VPWR VPWR _1089_
+ sky130_fd_sc_hd__a21oi_1
Xhold201 gencon_inst.add_calc.main.GENERATE_ADDER\[11\].thingy.in1 VGND VGND VPWR
+ VPWR net361 sky130_fd_sc_hd__dlygate4sd3_1
X_2786_ clknet_leaf_22_clk _0330_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[12\] sky130_fd_sc_hd__dfxtp_1
X_1806_ net188 _0971_ net41 VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_28_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1599_ net107 gencon_inst.add_calc.main.in2\[6\] VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__nand2_1
X_1668_ _0874_ _0877_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__or2_1
X_1737_ net339 _0932_ net111 VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__mux2_1
Xhold289 gencon_inst.ALU_out\[4\] VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold256 gencon_inst.ALU_in2\[8\] VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 gencon_inst.operand1\[15\] VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 input_ctrl_inst.debounce_cnt\[18\] VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_37_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold245 gencon_inst.mult_calc.adderSave\[11\] VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 input_ctrl_inst.col_index\[13\] VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 input_ctrl_inst.col_index\[9\] VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 _0177_ VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_55_Left_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_64_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2640_ clknet_leaf_35_clk _0189_ net129 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2571_ clknet_leaf_15_clk _0124_ net135 VGND VGND VPWR VPWR gencon_inst.operand2\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_1522_ _0738_ _0746_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__or2_1
X_1453_ net267 gencon_inst.mult_calc.INn2\[0\] net99 VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__mux2_1
XFILLER_55_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1384_ gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.cIn net86 net228 net88
+ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__a2bb2o_1
X_2005_ _1069_ _1070_ _1072_ VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__or3_1
XFILLER_50_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2769_ clknet_leaf_22_clk _0313_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[11\] sky130_fd_sc_hd__dfxtp_1
X_2838_ clknet_leaf_7_clk input_ctrl_inst.next_state\[1\] net131 VGND VGND VPWR VPWR
+ input_ctrl_inst.input_control_state\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2554_ clknet_leaf_14_clk _0107_ net135 VGND VGND VPWR VPWR gencon_inst.operand1\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_30_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2623_ clknet_leaf_36_clk _0172_ net129 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2485_ clknet_leaf_8_clk _0016_ net131 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_1367_ _1029_ _0680_ _1211_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__a21o_1
X_1436_ net86 net79 VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__nand2_1
X_1505_ gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in1
+ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__nand2_1
XFILLER_55_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1298_ gencon_inst.ALU_out\[13\] net70 net57 gencon_inst.mult_calc.out\[13\] _0565_
+ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_38_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1221_ _0379_ net56 _0382_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__a21oi_1
X_2270_ input_ctrl_inst.scan_timer\[4\] _0454_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__nand2_1
XFILLER_6_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1985_ input_ctrl_inst.input_control_state\[1\] input_ctrl_inst.input_control_state\[0\]
+ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__nor2_1
X_2606_ clknet_leaf_35_clk _0155_ net128 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2537_ clknet_leaf_38_clk _0098_ net121 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2468_ clknet_leaf_8_clk _0008_ net132 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_2399_ net58 _0500_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__or2_1
X_1419_ gencon_inst.mult_calc.out\[14\] net399 net105 VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__mux2_1
XFILLER_73_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire84 _1058_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_1
XFILLER_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout160 net5 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__buf_2
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1770_ gencon_inst.ALU_in2\[6\] gencon_inst.ALU_in1\[6\] net65 VGND VGND VPWR VPWR
+ _0949_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2184_ gencon_inst.gencon_state\[1\] gencon_inst.gencon_state\[0\] _1036_ _1037_
+ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__and4_4
X_2322_ _1205_ _0477_ _0483_ input_ctrl_inst.decoded_key\[3\] VGND VGND VPWR VPWR
+ _0487_ sky130_fd_sc_hd__a31o_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2253_ _1059_ _0437_ _0438_ _0442_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__or4_1
XFILLER_25_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1899_ gencon_inst.ALU_out\[2\] net68 net60 gencon_inst.mult_calc.out\[2\] VGND VGND
+ VPWR VPWR _1002_ sky130_fd_sc_hd__a22o_1
X_1968_ net103 VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__inv_2
XFILLER_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold5 gencon_inst.prev_read_input VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dlygate4sd3_1
X_1753_ net349 _0940_ net112 VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__mux2_1
X_1822_ net177 _0979_ net42 VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1684_ _0879_ _0881_ _0886_ _0890_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__or4_1
XFILLER_72_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2167_ _1207_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__inv_2
XFILLER_38_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2305_ _0475_ _0476_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_13_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2236_ net117 input_ctrl_inst.col_index\[1\] VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__nand2_1
XFILLER_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2098_ net35 _1151_ input_ctrl_inst.debounce_cnt\[9\] VGND VGND VPWR VPWR _1154_
+ sky130_fd_sc_hd__a21o_1
XFILLER_53_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2021_ gencon_inst.mult_calc.count.GENERATE_ADDER\[3\].thingy.in1 _1074_ VGND VGND
+ VPWR VPWR _1088_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_65_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold202 gencon_inst.add_calc.main.GENERATE_ADDER\[13\].thingy.in1 VGND VGND VPWR
+ VPWR net362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 gencon_inst.add_calc.main.GENERATE_ADDER\[14\].thingy.in1 VGND VGND VPWR
+ VPWR net373 sky130_fd_sc_hd__dlygate4sd3_1
X_1736_ gencon_inst.ALU_in1\[4\] gencon_inst.ALU_in2\[4\] net62 VGND VGND VPWR VPWR
+ _0932_ sky130_fd_sc_hd__mux2_1
X_2785_ clknet_leaf_21_clk _0329_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[11\] sky130_fd_sc_hd__dfxtp_1
X_1805_ gencon_inst.operand2\[3\] gencon_inst.operand1\[3\] net76 VGND VGND VPWR VPWR
+ _0971_ sky130_fd_sc_hd__mux2_1
Xhold224 gencon_inst.mult_calc.INn2\[5\] VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 gencon_inst.mult_calc.adderSave\[0\] VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__dlygate4sd3_1
X_1598_ net107 gencon_inst.add_calc.main.in2\[6\] VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__or2_1
Xhold279 gencon_inst.ALU_out\[14\] VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__dlygate4sd3_1
X_1667_ net449 _0878_ net114 VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__mux2_1
Xhold246 gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in2 VGND VGND VPWR
+ VPWR net406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 input_ctrl_inst.col_index\[20\] VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 input_ctrl_inst.col_index\[31\] VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2219_ input_ctrl_inst.col_index\[28\] input_ctrl_inst.col_index\[31\] input_ctrl_inst.col_index\[30\]
+ _0417_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__or4_1
XFILLER_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2570_ clknet_leaf_5_clk _0123_ net128 VGND VGND VPWR VPWR gencon_inst.operand2\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_10_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1521_ _0725_ _0731_ _0734_ _0739_ _0732_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__o311a_1
X_1452_ net170 net166 net100 VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__mux2_1
X_1383_ net100 net102 VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__nor2_1
XFILLER_35_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2004_ gencon_inst.mult_calc.INn2\[13\] gencon_inst.mult_calc.INn2\[12\] gencon_inst.mult_calc.INn2\[14\]
+ _1071_ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__or4_1
XFILLER_50_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2699_ clknet_leaf_19_clk _0243_ net158 VGND VGND VPWR VPWR gencon_inst.ALU_out\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1719_ net115 net437 _0920_ _0921_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__o22a_1
X_2768_ clknet_leaf_22_clk _0312_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[10\] sky130_fd_sc_hd__dfxtp_1
X_2837_ clknet_leaf_7_clk input_ctrl_inst.next_state\[0\] net131 VGND VGND VPWR VPWR
+ input_ctrl_inst.input_control_state\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_58_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2553_ clknet_leaf_2_clk net161 net123 VGND VGND VPWR VPWR input_ctrl_inst.RowSync\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_1504_ gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in1
+ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__nor2_1
X_2622_ clknet_leaf_36_clk _0171_ net126 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.a0.in2
+ sky130_fd_sc_hd__dfrtp_1
X_2484_ clknet_leaf_8_clk _0015_ net131 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_1366_ gencon_inst.operand2\[11\] gencon_inst.operand2\[10\] gencon_inst.operand2\[9\]
+ _0674_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__and4_1
XFILLER_28_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1435_ net97 gencon_inst.mult_calc.adderSave\[14\] net295 net80 VGND VGND VPWR VPWR
+ _0185_ sky130_fd_sc_hd__a22o_1
X_1297_ gencon_inst.operand1\[13\] _0622_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_38_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_1_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1220_ net72 net71 VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__nor2_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1984_ _1055_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_43_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2467_ clknet_leaf_2_clk _0030_ net124 VGND VGND VPWR VPWR input_ctrl_inst.decoded_key\[3\]
+ sky130_fd_sc_hd__dfstp_2
X_2605_ clknet_leaf_4_clk _0154_ net128 VGND VGND VPWR VPWR gencon_inst.mult_calc.diffSign
+ sky130_fd_sc_hd__dfrtp_1
X_2536_ clknet_leaf_37_clk _0097_ net127 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_1349_ gencon_inst.operand2\[6\] net55 _0670_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__o21a_1
X_2398_ _0524_ _0525_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__nor2_1
X_1418_ gencon_inst.mult_calc.out\[13\] net285 net105 VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__mux2_1
Xfanout150 net151 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2321_ net118 net299 _0482_ _0486_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__a22o_1
XFILLER_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2183_ _0384_ _0385_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__nand2_1
X_2252_ input_ctrl_inst.scan_timer\[10\] _0435_ _0436_ _0441_ VGND VGND VPWR VPWR
+ _0442_ sky130_fd_sc_hd__or4_1
XFILLER_33_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1898_ _1000_ _1001_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__or2_1
X_1967_ gencon_inst.mult_calc.compCount.in2\[14\] VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__inv_2
XFILLER_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2519_ clknet_leaf_0_clk _0080_ net122 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold6 gencon_inst.mult_calc.INn1\[14\] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1683_ net443 _0891_ net114 VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_10_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
X_1752_ gencon_inst.ALU_in1\[12\] gencon_inst.ALU_in2\[12\] net63 VGND VGND VPWR VPWR
+ _0940_ sky130_fd_sc_hd__mux2_1
X_1821_ gencon_inst.operand2\[11\] gencon_inst.operand1\[11\] net77 VGND VGND VPWR
+ VPWR _0979_ sky130_fd_sc_hd__mux2_1
X_2304_ input_ctrl_inst.scan_timer\[18\] _0473_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_68_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2097_ net424 net38 net35 _1153_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__a22o_1
XFILLER_53_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2166_ gencon_inst.gencon_state\[3\] _1037_ gencon_inst.gencon_state\[1\] VGND VGND
+ VPWR VPWR _1207_ sky130_fd_sc_hd__or3b_4
XFILLER_38_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2235_ net116 _0411_ _0429_ _0432_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__or4_1
XFILLER_53_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2020_ gencon_inst.mult_calc.compCount.in2\[11\] _1086_ VGND VGND VPWR VPWR _1087_
+ sky130_fd_sc_hd__and2_1
XFILLER_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1735_ net315 _0931_ net111 VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__mux2_1
X_1666_ _0875_ _0877_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__xnor2_1
Xhold225 gencon_inst.ALU_out\[8\] VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__dlygate4sd3_1
X_2784_ clknet_leaf_22_clk _0328_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold214 gencon_inst.mult_calc.INn2\[12\] VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__dlygate4sd3_1
X_1804_ net171 _0970_ net41 VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__mux2_1
Xhold203 input_ctrl_inst.scan_timer\[13\] VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 input_ctrl_inst.col_index\[10\] VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 input_ctrl_inst.col_index\[24\] VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 gencon_inst.mult_calc.compCount.in2\[8\] VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 gencon_inst.mult_calc.main.a0.in2 VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__dlygate4sd3_1
X_1597_ gencon_inst.add_calc.main.GENERATE_ADDER\[7\].thingy.in1 _0809_ _0810_ VGND
+ VGND VPWR VPWR _0812_ sky130_fd_sc_hd__nand3_1
X_2149_ _1033_ input_ctrl_inst.RowSync\[1\] input_ctrl_inst.RowSync\[3\] VGND VGND
+ VPWR VPWR _1193_ sky130_fd_sc_hd__o21a_1
X_2218_ input_ctrl_inst.col_index\[25\] input_ctrl_inst.col_index\[27\] input_ctrl_inst.col_index\[26\]
+ input_ctrl_inst.col_index\[29\] VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__or4_1
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1520_ _0743_ _0744_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_10_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1382_ gencon_inst.read_input net82 _1206_ _1043_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__a22o_1
X_1451_ net278 net219 net101 VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__mux2_1
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2003_ gencon_inst.mult_calc.INn2\[9\] gencon_inst.mult_calc.INn2\[8\] gencon_inst.mult_calc.INn2\[11\]
+ gencon_inst.mult_calc.INn2\[10\] VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__or4_1
X_2836_ clknet_leaf_4_clk net200 VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1649_ net85 _0862_ _0863_ _0861_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__o31a_1
X_2698_ clknet_leaf_17_clk _0242_ net153 VGND VGND VPWR VPWR gencon_inst.ALU_out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1718_ _0917_ _0919_ net115 VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__o21ai_1
X_2767_ clknet_leaf_22_clk _0311_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2483_ clknet_leaf_8_clk _0014_ net131 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_2621_ clknet_leaf_5_clk _0170_ net129 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_2552_ clknet_leaf_2_clk net162 net123 VGND VGND VPWR VPWR input_ctrl_inst.RowSync\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_1503_ net103 _0729_ _0730_ net289 net88 VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__a32o_1
X_1296_ gencon_inst.operand1\[13\] _0622_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__nand2_1
X_1365_ gencon_inst.operand2\[10\] _0682_ net55 VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__mux2_1
X_1434_ net97 gencon_inst.mult_calc.adderSave\[13\] net273 net81 VGND VGND VPWR VPWR
+ _0184_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_38_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2819_ clknet_leaf_5_clk gencon_inst.next_state\[2\] net134 VGND VGND VPWR VPWR gencon_inst.gencon_state\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_11_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2604_ clknet_leaf_13_clk net310 net136 VGND VGND VPWR VPWR gencon_inst.add_calc.sameSignVal
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_43_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1983_ input_ctrl_inst.RowSync\[2\] input_ctrl_inst.RowSync\[0\] input_ctrl_inst.RowSync\[1\]
+ input_ctrl_inst.RowSync\[3\] VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__and4_4
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2466_ clknet_leaf_2_clk _0029_ net124 VGND VGND VPWR VPWR input_ctrl_inst.decoded_key\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_1417_ gencon_inst.mult_calc.out\[12\] net301 net105 VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__mux2_1
X_2535_ clknet_leaf_37_clk _0096_ net127 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_68_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1279_ gencon_inst.operand1\[9\] _0606_ _0612_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__o21a_1
X_1348_ gencon_inst.mult_calc.out\[6\] net66 _0669_ net73 _0635_ VGND VGND VPWR VPWR
+ _0670_ sky130_fd_sc_hd__a221o_1
X_2397_ input_ctrl_inst.col_index\[19\] _0412_ _0520_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__and3_1
XFILLER_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout151 net160 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__buf_2
Xfanout140 net145 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
XFILLER_15_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2320_ gencon_inst.keypad_input\[0\] net83 _0484_ _0485_ VGND VGND VPWR VPWR _0486_
+ sky130_fd_sc_hd__o22a_1
X_2251_ input_ctrl_inst.scan_timer\[11\] input_ctrl_inst.scan_timer\[8\] input_ctrl_inst.scan_timer\[9\]
+ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__nand3b_1
XFILLER_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2182_ gencon_inst.operator_input\[2\] _0378_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_48_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1966_ net128 VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__inv_2
X_1897_ net52 _0969_ net40 net18 VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__a22o_1
X_2449_ clknet_leaf_4_clk _0037_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_2518_ clknet_leaf_0_clk _0079_ net122 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_54_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold7 gencon_inst.mult_calc.INn1\[7\] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__dlygate4sd3_1
X_1820_ net169 _0978_ net42 VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__mux2_1
XFILLER_30_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1682_ _0888_ _0890_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__xnor2_1
X_1751_ net331 _0939_ net113 VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__mux2_1
X_2303_ input_ctrl_inst.scan_timer\[18\] _0473_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__nand2_1
X_2234_ _0398_ _0429_ _0432_ VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__or3_1
X_2096_ _1151_ _1152_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__nor2_1
X_2165_ net351 _1206_ _1188_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__o21a_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1949_ gencon_inst.operand2\[9\] net50 net33 net298 VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2783_ clknet_leaf_22_clk _0327_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[9\] sky130_fd_sc_hd__dfxtp_1
X_1803_ gencon_inst.operand2\[2\] gencon_inst.operand1\[2\] net76 VGND VGND VPWR VPWR
+ _0970_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold204 gencon_inst.add_calc.main.GENERATE_ADDER\[3\].thingy.in1 VGND VGND VPWR VPWR
+ net364 sky130_fd_sc_hd__dlygate4sd3_1
X_1596_ _0809_ _0810_ gencon_inst.add_calc.main.GENERATE_ADDER\[7\].thingy.in1 VGND
+ VGND VPWR VPWR _0811_ sky130_fd_sc_hd__a21oi_1
X_1665_ _0840_ _0876_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__xnor2_1
X_1734_ gencon_inst.ALU_in1\[3\] gencon_inst.ALU_in2\[3\] net62 VGND VGND VPWR VPWR
+ _0931_ sky130_fd_sc_hd__mux2_1
Xhold248 net17 VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 gencon_inst.ALU_in1\[9\] VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 gencon_inst.operator_input\[1\] VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 input_ctrl_inst.scan_timer\[2\] VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 gencon_inst.mult_calc.adderSave\[4\] VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2217_ _0402_ _0407_ _0409_ _0410_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_64_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2079_ input_ctrl_inst.debounce_cnt\[1\] input_ctrl_inst.debounce_cnt\[0\] input_ctrl_inst.debounce_cnt\[2\]
+ input_ctrl_inst.debounce_cnt\[3\] VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__a31o_1
X_2148_ _1188_ _1192_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_24_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1450_ net220 net209 net101 VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__mux2_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1381_ gencon_inst.operand2\[14\] _0694_ net54 VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2002_ gencon_inst.mult_calc.INn2\[1\] gencon_inst.mult_calc.INn2\[0\] gencon_inst.mult_calc.INn2\[3\]
+ gencon_inst.mult_calc.INn2\[2\] VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__or4_1
X_2766_ clknet_leaf_16_clk _0310_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[8\] sky130_fd_sc_hd__dfxtp_1
X_2835_ clknet_leaf_26_clk _0375_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_1648_ _0781_ net32 _0860_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__a21oi_1
X_1579_ net108 gencon_inst.add_calc.main.in2\[11\] VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__nand2_1
X_2697_ clknet_leaf_18_clk _0241_ net154 VGND VGND VPWR VPWR gencon_inst.ALU_out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1717_ _0917_ _0919_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__and2_1
XFILLER_26_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2620_ clknet_leaf_33_clk _0169_ net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_2482_ clknet_leaf_8_clk _0013_ net131 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1433_ net97 gencon_inst.mult_calc.adderSave\[12\] net287 net81 VGND VGND VPWR VPWR
+ _0183_ sky130_fd_sc_hd__a22o_1
X_1502_ _0727_ _0728_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__nand2_1
X_2551_ clknet_leaf_1_clk net163 net123 VGND VGND VPWR VPWR input_ctrl_inst.RowSync\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_1295_ gencon_inst.operand1\[12\] net45 _0624_ _0625_ VGND VGND VPWR VPWR _0119_
+ sky130_fd_sc_hd__o22a_1
X_1364_ net74 _0680_ _0681_ net67 gencon_inst.mult_calc.out\[10\] VGND VGND VPWR VPWR
+ _0682_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_38_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2818_ clknet_leaf_6_clk gencon_inst.next_state\[1\] net134 VGND VGND VPWR VPWR gencon_inst.gencon_state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_2749_ clknet_leaf_27_clk _0293_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_72_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1982_ _1051_ _1053_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_43_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2534_ clknet_leaf_38_clk _0095_ net121 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_2603_ clknet_leaf_29_clk net217 net148 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_1347_ _0667_ _0668_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__nor2_1
X_2465_ clknet_leaf_3_clk _0028_ net124 VGND VGND VPWR VPWR input_ctrl_inst.decoded_key\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_1416_ gencon_inst.mult_calc.out\[11\] net405 net105 VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__mux2_1
XFILLER_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2396_ _0412_ _0520_ input_ctrl_inst.col_index\[19\] VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__a21oi_1
X_1278_ _0559_ _0611_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__nor2_1
XFILLER_28_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout152 net155 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_4
Xfanout141 net145 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_4
Xfanout130 net5 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__buf_2
XFILLER_19_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2250_ net124 _1055_ net84 input_ctrl_inst.scan_timer\[0\] VGND VGND VPWR VPWR _0440_
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_48_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2181_ gencon_inst.operator_input\[1\] _0378_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__nand2_1
X_1965_ gencon_inst.gencon_state\[2\] VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__inv_2
XFILLER_21_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1896_ gencon_inst.ALU_out\[1\] net68 net60 gencon_inst.mult_calc.out\[1\] VGND VGND
+ VPWR VPWR _1000_ sky130_fd_sc_hd__a22o_1
X_2517_ clknet_leaf_1_clk _0078_ net120 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_75_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2448_ clknet_leaf_4_clk _0036_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_2379_ input_ctrl_inst.col_index\[11\] _0513_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_54_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold8 gencon_inst.mult_calc.INn1\[1\] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__dlygate4sd3_1
X_1750_ gencon_inst.ALU_in1\[11\] gencon_inst.ALU_in2\[11\] net64 VGND VGND VPWR VPWR
+ _0939_ sky130_fd_sc_hd__mux2_1
XFILLER_30_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1681_ _0844_ _0889_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__xnor2_1
X_2164_ input_ctrl_inst.decoded_key\[0\] _1204_ _1205_ net83 VGND VGND VPWR VPWR _1206_
+ sky130_fd_sc_hd__o211a_1
X_2302_ _0473_ net202 VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__nor2_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2233_ _1044_ _0416_ _0430_ _0431_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__o31a_1
XFILLER_65_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2095_ input_ctrl_inst.debounce_cnt\[7\] _1147_ input_ctrl_inst.debounce_cnt\[8\]
+ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__a21oi_1
X_1879_ net192 gencon_inst.latched_keypad_input\[3\] _0961_ VGND VGND VPWR VPWR _0341_
+ sky130_fd_sc_hd__mux2_1
X_1948_ gencon_inst.operand2\[8\] net50 net33 net366 VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_43_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1733_ net316 _0930_ net110 VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__mux2_1
X_2782_ clknet_leaf_21_clk _0326_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[8\] sky130_fd_sc_hd__dfxtp_1
X_1802_ net168 _0969_ net41 VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__mux2_1
XFILLER_7_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1595_ net107 gencon_inst.add_calc.main.in2\[7\] VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__nand2_1
X_1664_ _0823_ _0824_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__nand2b_1
Xhold216 net11 VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 input_ctrl_inst.scan_timer\[10\] VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 gencon_inst.mult_calc.compCount.in2\[6\] VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 gencon_inst.mult_calc.compCount.in2\[9\] VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 gencon_inst.mult_calc.adderSave\[3\] VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2147_ input_ctrl_inst.decoded_key\[1\] net83 _1191_ VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__o21ai_1
X_2216_ _0402_ _0409_ _0414_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_64_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2078_ _1139_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__inv_2
XFILLER_53_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1380_ _0692_ _0693_ gencon_inst.mult_calc.out\[14\] net66 VGND VGND VPWR VPWR _0694_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2001_ gencon_inst.mult_calc.INn2\[5\] gencon_inst.mult_calc.INn2\[4\] gencon_inst.mult_calc.INn2\[7\]
+ gencon_inst.mult_calc.INn2\[6\] VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_61_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1716_ _0853_ _0918_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__xnor2_1
X_2696_ clknet_leaf_16_clk _0240_ net154 VGND VGND VPWR VPWR gencon_inst.ALU_out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2765_ clknet_leaf_16_clk _0309_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[7\] sky130_fd_sc_hd__dfxtp_1
X_2834_ clknet_leaf_26_clk _0374_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_1647_ _0781_ net32 _0860_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__and3_1
X_1578_ net108 gencon_inst.add_calc.main.in2\[11\] VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__or2_1
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2550_ clknet_leaf_2_clk net164 net123 VGND VGND VPWR VPWR input_ctrl_inst.RowSync\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_2481_ clknet_leaf_9_clk _0012_ net131 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1363_ gencon_inst.operand2\[9\] _0674_ gencon_inst.operand2\[10\] VGND VGND VPWR
+ VPWR _0681_ sky130_fd_sc_hd__a21o_1
X_1432_ net97 gencon_inst.mult_calc.adderSave\[11\] net336 net81 VGND VGND VPWR VPWR
+ _0182_ sky130_fd_sc_hd__a22o_1
X_1501_ _0727_ _0728_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__or2_1
X_1294_ gencon_inst.ALU_out\[12\] net69 net57 gencon_inst.mult_calc.out\[12\] _0565_
+ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_43_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2817_ clknet_leaf_6_clk gencon_inst.next_state\[0\] net134 VGND VGND VPWR VPWR gencon_inst.gencon_state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2748_ clknet_leaf_27_clk _0292_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_2679_ clknet_leaf_28_clk _0228_ net149 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Left_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1981_ input_ctrl_inst.input_control_state\[1\] input_ctrl_inst.input_control_state\[0\]
+ net92 VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__nand3b_4
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2602_ clknet_leaf_30_clk _0151_ net146 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_2533_ clknet_leaf_38_clk _0094_ net121 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1346_ gencon_inst.operand2\[6\] _0665_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__nor2_1
X_2464_ clknet_leaf_7_clk _0027_ net124 VGND VGND VPWR VPWR input_ctrl_inst.decoded_key\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_1415_ gencon_inst.mult_calc.out\[10\] net415 net105 VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__mux2_1
XFILLER_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2395_ net204 _0523_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__xnor2_1
X_1277_ gencon_inst.operand1\[7\] gencon_inst.operand1\[8\] gencon_inst.operand1\[9\]
+ _0598_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_31_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_22_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout131 net133 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_4
Xfanout120 net122 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_4
XFILLER_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout153 net155 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_4
Xfanout142 net145 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_30_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2180_ gencon_inst.operator_input\[2\] gencon_inst.operator_input\[1\] VGND VGND
+ VPWR VPWR _0383_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_48_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
X_1895_ _0999_ net376 net40 VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__mux2_1
X_1964_ gencon_inst.gencon_state\[3\] VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__inv_2
XFILLER_33_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2447_ clknet_leaf_3_clk _0035_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2516_ clknet_leaf_1_clk _0077_ net121 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1329_ gencon_inst.operand2\[3\] gencon_inst.latched_keypad_input\[3\] VGND VGND
+ VPWR VPWR _0654_ sky130_fd_sc_hd__nor2_1
X_2378_ input_ctrl_inst.col_index\[11\] _0513_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_54_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold9 gencon_inst.mult_calc.INn1\[10\] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1680_ _0811_ _0812_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__and2b_1
X_2301_ input_ctrl_inst.scan_timer\[16\] _0471_ net201 VGND VGND VPWR VPWR _0474_
+ sky130_fd_sc_hd__a21oi_1
X_2163_ input_ctrl_inst.decoded_key\[0\] input_ctrl_inst.decoded_key\[1\] VGND VGND
+ VPWR VPWR _1205_ sky130_fd_sc_hd__nand2_1
XFILLER_38_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_2_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
X_2232_ input_ctrl_inst.col_index\[24\] _0418_ _0416_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__or3b_1
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2094_ input_ctrl_inst.debounce_cnt\[7\] input_ctrl_inst.debounce_cnt\[8\] _1147_
+ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_16_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1878_ net282 gencon_inst.latched_keypad_input\[2\] _0961_ VGND VGND VPWR VPWR _0340_
+ sky130_fd_sc_hd__mux2_1
X_1947_ gencon_inst.operand2\[7\] net50 net33 net393 VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__a22o_1
XFILLER_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold217 gencon_inst.add_calc.main.GENERATE_ADDER\[5\].thingy.in1 VGND VGND VPWR VPWR
+ net377 sky130_fd_sc_hd__dlygate4sd3_1
X_1663_ net32 _0874_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__nand2_1
X_1732_ gencon_inst.ALU_in1\[2\] gencon_inst.ALU_in2\[2\] net62 VGND VGND VPWR VPWR
+ _0930_ sky130_fd_sc_hd__mux2_1
X_1801_ gencon_inst.operand2\[1\] gencon_inst.operand1\[1\] net76 VGND VGND VPWR VPWR
+ _0969_ sky130_fd_sc_hd__mux2_1
X_2781_ clknet_leaf_16_clk _0325_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[7\] sky130_fd_sc_hd__dfxtp_1
Xhold206 gencon_inst.mult_calc.INn2\[8\] VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_13_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1594_ net107 gencon_inst.add_calc.main.in2\[7\] VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__or2_1
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold239 gencon_inst.mult_calc.adderSave\[14\] VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold228 gencon_inst.mult_calc.compCount.in2\[12\] VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_64_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2077_ input_ctrl_inst.debounce_cnt\[1\] input_ctrl_inst.debounce_cnt\[0\] input_ctrl_inst.debounce_cnt\[3\]
+ input_ctrl_inst.debounce_cnt\[2\] VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__and4_1
X_2146_ input_ctrl_inst.col_index\[1\] _1055_ net82 VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__or3_1
X_2215_ input_ctrl_inst.col_index\[19\] _0411_ _0412_ _0413_ VGND VGND VPWR VPWR _0414_
+ sky130_fd_sc_hd__and4_1
XFILLER_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2000_ net96 net101 VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_18_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2833_ clknet_leaf_27_clk _0373_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_1646_ net114 gencon_inst.ALU_out\[1\] VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__or2_1
X_2695_ clknet_leaf_16_clk _0239_ net153 VGND VGND VPWR VPWR gencon_inst.ALU_out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1715_ _0787_ _0788_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__and2b_1
X_2764_ clknet_leaf_16_clk net223 VGND VGND VPWR VPWR gencon_inst.ALU_in2\[6\] sky130_fd_sc_hd__dfxtp_1
X_1577_ gencon_inst.add_calc.main.GENERATE_ADDER\[12\].thingy.in1 _0789_ _0790_ VGND
+ VGND VPWR VPWR _0792_ sky130_fd_sc_hd__nand3_1
X_2129_ input_ctrl_inst.debounce_cnt\[15\] net37 _1177_ _1178_ VGND VGND VPWR VPWR
+ _0014_ sky130_fd_sc_hd__a22o_1
XFILLER_54_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2480_ clknet_leaf_9_clk _0011_ net138 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1500_ _0718_ _0722_ _0719_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__o21a_1
XFILLER_9_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1293_ _0622_ _0623_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__nor2_1
X_1362_ gencon_inst.operand2\[10\] gencon_inst.operand2\[9\] _0674_ VGND VGND VPWR
+ VPWR _0680_ sky130_fd_sc_hd__nand3_1
X_1431_ net97 gencon_inst.mult_calc.adderSave\[10\] net329 net81 VGND VGND VPWR VPWR
+ _0181_ sky130_fd_sc_hd__a22o_1
XFILLER_63_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2816_ clknet_leaf_14_clk _0360_ net135 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_21_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1629_ _0815_ _0819_ _0842_ _0816_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__o31a_1
X_2747_ clknet_leaf_27_clk _0291_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_2678_ clknet_leaf_28_clk _0227_ net149 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1980_ input_ctrl_inst.input_control_state\[1\] input_ctrl_inst.input_control_state\[0\]
+ net92 VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_43_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2463_ clknet_leaf_2_clk net174 VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_2532_ clknet_leaf_38_clk _0093_ net121 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_2601_ clknet_leaf_30_clk _0150_ net146 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_21_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1276_ gencon_inst.operand1\[8\] net44 _0608_ _0610_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__o22a_1
X_1345_ gencon_inst.operand2\[6\] gencon_inst.operand2\[5\] gencon_inst.operand2\[4\]
+ _0658_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__and4_1
X_1414_ gencon_inst.mult_calc.out\[9\] net300 net105 VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__mux2_1
X_2394_ net284 _0521_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__xor2_1
XFILLER_51_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout154 net155 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__buf_2
Xfanout110 gencon_inst.add_calc.state\[2\] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_4
Xfanout132 net133 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__buf_2
Xfanout143 net145 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_4
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout121 net122 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_57_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1894_ gencon_inst.ALU_out\[0\] net68 net60 gencon_inst.mult_calc.out\[0\] _0996_
+ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__a221o_1
X_1963_ gencon_inst.gencon_state\[0\] VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__inv_2
X_2446_ clknet_leaf_3_clk _0034_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2515_ clknet_leaf_0_clk _0076_ net120 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_68_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1259_ gencon_inst.operand1\[5\] _0591_ _0592_ _0596_ VGND VGND VPWR VPWR _0597_
+ sky130_fd_sc_hd__o22a_1
X_1328_ gencon_inst.operand2\[3\] gencon_inst.latched_keypad_input\[3\] VGND VGND
+ VPWR VPWR _0653_ sky130_fd_sc_hd__and2_1
XFILLER_24_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2377_ _0512_ _0513_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__nor2_1
XFILLER_24_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2300_ input_ctrl_inst.scan_timer\[17\] input_ctrl_inst.scan_timer\[16\] _0471_ VGND
+ VGND VPWR VPWR _0473_ sky130_fd_sc_hd__and3_1
X_2231_ input_ctrl_inst.col_index\[25\] input_ctrl_inst.col_index\[27\] input_ctrl_inst.col_index\[26\]
+ _0428_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__nand4_1
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2093_ net35 _1149_ _1150_ net38 input_ctrl_inst.debounce_cnt\[7\] VGND VGND VPWR
+ VPWR _0024_ sky130_fd_sc_hd__a32o_1
XFILLER_53_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2162_ input_ctrl_inst.decoded_key\[3\] input_ctrl_inst.decoded_key\[2\] VGND VGND
+ VPWR VPWR _1204_ sky130_fd_sc_hd__nand2_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1877_ net271 gencon_inst.latched_keypad_input\[1\] _0961_ VGND VGND VPWR VPWR _0339_
+ sky130_fd_sc_hd__mux2_1
X_1946_ gencon_inst.operand2\[6\] net50 net33 net319 VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__a22o_1
XFILLER_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2429_ net423 net59 _0548_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__a21bo_1
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1800_ net180 _0968_ net41 VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__mux2_1
Xhold207 gencon_inst.add_calc.main.GENERATE_ADDER\[7\].thingy.in1 VGND VGND VPWR VPWR
+ net367 sky130_fd_sc_hd__dlygate4sd3_1
X_1662_ _0864_ _0866_ _0871_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__or3_1
X_1731_ net311 _0929_ net110 VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__mux2_1
X_2780_ clknet_leaf_16_clk _0324_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold229 input_ctrl_inst.scan_timer\[15\] VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 gencon_inst.mult_calc.compCount.in2\[2\] VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__dlygate4sd3_1
X_1593_ gencon_inst.add_calc.main.GENERATE_ADDER\[8\].thingy.in1 _0805_ _0806_ VGND
+ VGND VPWR VPWR _0808_ sky130_fd_sc_hd__nand3_1
X_2214_ input_ctrl_inst.col_index\[21\] input_ctrl_inst.col_index\[20\] input_ctrl_inst.col_index\[23\]
+ input_ctrl_inst.col_index\[22\] VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_64_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2076_ net36 _1137_ _1138_ net37 net448 VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__a32o_1
X_2145_ _1187_ _1190_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__nor2_1
XFILLER_19_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1929_ gencon_inst.operand1\[12\] _0378_ net60 gencon_inst.mult_calc.out\[12\] VGND
+ VGND VPWR VPWR _1022_ sky130_fd_sc_hd__a22o_1
XFILLER_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold90 gencon_inst.ALU_in2\[14\] VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_18_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2763_ clknet_leaf_16_clk _0307_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[5\] sky130_fd_sc_hd__dfxtp_1
X_2832_ clknet_leaf_27_clk _0372_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1645_ _0835_ _0859_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__xnor2_1
X_1576_ _0789_ _0790_ gencon_inst.add_calc.main.GENERATE_ADDER\[12\].thingy.in1 VGND
+ VGND VPWR VPWR _0791_ sky130_fd_sc_hd__a21oi_1
X_1714_ _0912_ _0915_ _0858_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__o21ai_1
X_2694_ clknet_leaf_16_clk _0238_ net153 VGND VGND VPWR VPWR gencon_inst.ALU_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2128_ input_ctrl_inst.debounce_cnt\[15\] _1171_ _1156_ VGND VGND VPWR VPWR _1178_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_34_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2059_ _1039_ _1084_ _1125_ VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__o21ai_1
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1430_ net97 net300 net406 net81 VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__a22o_1
X_1292_ gencon_inst.operand1\[12\] _0618_ net72 VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__o21ai_1
X_1361_ gencon_inst.operand2\[9\] net55 _0679_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__o21a_1
XFILLER_63_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2815_ clknet_leaf_22_clk _0359_ net157 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfrtp_1
X_2746_ clknet_leaf_27_clk _0290_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1628_ _0819_ _0842_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__nor2_1
X_2677_ clknet_leaf_26_clk _0226_ net150 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1559_ net399 net90 _0777_ net102 VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__a22o_1
XFILLER_54_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2600_ clknet_leaf_31_clk _0149_ net146 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2462_ clknet_leaf_2_clk _0050_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_1413_ gencon_inst.mult_calc.out\[8\] net391 net105 VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__mux2_1
XFILLER_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2531_ clknet_leaf_39_clk _0092_ net121 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_2393_ input_ctrl_inst.col_index\[17\] _0521_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__nand2_1
XFILLER_68_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1275_ gencon_inst.mult_calc.out\[8\] net57 net43 _0609_ VGND VGND VPWR VPWR _0610_
+ sky130_fd_sc_hd__a211o_1
X_1344_ gencon_inst.operand2\[5\] _0664_ _0666_ _0635_ VGND VGND VPWR VPWR _0127_
+ sky130_fd_sc_hd__o22a_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2729_ clknet_leaf_20_clk _0273_ net158 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[8\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
Xfanout111 gencon_inst.add_calc.state\[2\] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_2
Xfanout133 net138 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_4
Xfanout155 net160 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
Xfanout144 net145 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_2
Xfanout122 net130 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__buf_2
Xfanout100 gencon_inst.mult_calc.state\[3\] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1962_ net98 VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__inv_2
X_1893_ _0560_ net52 VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__nor2_1
XFILLER_68_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2445_ clknet_leaf_3_clk _0033_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2514_ clknet_leaf_1_clk _0075_ net123 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2376_ input_ctrl_inst.col_index\[9\] input_ctrl_inst.col_index\[10\] _0511_ VGND
+ VGND VPWR VPWR _0513_ sky130_fd_sc_hd__and3_1
XFILLER_68_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1258_ gencon_inst.operand1\[5\] _0559_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__nor2_1
X_1327_ _0646_ _0648_ _0647_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__a21boi_1
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_49_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_58_Left_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_67_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2230_ _0408_ _0415_ _0427_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__a21o_1
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2092_ input_ctrl_inst.debounce_cnt\[7\] _1147_ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__or2_1
XFILLER_38_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2161_ input_ctrl_inst.decoded_key\[3\] net82 _1187_ _1203_ VGND VGND VPWR VPWR _0030_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1945_ gencon_inst.operand2\[5\] net50 net33 net384 VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1876_ net299 gencon_inst.latched_keypad_input\[0\] _0961_ VGND VGND VPWR VPWR _0338_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2359_ _0444_ _0502_ _0501_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2428_ _0546_ _0547_ _0528_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__or3b_1
XFILLER_71_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1592_ _0805_ _0806_ gencon_inst.add_calc.main.GENERATE_ADDER\[8\].thingy.in1 VGND
+ VGND VPWR VPWR _0807_ sky130_fd_sc_hd__a21oi_1
X_1730_ gencon_inst.ALU_in1\[1\] gencon_inst.ALU_in2\[1\] net62 VGND VGND VPWR VPWR
+ _0929_ sky130_fd_sc_hd__mux2_1
X_1661_ _0873_ _0872_ net447 net85 VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__a2bb2o_1
Xhold219 gencon_inst.add_calc.main.GENERATE_ADDER\[12\].thingy.in1 VGND VGND VPWR
+ VPWR net379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold208 gencon_inst.add_calc.main.in2\[13\] VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__dlygate4sd3_1
X_2144_ input_ctrl_inst.decoded_key\[0\] net82 _1189_ VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__a21oi_1
X_2213_ input_ctrl_inst.col_index\[17\] input_ctrl_inst.col_index\[16\] input_ctrl_inst.col_index\[18\]
+ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_64_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2075_ input_ctrl_inst.debounce_cnt\[1\] input_ctrl_inst.debounce_cnt\[0\] input_ctrl_inst.debounce_cnt\[2\]
+ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__a21o_1
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1859_ gencon_inst.operand1\[3\] net224 net46 VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__mux2_1
X_1928_ _1020_ _1021_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__or2_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold80 _0362_ VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 gencon_inst.mult_calc.countSave\[1\] VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__dlygate4sd3_1
X_1713_ net422 _0916_ net115 VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__mux2_1
X_2762_ clknet_leaf_16_clk _0306_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[4\] sky130_fd_sc_hd__dfxtp_1
X_2831_ clknet_leaf_27_clk _0371_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1644_ gencon_inst.add_calc.main.GENERATE_ADDER\[1\].thingy.in1 _0833_ VGND VGND
+ VPWR VPWR _0859_ sky130_fd_sc_hd__xor2_1
X_2693_ clknet_leaf_17_clk _0237_ net153 VGND VGND VPWR VPWR gencon_inst.ALU_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1575_ net108 gencon_inst.add_calc.main.in2\[12\] VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__nand2_1
XFILLER_6_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2127_ net35 _1171_ input_ctrl_inst.debounce_cnt\[15\] VGND VGND VPWR VPWR _1177_
+ sky130_fd_sc_hd__a21o_1
XFILLER_25_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2058_ _1039_ _1084_ _1120_ _1124_ _1123_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__a221o_1
XFILLER_22_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1360_ gencon_inst.mult_calc.out\[9\] net67 _0678_ net74 _0635_ VGND VGND VPWR VPWR
+ _0679_ sky130_fd_sc_hd__a221o_1
X_1291_ gencon_inst.operand1\[12\] _0618_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__and2_1
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2814_ clknet_leaf_23_clk _0358_ net156 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfrtp_1
X_2745_ clknet_leaf_26_clk _0289_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_2676_ clknet_leaf_26_clk _0225_ net144 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_21_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1627_ _0823_ _0827_ _0839_ _0824_ _0820_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__o311a_1
X_1489_ gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in1
+ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__nor2_1
X_1558_ _0775_ _0776_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_34_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_60_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_25_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_26_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2530_ clknet_leaf_39_clk _0091_ net121 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1343_ _1211_ _0665_ net66 gencon_inst.mult_calc.out\[5\] VGND VGND VPWR VPWR _0666_
+ sky130_fd_sc_hd__a2bb2o_1
X_2461_ clknet_leaf_2_clk _0049_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_1412_ gencon_inst.mult_calc.out\[7\] net279 net105 VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__mux2_1
XFILLER_5_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2392_ _0521_ _0522_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__and2b_1
X_1274_ _1035_ gencon_inst.ALU_out\[8\] _0560_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_16_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
X_2728_ clknet_leaf_18_clk _0272_ net154 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[7\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2659_ clknet_leaf_33_clk _0208_ net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout112 gencon_inst.add_calc.state\[2\] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout134 net135 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_4
Xfanout156 net157 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_4
Xfanout123 net125 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_4
Xfanout145 net160 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_2
Xfanout101 gencon_inst.mult_calc.state\[3\] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_2
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1892_ _1035_ _0561_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__nor2_1
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1961_ input_ctrl_inst.RowSync\[2\] VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__inv_2
X_2513_ clknet_leaf_2_clk net4 net123 VGND VGND VPWR VPWR input_ctrl_inst.RowMid\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_68_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1326_ gencon_inst.operand2\[2\] _0651_ net54 VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_5_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
X_2444_ clknet_leaf_3_clk _0032_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2375_ input_ctrl_inst.col_index\[9\] _0511_ net429 VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__a21oi_1
XFILLER_64_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1257_ gencon_inst.ALU_out\[5\] net68 net56 gencon_inst.mult_calc.out\[5\] VGND VGND
+ VPWR VPWR _0595_ sky130_fd_sc_hd__a22o_1
XFILLER_59_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2160_ input_ctrl_inst.RowSync\[3\] _1197_ _1198_ _1202_ net83 VGND VGND VPWR VPWR
+ _1203_ sky130_fd_sc_hd__o311a_1
XFILLER_24_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2091_ input_ctrl_inst.debounce_cnt\[7\] _1147_ VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1875_ net215 _0384_ _0385_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__a21bo_1
X_1944_ gencon_inst.operand2\[4\] net50 net33 net355 VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2427_ input_ctrl_inst.col_index\[27\] _0544_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__and2_1
XFILLER_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1309_ gencon_inst.operand2\[0\] gencon_inst.latched_keypad_input\[0\] VGND VGND
+ VPWR VPWR _0637_ sky130_fd_sc_hd__or2_1
X_2289_ net411 _0464_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__nor2_1
X_2358_ net117 input_ctrl_inst.col_index\[1\] _1198_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__and3_1
XFILLER_71_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1591_ net107 gencon_inst.add_calc.main.in2\[8\] VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__nand2_1
X_1660_ net32 _0869_ _0871_ net85 VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__a31o_1
Xhold209 gencon_inst.ALU_finish VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_50_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2143_ input_ctrl_inst.col_index\[0\] net30 net83 VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__and3_1
X_2212_ _0397_ _0404_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_64_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2074_ input_ctrl_inst.debounce_cnt\[1\] input_ctrl_inst.debounce_cnt\[0\] input_ctrl_inst.debounce_cnt\[2\]
+ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__nand3_1
XFILLER_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1858_ gencon_inst.operand1\[2\] net207 net47 VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__mux2_1
X_1927_ net53 _0979_ net39 net13 VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__a22o_1
X_1789_ net277 net369 _0958_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__mux2_1
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold70 gencon_inst.ALU_in1\[12\] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 gencon_inst.ALU_in1\[14\] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 input_ctrl_inst.input_control_state\[0\] VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2830_ clknet_leaf_26_clk _0370_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2692_ clknet_leaf_12_clk _0236_ net137 VGND VGND VPWR VPWR gencon_inst.ALU_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1712_ _0913_ _0915_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__xnor2_1
X_1643_ _0784_ _0787_ _0854_ _0857_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__o31a_1
X_2761_ clknet_leaf_16_clk net261 VGND VGND VPWR VPWR gencon_inst.ALU_in2\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1 _1006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1574_ net108 gencon_inst.add_calc.main.in2\[12\] VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__or2_1
X_2126_ _1170_ _1172_ _1173_ _1176_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__a31o_1
XFILLER_39_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2057_ gencon_inst.mult_calc.compCount.in2\[12\] _1118_ _1122_ gencon_inst.mult_calc.compCount.in2\[13\]
+ VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_24_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1290_ gencon_inst.operand1\[11\] net45 _0620_ _0621_ VGND VGND VPWR VPWR _0118_
+ sky130_fd_sc_hd__o22a_1
XFILLER_36_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2813_ clknet_leaf_22_clk _0357_ net157 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfrtp_1
XFILLER_31_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1626_ _0823_ _0827_ _0839_ _0824_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__o31a_1
X_2744_ clknet_leaf_25_clk _0288_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2675_ clknet_leaf_34_clk _0224_ net144 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1557_ _0770_ _0772_ _0771_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__o21ba_1
X_1488_ net387 net91 _0717_ net103 VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__a22o_1
X_2109_ net37 _1161_ _1162_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_37_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2460_ clknet_leaf_3_clk _0048_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1273_ gencon_inst.operand1\[8\] _0602_ _0607_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__o21a_1
X_1342_ gencon_inst.operand2\[5\] gencon_inst.operand2\[4\] _0658_ VGND VGND VPWR
+ VPWR _0665_ sky130_fd_sc_hd__and3_1
X_1411_ gencon_inst.mult_calc.out\[6\] net440 net105 VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__mux2_1
XFILLER_5_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2391_ input_ctrl_inst.col_index\[15\] _0519_ input_ctrl_inst.col_index\[16\] VGND
+ VGND VPWR VPWR _0522_ sky130_fd_sc_hd__a21o_1
XFILLER_24_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2727_ clknet_leaf_18_clk _0271_ net154 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[6\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1609_ gencon_inst.add_calc.main.GENERATE_ADDER\[4\].thingy.in1 _0821_ _0822_ VGND
+ VGND VPWR VPWR _0824_ sky130_fd_sc_hd__nand3_1
Xfanout113 gencon_inst.add_calc.state\[2\] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_2
X_2589_ clknet_leaf_37_clk _0138_ net126 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2658_ clknet_leaf_32_clk _0207_ net140 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout102 net103 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__buf_2
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout157 net160 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_4
Xfanout135 net138 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_2
Xfanout124 net125 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
Xfanout146 net148 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_40_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1891_ _0561_ _0968_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__and2_1
X_1960_ input_ctrl_inst.debounce_cnt\[0\] VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__inv_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2443_ gencon_inst.gencon_state\[1\] _1035_ _1036_ _1037_ VGND VGND VPWR VPWR _0558_
+ sky130_fd_sc_hd__and4_1
X_2512_ clknet_leaf_2_clk net3 net123 VGND VGND VPWR VPWR input_ctrl_inst.RowMid\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1256_ gencon_inst.operand1\[4\] net44 _0593_ _0594_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__o22a_1
X_1325_ net73 _0649_ _0650_ net66 gencon_inst.mult_calc.out\[2\] VGND VGND VPWR VPWR
+ _0651_ sky130_fd_sc_hd__a32o_1
X_2374_ net394 _0511_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__xor2_1
XFILLER_64_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2090_ _1147_ _1148_ net433 net38 VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_38_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1874_ net270 _0385_ _0384_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__a21bo_1
X_1943_ gencon_inst.operand2\[3\] _0965_ net42 net265 VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_16_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2426_ input_ctrl_inst.col_index\[27\] _0544_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_67_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1239_ _0570_ _0572_ _0576_ _0578_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__o211a_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1308_ net73 _1213_ _0560_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__or3_1
X_2288_ input_ctrl_inst.scan_timer\[12\] _0464_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__and2_1
X_2357_ net116 _0496_ input_ctrl_inst.col_index\[3\] VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__a21oi_1
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1590_ net107 gencon_inst.add_calc.main.in2\[8\] VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__or2_1
XFILLER_50_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2073_ net36 _1135_ _1136_ net38 input_ctrl_inst.debounce_cnt\[1\] VGND VGND VPWR
+ VPWR _0018_ sky130_fd_sc_hd__a32o_1
X_2142_ _1051_ _1052_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__nand2_1
XFILLER_38_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2211_ net75 _0404_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_64_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1857_ gencon_inst.operand1\[1\] net272 net46 VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__mux2_1
X_1788_ net110 net114 VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__or2_1
X_1926_ gencon_inst.ALU_out\[11\] net69 net61 gencon_inst.mult_calc.out\[11\] VGND
+ VGND VPWR VPWR _1020_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_12_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2409_ input_ctrl_inst.col_index\[22\] net59 VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__nand2_1
XFILLER_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold71 gencon_inst.ALU_in2\[5\] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 gencon_inst.mult_calc.out\[15\] VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in1 VGND VGND VPWR
+ VPWR net220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 gencon_inst.mult_calc.countSave\[7\] VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__dlygate4sd3_1
X_2691_ clknet_leaf_12_clk _0235_ net137 VGND VGND VPWR VPWR gencon_inst.ALU_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1642_ _1045_ _0856_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__nor2_1
X_1711_ _0852_ _0914_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__xnor2_1
X_2760_ clknet_leaf_13_clk _0304_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_31_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_2 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1573_ gencon_inst.add_calc.main.GENERATE_ADDER\[13\].thingy.in1 _0785_ _0786_ VGND
+ VGND VPWR VPWR _0788_ sky130_fd_sc_hd__nand3_1
XFILLER_66_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2125_ input_ctrl_inst.debounce_cnt\[14\] _1047_ _1052_ net30 _1175_ VGND VGND VPWR
+ VPWR _1176_ sky130_fd_sc_hd__a41o_1
X_2056_ gencon_inst.mult_calc.compCount.in2\[13\] _1122_ VGND VGND VPWR VPWR _1123_
+ sky130_fd_sc_hd__nor2_1
X_1909_ net53 _0973_ net39 net22 VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__a22o_1
XFILLER_22_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2812_ clknet_leaf_27_clk _0356_ net151 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfrtp_1
X_2743_ clknet_leaf_25_clk _0287_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_1625_ _0827_ _0839_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__nor2_1
X_1556_ gencon_inst.mult_calc.main.GENERATE_ADDER\[14\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[14\].thingy.in1
+ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__xor2_1
X_2674_ clknet_leaf_34_clk _0223_ net142 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1487_ _0715_ _0716_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__xnor2_1
X_2108_ input_ctrl_inst.debounce_cnt\[10\] net35 _1155_ input_ctrl_inst.debounce_cnt\[11\]
+ VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_37_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2039_ gencon_inst.mult_calc.compCount.in2\[7\] _1105_ VGND VGND VPWR VPWR _1106_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_20_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_15_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1410_ gencon_inst.mult_calc.out\[5\] net289 net104 VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__mux2_1
X_1272_ _0559_ _0606_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__nor2_1
X_1341_ _0635_ _0663_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__nor2_1
X_2390_ input_ctrl_inst.col_index\[15\] input_ctrl_inst.col_index\[16\] _0519_ VGND
+ VGND VPWR VPWR _0521_ sky130_fd_sc_hd__and3_1
X_2726_ clknet_leaf_17_clk _0270_ net153 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[5\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1608_ _0821_ _0822_ gencon_inst.add_calc.main.GENERATE_ADDER\[4\].thingy.in1 VGND
+ VGND VPWR VPWR _0823_ sky130_fd_sc_hd__a21oi_1
Xfanout114 gencon_inst.add_calc.state\[1\] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_4
Xfanout136 net138 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_4
X_2588_ clknet_leaf_3_clk _0137_ net125 VGND VGND VPWR VPWR gencon_inst.read_input
+ sky130_fd_sc_hd__dfrtp_4
X_1539_ gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in1
+ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__nand2_1
Xfanout125 net130 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
X_2657_ clknet_leaf_33_clk _0206_ net140 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout103 gencon_inst.mult_calc.state\[2\] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_4
Xfanout147 net148 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_2
XFILLER_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout158 net160 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_4
XFILLER_50_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold190 gencon_inst.mult_calc.compCount.in2\[1\] VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1890_ _1036_ net10 _1215_ _0560_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__a31o_1
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2373_ _0510_ _0511_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__nor2_1
X_2442_ _0556_ _0557_ net417 VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__mux2_1
X_2511_ clknet_leaf_1_clk net2 net123 VGND VGND VPWR VPWR input_ctrl_inst.RowMid\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1255_ gencon_inst.ALU_out\[4\] net68 net56 gencon_inst.mult_calc.out\[4\] VGND VGND
+ VPWR VPWR _0594_ sky130_fd_sc_hd__a22o_1
X_1324_ _0647_ _0648_ _0646_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2709_ clknet_leaf_12_clk _0253_ net153 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1942_ gencon_inst.operand2\[2\] net51 net34 net308 VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_54_Left_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1873_ net302 gencon_inst.operator_input\[0\] _0386_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__mux2_1
X_2425_ net434 net58 _0545_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__a21bo_1
X_2356_ _0433_ _0497_ _0498_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_67_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1238_ _0576_ _0578_ _0570_ _0572_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__a211o_1
XFILLER_44_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1307_ _1213_ net66 VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__and2b_2
X_2287_ _0464_ _0465_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__and2b_1
XFILLER_52_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _0398_ _0399_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__nor2_1
X_2072_ input_ctrl_inst.debounce_cnt\[1\] input_ctrl_inst.debounce_cnt\[0\] VGND VGND
+ VPWR VPWR _1136_ sky130_fd_sc_hd__or2_1
X_2141_ _1051_ _1052_ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__and2_2
XFILLER_38_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1925_ net195 net39 _1019_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__a21o_1
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1787_ net373 _0957_ net112 VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__mux2_1
X_1856_ gencon_inst.operand1\[0\] net249 net46 VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__mux2_1
XFILLER_29_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2339_ net94 net235 net78 gencon_inst.mult_calc.count.GENERATE_ADDER\[6\].thingy.in1
+ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__a22o_1
X_2408_ input_ctrl_inst.col_index\[21\] net59 _0528_ _0533_ VGND VGND VPWR VPWR _0096_
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold50 gencon_inst.ALU_in1\[6\] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 gencon_inst.mult_calc.countSave\[12\] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 gencon_inst.mult_calc.countSave\[4\] VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 gencon_inst.mult_calc.countSave\[8\] VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 gencon_inst.mult_calc.countSave\[2\] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_61_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2690_ clknet_leaf_13_clk _0234_ net137 VGND VGND VPWR VPWR gencon_inst.ALU_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1710_ _0791_ _0792_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__nand2b_1
X_1572_ _0785_ _0786_ gencon_inst.add_calc.main.GENERATE_ADDER\[13\].thingy.in1 VGND
+ VGND VPWR VPWR _0787_ sky130_fd_sc_hd__a21oi_1
X_1641_ gencon_inst.add_calc.main.GENERATE_ADDER\[14\].thingy.in1 _0782_ _0783_ VGND
+ VGND VPWR VPWR _0856_ sky130_fd_sc_hd__and3_1
X_2124_ _1065_ _1174_ input_ctrl_inst.debounce_cnt\[14\] _1053_ VGND VGND VPWR VPWR
+ _1175_ sky130_fd_sc_hd__o211a_1
XFILLER_26_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2055_ _1082_ _1121_ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__nand2_1
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1839_ net118 net246 net46 VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__a21bo_1
X_1908_ gencon_inst.ALU_out\[5\] net70 net60 gencon_inst.mult_calc.out\[5\] VGND VGND
+ VPWR VPWR _1008_ sky130_fd_sc_hd__a22o_1
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_37_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_40_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_28_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_16_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2811_ clknet_leaf_22_clk _0355_ net156 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfrtp_1
X_2742_ clknet_leaf_35_clk _0286_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_1624_ _0831_ _0834_ _0836_ _0832_ _0828_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__o311a_1
X_1555_ net102 _0773_ _0774_ net285 net90 VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__a32o_1
X_2673_ clknet_leaf_33_clk _0222_ net140 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_19_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
X_2107_ _1156_ _1160_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__nor2_1
XFILLER_39_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1486_ _0707_ _0711_ _0708_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__o21ai_1
X_2038_ gencon_inst.mult_calc.count.GENERATE_ADDER\[7\].thingy.in1 _1077_ VGND VGND
+ VPWR VPWR _1105_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1340_ gencon_inst.mult_calc.out\[5\] net66 _0659_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__a21oi_1
X_1271_ gencon_inst.operand1\[7\] gencon_inst.operand1\[8\] _0598_ VGND VGND VPWR
+ VPWR _0606_ sky130_fd_sc_hd__and3_1
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2725_ clknet_leaf_17_clk _0269_ net153 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[4\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_8_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_42_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2656_ clknet_leaf_33_clk _0205_ net140 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1607_ net109 gencon_inst.add_calc.main.in2\[4\] VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__nand2_1
Xfanout115 gencon_inst.add_calc.state\[1\] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_2
Xfanout159 net160 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__buf_2
Xfanout137 net138 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__buf_2
X_2587_ clknet_leaf_11_clk _0005_ net136 VGND VGND VPWR VPWR gencon_inst.add_calc.next_finish
+ sky130_fd_sc_hd__dfrtp_1
X_1538_ gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in1
+ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__nor2_1
Xfanout126 net127 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_4
Xfanout148 net151 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_4
Xfanout104 gencon_inst.mult_calc.next_finish VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_4
X_1469_ gencon_inst.mult_calc.main.a0.in2 gencon_inst.mult_calc.main.a0.in1 VGND VGND
+ VPWR VPWR _0702_ sky130_fd_sc_hd__or2_1
XFILLER_63_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold180 gencon_inst.mult_calc.compCount.in2\[10\] VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 input_ctrl_inst.read_input_flag VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2510_ clknet_leaf_0_clk net1 net123 VGND VGND VPWR VPWR input_ctrl_inst.RowMid\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_1323_ _0646_ _0647_ _0648_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__nand3_1
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2372_ input_ctrl_inst.col_index\[8\] _0509_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__and2_1
X_2441_ _0451_ _0555_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__nand2b_1
X_1254_ gencon_inst.operand1\[4\] _0583_ _0586_ _0592_ VGND VGND VPWR VPWR _0593_
+ sky130_fd_sc_hd__o31a_1
X_2708_ clknet_leaf_12_clk _0252_ net137 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2639_ clknet_leaf_36_clk _0188_ net128 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1872_ net165 gencon_inst.read_input _0962_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__mux2_1
X_1941_ gencon_inst.operand2\[1\] _0965_ net41 net239 VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__o22a_1
XFILLER_69_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1306_ net73 _0560_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__nor2_1
X_2286_ input_ctrl_inst.scan_timer\[9\] input_ctrl_inst.scan_timer\[10\] _0461_ input_ctrl_inst.scan_timer\[11\]
+ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__a31o_1
X_2424_ _0527_ _0543_ _0544_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__or3_1
X_2355_ _0434_ _0499_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_67_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1237_ gencon_inst.operand1\[2\] gencon_inst.latched_keypad_input\[2\] VGND VGND
+ VPWR VPWR _0578_ sky130_fd_sc_hd__or2_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ net427 net37 net36 _1186_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__a22o_1
X_2071_ input_ctrl_inst.debounce_cnt\[1\] input_ctrl_inst.debounce_cnt\[0\] VGND VGND
+ VPWR VPWR _1135_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_29_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1855_ gencon_inst.operand2\[15\] net218 net46 VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__mux2_1
X_1924_ gencon_inst.operand2\[10\] _0387_ net69 gencon_inst.ALU_out\[10\] _1018_ VGND
+ VGND VPWR VPWR _1019_ sky130_fd_sc_hd__a221o_1
X_1786_ gencon_inst.ALU_in2\[14\] gencon_inst.ALU_in1\[14\] net63 VGND VGND VPWR VPWR
+ _0957_ sky130_fd_sc_hd__mux2_1
X_2269_ _0454_ _0455_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__and2b_1
X_2338_ net94 net237 net78 gencon_inst.mult_calc.count.GENERATE_ADDER\[5\].thingy.in1
+ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__a22o_1
X_2407_ input_ctrl_inst.col_index\[21\] _0530_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__xor2_1
XFILLER_71_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_73_Left_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold40 _0376_ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold51 gencon_inst.ALU_in2\[11\] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_61_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold62 gencon_inst.ALU_in2\[6\] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold84 _0064_ VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 _0068_ VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 gencon_inst.mult_calc.countSave\[13\] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1640_ _0787_ _0854_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__nor2_1
X_1571_ net107 gencon_inst.add_calc.main.in2\[13\] VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__nand2_1
XFILLER_6_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2123_ _1046_ net30 VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__nor2_1
XFILLER_39_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2054_ gencon_inst.mult_calc.count.GENERATE_ADDER\[13\].thingy.in1 _1081_ VGND VGND
+ VPWR VPWR _1121_ sky130_fd_sc_hd__or2_1
XFILLER_22_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1907_ _1006_ _1007_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__or2_1
XFILLER_41_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1838_ net184 _0987_ _0962_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__mux2_1
XFILLER_22_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1769_ net377 _0948_ net111 VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__mux2_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput30 net30 VGND VGND VPWR VPWR key_pressed sky130_fd_sc_hd__buf_2
Xoutput6 net6 VGND VGND VPWR VPWR ColOut[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_74_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2810_ clknet_leaf_22_clk _0354_ net156 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dfrtp_1
X_2741_ clknet_leaf_35_clk _0285_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_2672_ clknet_leaf_35_clk _0221_ net143 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1623_ _0831_ _0834_ _0836_ _0832_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__o31a_1
X_1485_ _0713_ _0714_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__nand2b_1
X_1554_ _0770_ _0771_ _0772_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__o21ai_1
.ends


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO outel8227
  CLASS BLOCK ;
  FOREIGN outel8227 ;
  ORIGIN 0.000 0.000 ;
  SIZE 208.785 BY 219.505 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 206.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 206.960 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 206.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 206.960 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END clk
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END cs
  PIN dataBusIn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 204.785 119.040 208.785 119.640 ;
    END
  END dataBusIn[0]
  PIN dataBusIn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 154.650 215.505 154.930 219.505 ;
    END
  END dataBusIn[1]
  PIN dataBusIn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 204.785 122.440 208.785 123.040 ;
    END
  END dataBusIn[2]
  PIN dataBusIn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END dataBusIn[3]
  PIN dataBusIn[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 204.785 132.640 208.785 133.240 ;
    END
  END dataBusIn[4]
  PIN dataBusIn[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 204.785 88.440 208.785 89.040 ;
    END
  END dataBusIn[5]
  PIN dataBusIn[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 204.785 136.040 208.785 136.640 ;
    END
  END dataBusIn[6]
  PIN dataBusIn[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 204.785 129.240 208.785 129.840 ;
    END
  END dataBusIn[7]
  PIN dataBusOut[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END dataBusOut[0]
  PIN dataBusOut[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END dataBusOut[1]
  PIN dataBusOut[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END dataBusOut[2]
  PIN dataBusOut[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END dataBusOut[3]
  PIN dataBusOut[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END dataBusOut[4]
  PIN dataBusOut[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END dataBusOut[5]
  PIN dataBusOut[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END dataBusOut[6]
  PIN dataBusOut[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END dataBusOut[7]
  PIN dataBusSelect
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END dataBusSelect
  PIN gpio[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END gpio[0]
  PIN gpio[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 119.230 215.505 119.510 219.505 ;
    END
  END gpio[10]
  PIN gpio[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 132.110 215.505 132.390 219.505 ;
    END
  END gpio[11]
  PIN gpio[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 122.450 215.505 122.730 219.505 ;
    END
  END gpio[12]
  PIN gpio[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 125.670 215.505 125.950 219.505 ;
    END
  END gpio[13]
  PIN gpio[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 141.770 215.505 142.050 219.505 ;
    END
  END gpio[14]
  PIN gpio[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 128.890 215.505 129.170 219.505 ;
    END
  END gpio[15]
  PIN gpio[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END gpio[16]
  PIN gpio[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END gpio[17]
  PIN gpio[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END gpio[18]
  PIN gpio[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END gpio[19]
  PIN gpio[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END gpio[1]
  PIN gpio[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END gpio[20]
  PIN gpio[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.741500 ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER met3 ;
        RECT 204.785 81.640 208.785 82.240 ;
    END
  END gpio[21]
  PIN gpio[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.431000 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END gpio[22]
  PIN gpio[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END gpio[23]
  PIN gpio[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END gpio[24]
  PIN gpio[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END gpio[25]
  PIN gpio[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END gpio[2]
  PIN gpio[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END gpio[3]
  PIN gpio[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END gpio[4]
  PIN gpio[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 35.510 215.505 35.790 219.505 ;
    END
  END gpio[5]
  PIN gpio[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END gpio[6]
  PIN gpio[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END gpio[7]
  PIN gpio[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 138.550 215.505 138.830 219.505 ;
    END
  END gpio[8]
  PIN gpio[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 135.330 215.505 135.610 219.505 ;
    END
  END gpio[9]
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 204.785 17.040 208.785 17.640 ;
    END
  END nrst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 203.050 206.805 ;
      LAYER li1 ;
        RECT 5.520 10.795 202.860 206.805 ;
      LAYER met1 ;
        RECT 4.210 10.640 202.860 206.960 ;
      LAYER met2 ;
        RECT 4.230 215.225 35.230 215.505 ;
        RECT 36.070 215.225 118.950 215.505 ;
        RECT 119.790 215.225 122.170 215.505 ;
        RECT 123.010 215.225 125.390 215.505 ;
        RECT 126.230 215.225 128.610 215.505 ;
        RECT 129.450 215.225 131.830 215.505 ;
        RECT 132.670 215.225 135.050 215.505 ;
        RECT 135.890 215.225 138.270 215.505 ;
        RECT 139.110 215.225 141.490 215.505 ;
        RECT 142.330 215.225 154.370 215.505 ;
        RECT 155.210 215.225 201.390 215.505 ;
        RECT 4.230 4.280 201.390 215.225 ;
        RECT 4.230 4.000 57.770 4.280 ;
        RECT 58.610 4.000 60.990 4.280 ;
        RECT 61.830 4.000 64.210 4.280 ;
        RECT 65.050 4.000 67.430 4.280 ;
        RECT 68.270 4.000 70.650 4.280 ;
        RECT 71.490 4.000 73.870 4.280 ;
        RECT 74.710 4.000 77.090 4.280 ;
        RECT 77.930 4.000 80.310 4.280 ;
        RECT 81.150 4.000 83.530 4.280 ;
        RECT 84.370 4.000 89.970 4.280 ;
        RECT 90.810 4.000 96.410 4.280 ;
        RECT 97.250 4.000 102.850 4.280 ;
        RECT 103.690 4.000 106.070 4.280 ;
        RECT 106.910 4.000 109.290 4.280 ;
        RECT 110.130 4.000 115.730 4.280 ;
        RECT 116.570 4.000 118.950 4.280 ;
        RECT 119.790 4.000 201.390 4.280 ;
      LAYER met3 ;
        RECT 3.990 194.840 204.785 206.885 ;
        RECT 4.400 193.440 204.785 194.840 ;
        RECT 3.990 181.240 204.785 193.440 ;
        RECT 4.400 179.840 204.785 181.240 ;
        RECT 3.990 174.440 204.785 179.840 ;
        RECT 4.400 173.040 204.785 174.440 ;
        RECT 3.990 171.040 204.785 173.040 ;
        RECT 4.400 169.640 204.785 171.040 ;
        RECT 3.990 167.640 204.785 169.640 ;
        RECT 4.400 166.240 204.785 167.640 ;
        RECT 3.990 164.240 204.785 166.240 ;
        RECT 4.400 162.840 204.785 164.240 ;
        RECT 3.990 157.440 204.785 162.840 ;
        RECT 4.400 156.040 204.785 157.440 ;
        RECT 3.990 154.040 204.785 156.040 ;
        RECT 4.400 152.640 204.785 154.040 ;
        RECT 3.990 150.640 204.785 152.640 ;
        RECT 4.400 149.240 204.785 150.640 ;
        RECT 3.990 137.040 204.785 149.240 ;
        RECT 3.990 135.640 204.385 137.040 ;
        RECT 3.990 133.640 204.785 135.640 ;
        RECT 3.990 132.240 204.385 133.640 ;
        RECT 3.990 130.240 204.785 132.240 ;
        RECT 3.990 128.840 204.385 130.240 ;
        RECT 3.990 123.440 204.785 128.840 ;
        RECT 3.990 122.040 204.385 123.440 ;
        RECT 3.990 120.040 204.785 122.040 ;
        RECT 3.990 118.640 204.385 120.040 ;
        RECT 3.990 89.440 204.785 118.640 ;
        RECT 3.990 88.040 204.385 89.440 ;
        RECT 3.990 82.640 204.785 88.040 ;
        RECT 3.990 81.240 204.385 82.640 ;
        RECT 3.990 55.440 204.785 81.240 ;
        RECT 4.400 54.040 204.785 55.440 ;
        RECT 3.990 18.040 204.785 54.040 ;
        RECT 3.990 16.640 204.385 18.040 ;
        RECT 3.990 10.715 204.785 16.640 ;
      LAYER met4 ;
        RECT 23.295 19.215 23.940 176.625 ;
        RECT 26.340 19.215 174.240 176.625 ;
        RECT 176.640 19.215 177.540 176.625 ;
        RECT 179.940 19.215 192.905 176.625 ;
  END
END outel8227
END LIBRARY


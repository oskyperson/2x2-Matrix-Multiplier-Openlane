* NGSPICE file created from outel8227.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

.subckt outel8227 VGND VPWR clk cs dataBusIn[0] dataBusIn[1] dataBusIn[2] dataBusIn[3]
+ dataBusIn[4] dataBusIn[5] dataBusIn[6] dataBusIn[7] dataBusOut[0] dataBusOut[1]
+ dataBusOut[2] dataBusOut[3] dataBusOut[4] dataBusOut[5] dataBusOut[6] dataBusOut[7]
+ dataBusSelect gpio[0] gpio[10] gpio[11] gpio[12] gpio[13] gpio[14] gpio[15] gpio[16]
+ gpio[17] gpio[18] gpio[19] gpio[1] gpio[20] gpio[21] gpio[22] gpio[23] gpio[24]
+ gpio[25] gpio[2] gpio[3] gpio[4] gpio[5] gpio[6] gpio[7] gpio[8] gpio[9] nrst
X_2106_ top8227.internalDataflow.addressLowBusModule.busInputs\[35\] _1277_ _1282_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[19\] VGND VGND VPWR VPWR
+ _0161_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2037_ _1245_ _1307_ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1606_ _0882_ _0885_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__or2_1
X_2724_ clknet_4_2_0_clk top8227.instructionLoader.interruptInjector.interruptRequest
+ net132 VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.irqSync.nextQ2
+ sky130_fd_sc_hd__dfrtp_1
X_2655_ _0284_ _0285_ _0288_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__nand3_1
XFILLER_0_13_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout138 net139 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_4
X_1537_ net2 net1 net62 VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__o21ai_2
Xfanout127 top8227.demux.state_machine.timeState\[0\] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_38_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout105 net107 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__buf_2
Xfanout116 top8227.demux.state_machine.timeState\[2\] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_4
X_1468_ net79 net76 VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__and2_2
X_2586_ _0241_ _0252_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__xor2_1
X_1399_ top8227.demux.state_machine.currentInstruction\[5\] top8227.demux.state_machine.currentInstruction\[4\]
+ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__nand2_2
XFILLER_0_64_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2440_ net25 _0437_ _0440_ _0455_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__or4_1
XFILLER_0_59_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2371_ _1286_ _0402_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_19_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_12_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2569_ _1237_ top8227.internalDataflow.accRegToDB\[7\] _0552_ VGND VGND VPWR VPWR
+ _0090_ sky130_fd_sc_hd__mux2_1
X_2707_ clknet_4_10_0_clk _0021_ net142 VGND VGND VPWR VPWR top8227.demux.state_machine.currentInstruction\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2638_ _0120_ _0566_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_53_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1871_ net31 _1139_ _1142_ VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1940_ _0724_ _0746_ _1062_ VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_16_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2423_ _0447_ _0450_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2354_ _0363_ _0385_ _0362_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__o21a_1
X_2285_ _0649_ net159 top8227.demux.nmi VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2070_ top8227.internalDataflow.addressHighBusModule.busInputs\[20\] _1227_ _1228_
+ net148 _1234_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_64_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1854_ _1126_ _1122_ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__and2b_1
X_1785_ top8227.branchBackward _1034_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__and2_1
X_1923_ _0751_ _0797_ net73 VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2406_ _0433_ _0434_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2337_ top8227.internalDataflow.addressLowBusModule.busInputs\[20\] net23 VGND VGND
+ VPWR VPWR _0369_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2268_ net117 net57 _0765_ _0318_ _0646_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__a311o_1
X_2199_ _0200_ _0209_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__xor2_2
XFILLER_0_62_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold52 top8227.internalDataflow.accRegToDB\[1\] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 top8227.internalDataflow.addressLowBusModule.busInputs\[33\] VGND VGND VPWR
+ VPWR net189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 top8227.internalDataflow.stackBusModule.busInputs\[46\] VGND VGND VPWR VPWR
+ net178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1570_ net2 _0853_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2053_ _1142_ _1319_ _1318_ _1143_ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__a2bb2o_1
X_2122_ net30 _0176_ _0170_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_29_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1906_ net53 _1158_ _1178_ _1148_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__a211o_1
X_1768_ _0684_ _0750_ net119 VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__o21a_1
X_1837_ net116 net64 _1015_ _1036_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__a211o_1
X_1699_ net29 _0826_ _0835_ _0976_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2740_ clknet_4_13_0_clk _0046_ net138 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[20\]
+ sky130_fd_sc_hd__dfrtp_2
X_1622_ net87 net80 net36 _0884_ _0889_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__a32o_1
X_2671_ net187 _0225_ _0637_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__mux2_1
X_1553_ _0843_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__inv_2
X_1484_ _0775_ _0777_ _0784_ net109 VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__o31a_1
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2036_ _1256_ _1253_ _1308_ VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__mux2_1
X_2105_ _1253_ _1256_ _0158_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_39_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_48_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2723_ clknet_4_8_0_clk net156 net141 VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.irqGenerated
+ sky130_fd_sc_hd__dfrtp_1
X_2585_ gpio[7] _0560_ _1286_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__a21o_1
X_1536_ net2 net61 VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__nand2_1
X_1605_ _0776_ net39 _0881_ _0884_ _0880_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2654_ _0291_ _0293_ _0286_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__a21oi_1
Xfanout128 top8227.demux.state_machine.currentAddress\[1\] VGND VGND VPWR VPWR net128
+ sky130_fd_sc_hd__clkbuf_4
Xfanout106 net107 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__buf_2
Xfanout139 net140 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1467_ _0765_ _0767_ net109 VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__o21a_1
Xfanout117 net118 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__buf_2
X_1398_ top8227.demux.state_machine.currentInstruction\[5\] top8227.demux.state_machine.currentInstruction\[4\]
+ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2019_ _1289_ _1290_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__nor2_2
XFILLER_0_60_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2370_ _1307_ _1334_ _0401_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_19_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2706_ clknet_4_11_0_clk _0020_ net142 VGND VGND VPWR VPWR top8227.demux.state_machine.currentInstruction\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2499_ _0504_ _0505_ net50 _0502_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__a211o_2
X_2568_ _1303_ top8227.internalDataflow.accRegToDB\[6\] _0552_ VGND VGND VPWR VPWR
+ _0089_ sky130_fd_sc_hd__mux2_1
X_1519_ top8227.demux.state_machine.currentAddress\[6\] _0810_ _0813_ _0817_ _0818_
+ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__a2111o_2
X_2637_ _0607_ top8227.internalDataflow.addressLowBusModule.busInputs\[28\] _0576_
+ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1870_ net31 _1139_ _1142_ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_43_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2422_ _0422_ _0448_ _0449_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__a21oi_1
X_2353_ _0366_ _0384_ _0365_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_24_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2284_ _0311_ _0326_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1999_ _1268_ _1270_ _1259_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_11_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_56_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1922_ _0671_ _0697_ _0768_ _0785_ _1194_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1784_ _1049_ _1052_ _1053_ _1056_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__a31o_1
X_1853_ _0665_ _1058_ _1125_ net59 VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__o31a_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2405_ top8227.internalDataflow.addressHighBusModule.busInputs\[18\] net26 _0423_
+ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__a21oi_1
X_2336_ _0366_ _0367_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2267_ _1062_ _1108_ net57 VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__o21a_1
X_2198_ _0240_ _0252_ _0239_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold42 top8227.demux.state_machine.currentAddress\[11\] VGND VGND VPWR VPWR net190
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 top8227.demux.state_machine.currentAddress\[3\] VGND VGND VPWR VPWR net179
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 top8227.internalDataflow.stackBusModule.busInputs\[47\] VGND VGND VPWR VPWR
+ net168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 top8227.internalDataflow.addressLowBusModule.busInputs\[24\] VGND VGND VPWR
+ VPWR net201 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_61_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2121_ _1144_ _0174_ _0175_ _1142_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__o22a_1
X_2052_ _1324_ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1905_ _0653_ _0712_ _1177_ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__or3b_1
X_1698_ net80 net75 net41 _0975_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__a31o_1
X_1767_ _0682_ net77 net78 net122 VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1836_ _1014_ _1059_ _1062_ _1108_ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__or4_1
X_2319_ net124 _0811_ _1020_ _0349_ _0350_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_67_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput10 net10 VGND VGND VPWR VPWR dataBusOut[0] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1552_ net148 net4 net3 net62 VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__o31a_1
X_1621_ net64 net39 _0827_ _0866_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2670_ _0752_ _0759_ _0636_ net60 VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__o31a_4
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1483_ _0656_ net78 _0779_ _0781_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__a211o_1
X_2104_ _0158_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2035_ _1128_ _1295_ _1300_ _1091_ VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1819_ _1091_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__inv_2
X_2799_ clknet_4_1_0_clk _0105_ net130 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2722_ clknet_4_2_0_clk net160 net132 VGND VGND VPWR VPWR top8227.demux.nmi sky130_fd_sc_hd__dfrtp_2
XFILLER_0_13_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2584_ gpio[6] _0560_ _1307_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__a21o_1
X_1535_ net2 net61 VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__and2_1
X_1604_ net29 _0883_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__and2_1
Xfanout107 top8227.demux.state_machine.timeState\[6\] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__buf_2
X_2653_ _0618_ _0621_ _0270_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__a21o_1
Xfanout129 net130 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_4
Xfanout118 net122 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
X_1466_ net90 _0766_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__and2_1
X_1397_ _0665_ _0670_ _0676_ _0681_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__o31a_1
XFILLER_0_49_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2018_ _1290_ VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2705_ clknet_4_12_0_clk _0026_ net138 VGND VGND VPWR VPWR top8227.branchForward
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_42_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2636_ _0605_ _0606_ _0270_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2498_ _0811_ _1018_ _1037_ _1050_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__a22oi_1
X_1518_ top8227.demux.state_machine.currentAddress\[12\] _0810_ VGND VGND VPWR VPWR
+ _0818_ sky130_fd_sc_hd__and2_1
X_2567_ _1327_ top8227.internalDataflow.accRegToDB\[5\] _0552_ VGND VGND VPWR VPWR
+ _0088_ sky130_fd_sc_hd__mux2_1
X_1449_ net80 _0717_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__and2_2
XFILLER_0_10_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2421_ top8227.internalDataflow.addressHighBusModule.busInputs\[19\] top8227.internalDataflow.addressHighBusModule.busInputs\[17\]
+ top8227.internalDataflow.addressHighBusModule.busInputs\[18\] top8227.internalDataflow.addressHighBusModule.busInputs\[16\]
+ net26 VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__o41a_1
X_2352_ _0369_ _0383_ _0368_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__o21a_1
X_2283_ net49 _0825_ top8227.demux.setInterruptFlag VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_10_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1998_ _1268_ _1270_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__and2_1
X_2619_ _0257_ _0565_ _0567_ _0187_ net32 VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_7_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1852_ _1029_ _1044_ _1123_ _1124_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1921_ _0708_ _0742_ _0795_ net73 VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__o31a_1
X_1783_ top8227.branchForward _1034_ _1055_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2404_ top8227.internalDataflow.addressHighBusModule.busInputs\[19\] net25 VGND VGND
+ VPWR VPWR _0433_ sky130_fd_sc_hd__xor2_1
X_2335_ top8227.internalDataflow.addressLowBusModule.busInputs\[21\] net23 VGND VGND
+ VPWR VPWR _0367_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2266_ _0268_ _0269_ _0316_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__and3_1
X_2197_ net49 _0251_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold54 top8227.demux.state_machine.currentAddress\[5\] VGND VGND VPWR VPWR net202
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 top8227.internalDataflow.addressLowBusModule.busInputs\[32\] VGND VGND VPWR
+ VPWR net191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 top8227.internalDataflow.stackBusModule.busInputs\[44\] VGND VGND VPWR VPWR
+ net169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 net12 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 top8227.pulse_slower.nextEnableState\[1\] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2120_ top8227.internalDataflow.addressHighBusModule.busInputs\[18\] _1227_ _1228_
+ net3 _1234_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__a221oi_2
X_2051_ _1320_ _1321_ _1323_ _1127_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1904_ _1026_ _1044_ _1176_ _1175_ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__o31a_1
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1835_ net77 net74 net116 net88 VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__o211a_1
X_1697_ _0700_ net75 net41 _0827_ _0862_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__a32o_1
XFILLER_0_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1766_ _0685_ _0769_ _0797_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__or3_1
XFILLER_0_57_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2318_ top8227.demux.state_machine.currentAddress\[6\] _1037_ VGND VGND VPWR VPWR
+ _0350_ sky130_fd_sc_hd__and2_1
X_2249_ net119 _0792_ _1150_ _1155_ _0302_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_67_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_10_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
Xoutput11 net11 VGND VGND VPWR VPWR dataBusOut[1] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1551_ net54 _0804_ _0830_ _0841_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__and4_1
X_1620_ _0886_ _0891_ _0899_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__or3_1
X_1482_ _0700_ net76 VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__and2_1
X_2103_ _1092_ _0150_ _0155_ _1128_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__o22a_2
XFILLER_0_27_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2034_ _1280_ _1306_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__or2_2
XFILLER_0_43_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1818_ _1089_ _1090_ net50 _1088_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_4_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2798_ clknet_4_0_0_clk _0104_ net130 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1749_ _0806_ _0811_ _1021_ net67 VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__a211o_1
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2721_ clknet_4_2_0_clk _0031_ net132 VGND VGND VPWR VPWR top8227.demux.setInterruptFlag
+ sky130_fd_sc_hd__dfrtp_1
X_2652_ _1313_ _0563_ _0619_ _0620_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__a211o_1
X_2583_ gpio[5] _0560_ _1334_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__a21o_1
X_1534_ net147 net29 _0826_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__and3_2
X_1603_ net147 net7 net62 net146 VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__and4b_2
Xfanout119 net120 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__buf_2
XFILLER_0_22_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout108 net110 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__buf_2
X_1465_ net99 net104 net93 net96 VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__and4_1
X_2017_ _1238_ _1288_ VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__and2_1
X_1396_ _0686_ _0691_ _0694_ _0697_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__or4_1
XFILLER_0_64_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2635_ _0146_ _0282_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__xnor2_1
X_2704_ clknet_4_11_0_clk _0019_ net141 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2497_ _0805_ _0503_ _1260_ net71 VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__o211a_1
X_1517_ net126 top8227.demux.state_machine.currentAddress\[5\] _0814_ _0816_ _0815_
+ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__a221o_4
X_2566_ _0133_ top8227.internalDataflow.accRegToDB\[4\] _0552_ VGND VGND VPWR VPWR
+ _0087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1448_ _0745_ _0746_ _0747_ _0748_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__or4_1
XFILLER_0_65_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1379_ top8227.demux.reset _0679_ net84 net86 VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_2_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2420_ _0420_ _0433_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout90 net91 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_2
XFILLER_0_10_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2351_ _0372_ _0382_ _0371_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__o21a_1
X_2282_ gpio[20] net153 net49 VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1997_ net67 _0653_ _0712_ _1269_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_15_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2549_ _0402_ _0539_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2618_ net28 _0157_ _0272_ _0590_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_7_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1920_ _1185_ _1192_ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__nand2_1
X_1851_ net120 net79 net76 VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__and3_1
X_2403_ net19 _0425_ _0426_ _0432_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__o211a_1
X_1782_ net63 _1037_ _1054_ _1032_ _1036_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2334_ top8227.internalDataflow.addressLowBusModule.busInputs\[21\] net23 VGND VGND
+ VPWR VPWR _0366_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2196_ _0242_ _0244_ _0250_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__a21oi_1
X_2265_ _1289_ _1290_ _0315_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold22 top8227.internalDataflow.stackBusModule.busInputs\[40\] VGND VGND VPWR VPWR
+ net170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold11 top8227.instructionLoader.interruptInjector.nmiGeneratedFF.synchronizedNMI
+ VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 top8227.branchBackward VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 top8227.internalDataflow.stackBusModule.busInputs\[35\] VGND VGND VPWR VPWR
+ net181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2050_ _1132_ _1322_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1834_ top8227.demux.state_machine.currentAddress\[12\] top8227.demux.state_machine.currentAddress\[6\]
+ _1018_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1765_ net66 _0809_ _1037_ net63 _1036_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__a221o_1
X_1903_ _0781_ _0796_ net121 VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1696_ _0887_ _0908_ _0850_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2317_ net112 top8227.demux.state_machine.currentAddress\[7\] net81 _0720_ VGND VGND
+ VPWR VPWR _0349_ sky130_fd_sc_hd__and4_1
X_2179_ net105 _0716_ _1036_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__or3b_1
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2248_ _0747_ _1073_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput12 net12 VGND VGND VPWR VPWR dataBusOut[2] sky130_fd_sc_hd__buf_2
X_1550_ _0832_ _0838_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1481_ _0662_ _0701_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__nor2_1
X_2102_ _0152_ _0156_ net30 VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__mux2_2
X_2033_ net7 _1281_ _1282_ top8227.internalDataflow.addressLowBusModule.busInputs\[22\]
+ _1305_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1748_ net128 _0809_ _0816_ net124 _1020_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2797_ clknet_4_1_0_clk _0103_ net129 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1817_ net101 _0692_ net78 _0817_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__nand4_4
X_1679_ net78 _0717_ net37 _0863_ _0897_ VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__a32o_1
XFILLER_0_67_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2582_ gpio[4] _0560_ _0140_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1602_ _0767_ net39 _0827_ _0881_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__a22o_1
X_2720_ clknet_4_2_0_clk _0030_ net132 VGND VGND VPWR VPWR top8227.negEdgeDetector.q1
+ sky130_fd_sc_hd__dfrtp_1
X_2651_ _1239_ _0272_ _0567_ _1312_ net32 VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__a221o_1
X_1533_ _0648_ net7 net61 VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__and3_2
Xfanout109 net110 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_2
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1464_ _0673_ _0693_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__nor2_2
X_1395_ _0669_ _0696_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__nor2_2
XFILLER_0_49_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2016_ _1238_ _1288_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1516_ top8227.demux.state_machine.currentAddress\[11\] top8227.demux.state_machine.currentAddress\[3\]
+ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__or2_2
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2565_ _0157_ top8227.internalDataflow.accRegToDB\[3\] _0552_ VGND VGND VPWR VPWR
+ _0086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2634_ net32 _0262_ _0602_ _0604_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__a31o_1
X_2703_ clknet_4_8_0_clk _0018_ net141 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2496_ net125 top8227.demux.state_machine.currentAddress\[5\] top8227.demux.state_machine.currentAddress\[7\]
+ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__a21oi_1
X_1378_ net106 _0678_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1447_ net116 net88 _0661_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout80 net81 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_2
Xfanout91 _0654_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2350_ _0375_ _0381_ _0374_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__o21a_1
X_2281_ top8227.demux.nmi net49 _0325_ _0311_ net174 VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__o32a_1
XFILLER_0_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1996_ top8227.demux.state_machine.currentAddress\[5\] net128 net125 VGND VGND VPWR
+ VPWR _1269_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_50_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2548_ _1306_ _0392_ net23 VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2617_ _0256_ _0564_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_7_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2479_ net170 _0225_ _0494_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload0 clknet_4_0_0_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__inv_6
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1781_ net123 _0787_ _1026_ _1041_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_12_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1850_ net121 _0657_ net79 VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__and3_2
X_2333_ _0363_ _0364_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__nor2_1
X_2402_ _0428_ _0430_ _0431_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2195_ top8227.PSRCurrentValue\[0\] net68 _0247_ _0249_ VGND VGND VPWR VPWR _0250_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2264_ _1312_ _0265_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1979_ _0735_ _1034_ _1249_ _1251_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold45 top8227.internalDataflow.addressLowBusModule.busInputs\[38\] VGND VGND VPWR
+ VPWR net193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 top8227.internalDataflow.stackBusModule.busInputs\[36\] VGND VGND VPWR VPWR
+ net171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 top8227.internalDataflow.stackBusModule.busInputs\[37\] VGND VGND VPWR VPWR
+ net182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 _0032_ VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1902_ _0695_ net78 _0817_ _1174_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1833_ net59 _1097_ _1105_ _0712_ _0653_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__a2111o_1
X_1764_ net123 net106 _0678_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__or3_2
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2316_ _0344_ _0347_ net60 VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__o21a_1
X_1695_ _0663_ net38 _0889_ _0909_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__a22o_1
X_2178_ net1 _1281_ _1284_ top8227.internalDataflow.addressLowBusModule.busInputs\[24\]
+ _0232_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2247_ _1017_ _0295_ _0300_ _0301_ VGND VGND VPWR VPWR top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[0\]
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_23_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput13 net13 VGND VGND VPWR VPWR dataBusOut[3] sky130_fd_sc_hd__buf_2
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1480_ _0674_ net78 VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2101_ _1127_ _0155_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__nor2_1
X_2032_ top8227.internalDataflow.addressLowBusModule.busInputs\[38\] _1277_ _1284_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[30\] VGND VGND VPWR VPWR
+ _1305_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1747_ net124 top8227.demux.state_machine.currentAddress\[7\] VGND VGND VPWR VPWR
+ _1020_ sky130_fd_sc_hd__and2_1
X_1816_ top8227.demux.state_machine.currentAddress\[12\] _0814_ net67 VGND VGND VPWR
+ VPWR _1089_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1678_ _0750_ net35 _0889_ _0956_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_15_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2796_ clknet_4_1_0_clk _0102_ net130 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2581_ gpio[3] _0560_ _0163_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__a21o_1
X_1601_ net5 _0830_ _0839_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__and3_2
XFILLER_0_22_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1532_ top8227.instructionLoader.interruptInjector.resetDetected _0824_ VGND VGND
+ VPWR VPWR _0825_ sky130_fd_sc_hd__and2b_2
XFILLER_0_10_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2650_ _1314_ _0566_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__nor2_1
X_1463_ _0758_ _0763_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__or2_1
X_1394_ net92 net95 net98 net102 VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_54_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2015_ _1257_ _1287_ _1246_ VGND VGND VPWR VPWR _1288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2779_ clknet_4_6_0_clk _0085_ net134 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2702_ clknet_4_11_0_clk _0017_ net142 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_1515_ net125 net113 top8227.demux.state_machine.currentAddress\[7\] VGND VGND VPWR
+ VPWR _0815_ sky130_fd_sc_hd__and3b_1
X_2564_ _0177_ top8227.internalDataflow.accRegToDB\[2\] _0552_ VGND VGND VPWR VPWR
+ _0085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2495_ _0501_ _1274_ _0497_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__and3b_1
X_2633_ _0145_ _0565_ _0567_ _0143_ _0603_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1377_ net115 net112 net105 VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__nor3_1
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1446_ net108 net88 _0695_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout70 net72 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_54_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout81 net82 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_2
Xfanout92 net94 VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_63_Left_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2280_ _0649_ _0324_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1995_ _0653_ _0712_ _1267_ VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__or3_2
XFILLER_0_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2616_ _0587_ _0588_ _0261_ _0280_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__a211o_1
X_2547_ _1307_ _0392_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2478_ net48 _0493_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_7_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1429_ top8227.PSRCurrentValue\[6\] net83 _0674_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_66_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload1 clknet_4_1_0_clk VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__inv_6
XPHY_EDGE_ROW_3_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1780_ _1018_ _1050_ _1020_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_12_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2332_ top8227.internalDataflow.addressLowBusModule.busInputs\[22\] net23 VGND VGND
+ VPWR VPWR _0364_ sky130_fd_sc_hd__nor2_1
X_2401_ _0428_ _0430_ net46 VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2194_ top8227.freeCarry net70 _0248_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2263_ top8227.PSRCurrentValue\[3\] _0298_ _0313_ _0314_ _0312_ VGND VGND VPWR VPWR
+ top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[3\] sky130_fd_sc_hd__a311o_1
XFILLER_0_47_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1978_ _1028_ _1123_ _1247_ _1250_ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold46 top8227.internalDataflow.addressLowBusModule.busInputs\[37\] VGND VGND VPWR
+ VPWR net194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 net16 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 net11 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 net13 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1901_ net128 _0814_ _1173_ net126 net68 VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__a221o_1
X_1832_ _1100_ _1104_ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1763_ top8227.demux.state_machine.timeState\[1\] net86 net84 VGND VGND VPWR VPWR
+ _1036_ sky130_fd_sc_hd__and3_2
X_1694_ _0771_ net35 _0836_ _0956_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2315_ _0338_ _0346_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__nand2_1
X_2246_ _0228_ _0298_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__nor2_1
X_2177_ top8227.internalDataflow.addressLowBusModule.busInputs\[16\] _1271_ _1278_
+ _1277_ top8227.internalDataflow.addressLowBusModule.busInputs\[32\] VGND VGND VPWR
+ VPWR _0232_ sky130_fd_sc_hd__a32o_1
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput14 net14 VGND VGND VPWR VPWR dataBusOut[4] sky130_fd_sc_hd__buf_2
XFILLER_0_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2100_ top8227.internalDataflow.addressLowBusModule.busInputs\[19\] _1129_ _0154_
+ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2031_ net28 _1303_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2795_ clknet_4_4_0_clk _0101_ net129 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_1815_ _1079_ _1080_ _1087_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__nor3_2
XTAP_TAPCELL_ROW_20_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1746_ top8227.demux.state_machine.currentAddress\[6\] _1018_ VGND VGND VPWR VPWR
+ _1019_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1677_ net44 _0938_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2229_ _0118_ _0283_ _1314_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2580_ gpio[2] _0560_ _0185_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__a21o_1
X_1600_ _0875_ _0878_ _0879_ _0867_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__a211o_1
X_1462_ _0759_ _0760_ _0761_ _0762_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1531_ top8227.demux.nmi top8227.instructionLoader.interruptInjector.irqGenerated
+ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__nor2_2
X_1393_ net94 net97 net100 net104 VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_70_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2014_ _1286_ VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2778_ clknet_4_6_0_clk _0084_ net135 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1729_ _0943_ _0979_ _1002_ _0830_ _1003_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2632_ _1328_ _0273_ _0564_ _0144_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2701_ clknet_4_11_0_clk _0016_ net141 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1514_ net126 net113 VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__and2b_2
X_2563_ _0199_ net200 _0552_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__mux2_1
X_2494_ net71 _0758_ _0498_ _0500_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1445_ net108 net83 net74 VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__and3_1
X_1376_ net114 net111 VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__or2_2
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout71 net72 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_2
XFILLER_0_51_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout60 _0715_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_4
Xfanout93 net94 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_1
Xfanout82 _0672_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_59_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1994_ _1034_ _1266_ _1261_ _1224_ VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_35_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2615_ _0277_ _0586_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__nand2_1
X_2546_ _1334_ _0401_ _1307_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2477_ net127 _0492_ _1197_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_7_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1428_ _0645_ _0669_ net76 VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_66_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1359_ net98 net102 net92 net95 VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__nor4b_1
Xclkload2 clknet_4_2_0_clk VGND VGND VPWR VPWR clkload2/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2400_ _0174_ _0396_ _0429_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2331_ top8227.internalDataflow.addressLowBusModule.busInputs\[22\] net23 VGND VGND
+ VPWR VPWR _0363_ sky130_fd_sc_hd__and2_1
X_2262_ _0313_ _0297_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2193_ net115 top8227.demux.state_machine.currentAddress\[1\] _0805_ _0811_ _0814_
+ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1977_ net64 _0808_ _1029_ _1036_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__a211o_1
XFILLER_0_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2529_ net47 _0383_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__nor2_1
Xhold47 top8227.internalDataflow.addressLowBusModule.busInputs\[34\] VGND VGND VPWR
+ VPWR net195 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 top8227.internalDataflow.stackBusModule.busInputs\[42\] VGND VGND VPWR VPWR
+ net173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 top8227.internalDataflow.stackBusModule.busInputs\[43\] VGND VGND VPWR VPWR
+ net184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 net14 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1900_ top8227.demux.state_machine.currentAddress\[3\] top8227.demux.state_machine.currentAddress\[10\]
+ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__or2_1
X_1831_ _1101_ _1103_ net67 VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1762_ net66 _0809_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1693_ _0925_ _0971_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__or2_1
X_2314_ _1198_ _0345_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__nor2_1
X_2176_ _0226_ _0227_ _1253_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__a21boi_1
X_2245_ _0299_ _0297_ _0296_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput15 net15 VGND VGND VPWR VPWR dataBusOut[5] sky130_fd_sc_hd__buf_2
XFILLER_0_66_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2030_ net31 _1302_ _1296_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_27_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1745_ _0807_ _0814_ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__nor2_1
X_1814_ net118 _0787_ _1081_ _1082_ _1086_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_17_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2794_ clknet_4_1_0_clk _0100_ net129 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1676_ _0742_ net37 net21 _0883_ _0954_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2159_ _0211_ _0212_ _0213_ _1184_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2228_ _0263_ _0281_ _0120_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1461_ _0674_ _0755_ net111 net90 VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__o211a_1
X_1530_ net107 net49 _0820_ net116 VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__a22o_1
X_1392_ _0655_ _0693_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__nor2_4
X_2013_ _1280_ _1285_ VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__or2_4
XFILLER_0_38_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1728_ _0882_ _0888_ _0894_ _0901_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__or4_1
X_2777_ clknet_4_3_0_clk _0083_ net133 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1659_ _0684_ net40 _0874_ _0938_ _0937_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2562_ _0225_ top8227.internalDataflow.accRegToDB\[0\] _0552_ VGND VGND VPWR VPWR
+ _0083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2631_ _0145_ _0261_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2700_ clknet_4_8_0_clk _0015_ net141 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1375_ net115 net112 VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1513_ net115 _0805_ _0811_ _0810_ net128 VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__a32o_1
X_2493_ net106 _0667_ _0675_ _0499_ _1205_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__a221o_1
X_1444_ net108 net79 _0705_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout72 _0651_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_2
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout61 _0825_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_2
Xfanout50 net52 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_4
XFILLER_0_36_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout83 net84 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
Xfanout94 top8227.demux.state_machine.currentInstruction\[3\] VGND VGND VPWR VPWR
+ net94 sky130_fd_sc_hd__buf_2
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1993_ _1262_ _1264_ _1265_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2545_ _0385_ _0537_ net19 VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_42_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2614_ _0277_ _0586_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__or2_1
X_2476_ net80 _0766_ _0782_ _0783_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__a211o_1
X_1427_ top8227.PSRCurrentValue\[7\] _0669_ net77 VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__or3b_1
X_1358_ net100 net103 VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_66_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload3 clknet_4_3_0_clk VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__inv_6
XFILLER_0_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2330_ _0360_ _0361_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__nor2_1
X_2261_ _0756_ _0776_ _1240_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__o21bai_2
X_2192_ _1015_ _0246_ _0245_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__or3b_1
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1976_ _1042_ _1059_ _1063_ _1248_ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2528_ top8227.internalDataflow.addressLowBusModule.busInputs\[19\] _0523_ net20
+ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__mux2_1
X_2459_ net25 _0478_ _0466_ _0465_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__a211oi_1
Xhold48 top8227.internalDataflow.addressLowBusModule.busInputs\[39\] VGND VGND VPWR
+ VPWR net196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 top8227.internalDataflow.stackBusModule.busInputs\[41\] VGND VGND VPWR VPWR
+ net163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 top8227.internalDataflow.stackBusModule.busInputs\[38\] VGND VGND VPWR VPWR
+ net185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 top8227.instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning VGND
+ VGND VPWR VPWR net174 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1761_ _0732_ _0733_ net111 VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1830_ net120 _0663_ _1040_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2313_ _0759_ _0760_ _1203_ _1204_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1692_ _0960_ _0965_ _0969_ _0970_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_69_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2175_ _1256_ _0226_ _0227_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__and3_1
X_2244_ _1017_ _0298_ top8227.PSRCurrentValue\[0\] VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__and3b_1
XFILLER_0_28_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1959_ net65 _0787_ net111 VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput16 net16 VGND VGND VPWR VPWR dataBusOut[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_39_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1813_ net72 _0747_ _1083_ _1085_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__or4b_1
X_2793_ clknet_4_3_0_clk _0099_ net132 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_1744_ _1012_ _1013_ _1014_ _1016_ net58 VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__o41a_1
XFILLER_0_68_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1675_ _0707_ net40 _0874_ _0887_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2158_ top8227.internalDataflow.stackBusModule.busInputs\[40\] _1186_ _1188_ top8227.internalDataflow.addressLowBusModule.busInputs\[32\]
+ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__a22oi_1
X_2089_ _0141_ _0142_ _0134_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2227_ _0261_ _0280_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_48_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1460_ net112 net84 _0755_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__and3_1
X_1391_ net99 net93 net96 net104 VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__or4b_4
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2012_ net146 _1281_ _1284_ top8227.internalDataflow.addressLowBusModule.busInputs\[31\]
+ _1283_ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2776_ clknet_4_7_0_clk _0082_ net137 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_1727_ _0856_ _0917_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__and2b_1
X_1658_ _0887_ _0914_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__nor2_2
X_1589_ net29 _0852_ _0866_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1512_ net115 _0805_ _0811_ _0810_ net128 VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__a32oi_4
X_2492_ net112 net105 _1201_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__or3_1
X_2561_ _0302_ _0550_ _0551_ net60 VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__o31ai_4
X_2630_ _0597_ _0598_ _0601_ _0576_ top8227.internalDataflow.addressLowBusModule.busInputs\[27\]
+ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__a32o_1
X_1443_ _0668_ net74 VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__and2_1
X_1374_ _0671_ net80 _0674_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2759_ clknet_4_4_0_clk _0065_ net130 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout73 _0806_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_4
Xfanout62 _0825_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_2
Xfanout40 net43 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_2
Xfanout51 net52 VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_1_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout84 _0668_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_2
Xfanout95 top8227.demux.state_machine.currentInstruction\[2\] VGND VGND VPWR VPWR
+ net95 sky130_fd_sc_hd__buf_2
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1992_ net114 net65 _0787_ net111 net70 VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload10 clknet_4_11_0_clk VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__inv_6
X_2544_ _0365_ _0366_ _0384_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__nor3_1
X_2475_ net196 _1237_ _0491_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__mux2_1
X_2613_ _1256_ _0245_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_50_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1426_ top8227.PSRCurrentValue\[0\] _0657_ net84 VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__and3_1
X_1357_ _0655_ _0658_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__nor2_2
Xclkload4 clknet_4_5_0_clk VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_33_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2260_ _0158_ _0298_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__nor2_1
X_2191_ net77 net75 net119 net78 VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_63_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1975_ net120 net107 net63 _1124_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2458_ _0481_ _0482_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__xnor2_1
X_2527_ _0521_ _0522_ net47 VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__mux2_1
Xhold38 top8227.demux.state_machine.currentAddress\[9\] VGND VGND VPWR VPWR net186
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold16 top8227.internalDataflow.stackBusModule.busInputs\[39\] VGND VGND VPWR VPWR
+ net164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 net15 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1409_ _0699_ _0708_ _0709_ _0710_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__o31a_2
X_2389_ top8227.internalDataflow.addressHighBusModule.busInputs\[17\] _0419_ net20
+ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__mux2_1
Xhold49 top8227.demux.state_machine.currentAddress\[10\] VGND VGND VPWR VPWR net197
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1760_ _1011_ _1028_ _1030_ _1032_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__or4_1
X_1691_ _0952_ _0953_ _0955_ _0967_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__or4_1
XFILLER_0_57_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2312_ _1195_ _1210_ _0340_ _0343_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__or4b_1
XFILLER_0_12_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2174_ _0228_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__inv_2
X_2243_ net57 _1108_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__nand2_2
XFILLER_0_28_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1958_ _1095_ _1230_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__or2_1
X_1889_ _0707_ _0817_ _1161_ net68 VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_31_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput17 net17 VGND VGND VPWR VPWR dataBusOut[7] sky130_fd_sc_hd__buf_2
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2792_ clknet_4_7_0_clk _0098_ net137 VGND VGND VPWR VPWR gpio[7] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_40_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1812_ net123 _1084_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1674_ net85 net76 net34 _0850_ _0938_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__a32o_1
X_1743_ net120 _0694_ _1015_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2226_ _0146_ _0278_ _0279_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__or3b_1
XFILLER_0_48_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2157_ top8227.internalDataflow.stackBusModule.busInputs\[32\] _1182_ _1187_ top8227.internalDataflow.accRegToDB\[0\]
+ _1183_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__a221oi_2
X_2088_ _0134_ _0141_ _0142_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1390_ net92 net95 VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_58_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2011_ _1276_ _1272_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_33_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2775_ clknet_4_7_0_clk _0081_ net137 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[22\]
+ sky130_fd_sc_hd__dfrtp_2
X_1588_ net197 net42 _0837_ _0869_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1657_ _0828_ _0840_ _0843_ _0915_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__and4_1
X_1726_ top8227.demux.state_machine.currentInstruction\[5\] _0702_ net40 _0842_ _0992_
+ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__a311o_1
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2209_ _0120_ _0263_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1511_ top8227.demux.state_machine.currentAddress\[4\] top8227.demux.state_machine.currentAddress\[10\]
+ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__or2_4
XFILLER_0_50_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2491_ _0667_ net63 _1201_ net127 VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2560_ _0780_ _0781_ _0791_ net121 VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__o31a_1
X_1442_ net93 net97 net100 net103 VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__and4b_1
XFILLER_0_10_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1373_ net80 _0674_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2758_ clknet_4_4_0_clk _0064_ net134 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2689_ clknet_4_14_0_clk _0007_ net144 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1709_ net94 _0660_ net85 net34 VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_69_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout41 net43 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_2
Xfanout30 _1136_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout63 _0739_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout52 _0714_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_2
Xfanout74 _0743_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_2
Xfanout96 top8227.demux.state_machine.currentInstruction\[2\] VGND VGND VPWR VPWR
+ net96 sky130_fd_sc_hd__buf_1
Xfanout85 _0668_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_2
XFILLER_0_51_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload11 clknet_4_12_0_clk VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__inv_6
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1991_ top8227.demux.state_machine.timeState\[5\] _0678_ net66 VGND VGND VPWR VPWR
+ _1264_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_15_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2612_ _0270_ _0584_ _0585_ _0583_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__a211o_1
X_2543_ top8227.internalDataflow.addressLowBusModule.busInputs\[21\] net20 _0533_
+ _0534_ _0536_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__o221a_1
XFILLER_0_55_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2474_ net193 _1303_ _0491_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__mux2_1
X_1425_ top8227.PSRCurrentValue\[0\] _0662_ _0669_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__or3_1
X_1356_ net99 net93 net96 net102 VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_65_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload5 clknet_4_6_0_clk VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2190_ _0771_ _0793_ net121 VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_71_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_23_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1974_ _1043_ _1064_ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2388_ _0412_ _0418_ net46 VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__mux2_1
X_2457_ top8227.internalDataflow.addressHighBusModule.busInputs\[23\] net25 VGND VGND
+ VPWR VPWR _0482_ sky130_fd_sc_hd__xnor2_1
X_2526_ _0164_ _0519_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold17 top8227.internalDataflow.stackBusModule.busInputs\[45\] VGND VGND VPWR VPWR
+ net165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 top8227.internalDataflow.stackBusModule.busInputs\[32\] VGND VGND VPWR VPWR
+ net187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 net17 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1408_ _0696_ _0703_ _0706_ _0701_ net121 VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__a311o_1
X_1339_ net128 VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1690_ _0791_ net35 net21 _0878_ _0968_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__a221o_1
X_2311_ _1220_ _0341_ _0342_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__and3_1
X_2242_ top8227.demux.setInterruptFlag net69 _1219_ top8227.demux.state_machine.currentInstruction\[5\]
+ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__a31o_1
X_2173_ _0226_ _0227_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1957_ net119 _0664_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_31_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2509_ _0355_ _0507_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__xnor2_1
X_1888_ top8227.demux.state_machine.currentAddress\[11\] top8227.demux.state_machine.currentAddress\[12\]
+ top8227.demux.state_machine.currentAddress\[4\] net126 VGND VGND VPWR VPWR _1161_
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_43_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput18 net18 VGND VGND VPWR VPWR dataBusSelect sky130_fd_sc_hd__buf_2
XFILLER_0_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2791_ clknet_4_7_0_clk _0097_ net136 VGND VGND VPWR VPWR gpio[6] sky130_fd_sc_hd__dfrtp_4
X_1811_ net86 net77 net90 VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__o21a_1
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1673_ net85 _0717_ net34 _0850_ _0922_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__a32o_1
X_1742_ _0682_ _0687_ net119 net88 VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2225_ _0278_ _0279_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2156_ top8227.internalDataflow.addressLowBusModule.busInputs\[24\] _1189_ VGND VGND
+ VPWR VPWR _0211_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_36_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2087_ _1245_ _0137_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2010_ top8227.internalDataflow.addressLowBusModule.busInputs\[39\] _1277_ _1282_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] VGND VGND VPWR VPWR
+ _1283_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_58_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2774_ clknet_4_7_0_clk _0080_ net136 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1725_ _0954_ _0961_ _0964_ _0966_ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__or4_1
X_1587_ net5 _0839_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__and2_1
X_1656_ _0723_ net34 _0850_ _0883_ _0935_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2139_ top8227.internalDataflow.accRegToDB\[1\] _1187_ _1188_ top8227.internalDataflow.addressLowBusModule.busInputs\[33\]
+ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2208_ _0145_ _0261_ _0143_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1510_ net126 net114 net112 net105 VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__nor4b_2
X_2490_ _1195_ _0342_ _0346_ _0496_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__and4b_1
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1441_ _0673_ _0706_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__nor2_2
XFILLER_0_65_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1372_ net99 net103 net93 net96 VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__and4b_4
XFILLER_0_18_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2688_ clknet_4_15_0_clk _0006_ net143 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2757_ clknet_4_4_0_clk _0063_ net129 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1708_ _0751_ net37 net21 _0908_ _0984_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__a221o_1
X_1639_ _0835_ _0913_ _0918_ _0895_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout20 _0408_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_4
Xfanout42 net43 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_52_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout31 _1136_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_4
Xfanout53 net55 VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_2
Xfanout86 net87 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_2
Xfanout64 _0738_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_4
Xfanout97 top8227.demux.state_machine.currentInstruction\[2\] VGND VGND VPWR VPWR
+ net97 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_17_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout75 _0720_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1990_ net114 net65 net72 VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2542_ _0384_ _0535_ net19 VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__o21bai_1
Xclkload12 clknet_4_13_0_clk VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_42_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2611_ top8227.internalDataflow.addressLowBusModule.busInputs\[25\] _0576_ VGND VGND
+ VPWR VPWR _0585_ sky130_fd_sc_hd__and2_1
X_2473_ net194 _1327_ _0491_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__mux2_1
X_1355_ net100 top8227.demux.state_machine.currentInstruction\[3\] net97 net103 VGND
+ VGND VPWR VPWR _0657_ sky130_fd_sc_hd__and4bb_2
X_1424_ top8227.PSRCurrentValue\[7\] net83 _0687_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload6 clknet_4_7_0_clk VGND VGND VPWR VPWR clkload6/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2809_ clknet_4_4_0_clk _0113_ net129 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1973_ _1245_ VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2525_ _0382_ _0520_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2387_ _0415_ _0417_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__xnor2_1
X_2456_ _0460_ _0471_ _0472_ net25 top8227.internalDataflow.addressHighBusModule.busInputs\[22\]
+ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__a32o_1
X_1338_ net115 VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold18 top8227.internalDataflow.stackBusModule.busInputs\[33\] VGND VGND VPWR VPWR
+ net166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 net10 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1407_ _0686_ _0691_ _0694_ _0697_ _0678_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__o41a_1
XFILLER_0_34_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2172_ _1091_ _0223_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__or2_1
X_2310_ _0771_ net73 _0761_ _0762_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__a211oi_1
XPHY_EDGE_ROW_29_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2241_ net117 net57 _0757_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_38_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1956_ net106 top8227.demux.state_machine.timeState\[1\] net66 net59 VGND VGND VPWR
+ VPWR _1229_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_31_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1887_ net53 _1158_ _1148_ VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2508_ top8227.internalDataflow.addressLowBusModule.busInputs\[16\] _0236_ net46
+ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2439_ _0452_ _0455_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2790_ clknet_4_7_0_clk _0096_ net136 VGND VGND VPWR VPWR gpio[5] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_45_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1741_ _0661_ _0695_ _0705_ net79 net118 VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__o311a_2
X_1810_ _0684_ _0694_ net108 VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1672_ _0925_ _0941_ _0951_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__or3_1
X_2224_ _0258_ _0260_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__xor2_1
X_2155_ _0200_ _0209_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2086_ _1245_ _0140_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1939_ _1195_ _1211_ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2773_ clknet_4_7_0_clk _0079_ net136 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[20\]
+ sky130_fd_sc_hd__dfrtp_2
X_1724_ _0880_ _0921_ _0997_ _0999_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1586_ net190 net41 _0857_ _0858_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__a22o_1
X_1655_ _0682_ _0907_ _0922_ _0863_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2069_ _0121_ _0122_ _0123_ _1185_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__o31a_2
X_2138_ top8227.internalDataflow.stackBusModule.busInputs\[33\] _1182_ _1183_ VGND
+ VGND VPWR VPWR _0193_ sky130_fd_sc_hd__a21o_1
X_2207_ _0145_ _0261_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1440_ _0738_ _0740_ top8227.demux.state_machine.timeState\[5\] VGND VGND VPWR VPWR
+ _0741_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1371_ top8227.demux.state_machine.currentInstruction\[5\] top8227.demux.state_machine.currentInstruction\[4\]
+ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__nand2b_4
XTAP_TAPCELL_ROW_18_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2687_ clknet_4_14_0_clk _0005_ net144 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1638_ net8 _0876_ _0896_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__a21oi_1
X_2756_ clknet_4_4_0_clk _0062_ net129 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[44\]
+ sky130_fd_sc_hd__dfrtp_1
X_1707_ net44 _0871_ _0887_ net37 _0779_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__a32o_1
XFILLER_0_26_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1569_ _0803_ _0856_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout21 _0837_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_1_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout54 net55 VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_2
Xfanout43 _0821_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout65 _0675_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout32 _1048_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
Xfanout87 _0666_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_2
Xfanout98 net101 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_2
Xfanout76 _0718_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2541_ _0368_ _0369_ _0383_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__nor3_1
Xclkload13 clknet_4_14_0_clk VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_50_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2472_ net188 _0133_ _0491_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2610_ _0277_ _0577_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__xnor2_1
X_1423_ _0719_ _0721_ _0722_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__or3_4
X_1354_ net92 net95 VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_66_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2808_ clknet_4_4_0_clk _0112_ net129 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[37\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload7 clknet_4_8_0_clk VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__inv_6
X_2739_ clknet_4_13_0_clk _0045_ net138 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_6_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1972_ _1025_ _1243_ _1244_ net48 VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__a31o_2
XFILLER_0_7_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2455_ top8227.internalDataflow.addressHighBusModule.busInputs\[22\] _0408_ _0474_
+ _0356_ _0480_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__o221a_1
X_2524_ _0374_ _0375_ _0381_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2386_ _0393_ _0399_ _0416_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold19 top8227.internalDataflow.stackBusModule.busInputs\[34\] VGND VGND VPWR VPWR
+ net167 sky130_fd_sc_hd__dlygate4sd3_1
X_1337_ net95 VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__inv_2
X_1406_ net101 _0692_ net78 _0704_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__a31o_1
XFILLER_0_52_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2171_ _0211_ _0212_ _0213_ _1184_ _1092_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__a311o_1
X_2240_ _0292_ _0294_ _0275_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__o21a_2
X_1955_ _1218_ _1226_ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__and2_4
X_1886_ net53 _1158_ _1148_ VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_31_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2507_ _0487_ gpio[15] _0506_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__mux2_1
X_2438_ _1318_ _0395_ _0464_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__a21bo_2
X_2369_ _0140_ _0163_ _0400_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1671_ _0947_ _0948_ _0949_ _0950_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__or4_1
X_1740_ _0697_ _0793_ net118 VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2085_ _1280_ _0139_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_36_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2154_ _0203_ _0208_ _1246_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__mux2_2
X_2223_ _0276_ _0277_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1869_ net70 _1076_ _1139_ _1140_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__or4_4
X_1938_ _0764_ _1198_ _1208_ _1210_ VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_57_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_66_Left_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2772_ clknet_4_6_0_clk _0078_ net136 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[19\]
+ sky130_fd_sc_hd__dfrtp_2
X_1723_ _0881_ _0909_ _0939_ _0998_ _0891_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__a2111o_1
X_1654_ _0928_ _0932_ _0933_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__or3_1
X_1585_ top8227.demux.state_machine.currentAddress\[12\] net42 _0837_ _0844_ VGND
+ VGND VPWR VPWR _0003_ sky130_fd_sc_hd__a22o_1
X_2206_ _0258_ _0260_ _0166_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2137_ net30 _0191_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__nand2_1
X_2068_ top8227.internalDataflow.stackBusModule.busInputs\[44\] _1186_ _1189_ top8227.internalDataflow.addressLowBusModule.busInputs\[28\]
+ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1370_ top8227.demux.state_machine.currentInstruction\[5\] top8227.demux.state_machine.currentInstruction\[4\]
+ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__and2b_1
XFILLER_0_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2686_ clknet_4_14_0_clk _0004_ net144 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1637_ _0803_ _0887_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2755_ clknet_4_4_0_clk _0061_ net134 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_1706_ _0934_ _0947_ _0953_ _0983_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__or4_1
X_1568_ net4 net50 _0832_ net148 VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__or4b_1
X_1499_ _0708_ _0784_ _0792_ _0797_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__or4_1
XFILLER_0_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout22 net27 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_52_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout55 net56 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
Xfanout44 _0804_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout33 _1048_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_32_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout66 _0670_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_4
Xfanout77 _0717_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_4
Xfanout88 net89 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_2
Xfanout99 net101 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_1
XFILLER_0_17_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2540_ _1334_ _0526_ _0532_ net47 VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__o31ai_1
Xclkload14 clknet_4_15_0_clk VGND VGND VPWR VPWR clkload14/Y sky130_fd_sc_hd__inv_6
XFILLER_0_50_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2471_ net198 _0157_ _0491_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__mux2_1
X_1422_ _0669_ _0683_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__nor2_1
X_1353_ top8227.demux.state_machine.currentInstruction\[4\] top8227.demux.state_machine.currentInstruction\[5\]
+ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__nand2b_4
XTAP_TAPCELL_ROW_66_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2738_ clknet_4_7_0_clk _0044_ net138 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_61_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2807_ clknet_4_4_0_clk _0111_ net129 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload8 clknet_4_9_0_clk VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__inv_8
X_2669_ _0778_ _0789_ net121 VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1971_ net111 net64 net63 _0678_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__a22oi_1
X_2385_ _1286_ _0358_ _0399_ _0402_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__and4_1
X_2454_ _0476_ _0478_ _0479_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__a21o_1
X_2523_ _0390_ _0400_ _0358_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1405_ _0701_ _0706_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__nor2_1
Xinput1 dataBusIn[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_2
X_1336_ net98 VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2170_ net30 _0215_ _0219_ _0224_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__o31a_2
X_1954_ _1218_ _1226_ VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__nor2_4
XFILLER_0_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1885_ _0812_ _1089_ _1140_ _1157_ VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_31_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2506_ _0478_ gpio[14] _0506_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__mux2_1
X_2437_ _1319_ _0394_ _0397_ _1324_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__o22a_1
X_2368_ _0185_ _0207_ _0236_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2299_ _1255_ net176 _0331_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1670_ net6 _0826_ net21 _0793_ net34 VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__a32o_1
X_2222_ _0253_ _0254_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__xnor2_2
X_2153_ _0207_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__inv_2
X_2084_ net148 _1281_ _1284_ top8227.internalDataflow.addressLowBusModule.busInputs\[28\]
+ _0138_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_36_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1937_ net90 _0671_ net76 _1209_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__a31o_1
X_1868_ net70 _0812_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__nand2_1
X_1799_ net28 VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2771_ clknet_4_7_0_clk _0077_ net137 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_41_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1584_ net146 net29 net61 _0866_ _0868_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__a41o_1
X_1722_ top8227.demux.state_machine.currentInstruction\[4\] _0702_ net40 _0955_ _0992_
+ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__a311o_1
X_1653_ _0927_ _0930_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2205_ _0166_ _0259_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__and2b_1
X_2136_ _1127_ _0190_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__nor2_1
X_2067_ top8227.internalDataflow.accRegToDB\[4\] _1187_ _1188_ top8227.internalDataflow.addressLowBusModule.busInputs\[36\]
+ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_14_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2754_ clknet_4_5_0_clk _0060_ net134 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1705_ _0900_ _0965_ _0981_ _0982_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__or4_1
X_2685_ clknet_4_14_0_clk _0000_ net144 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_1567_ net44 _0854_ _0855_ net41 net202 VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__a32o_1
X_1636_ net80 _0695_ net40 _0866_ _0915_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__a32o_1
XFILLER_0_41_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2119_ _0171_ _0172_ _0173_ _1185_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__o31ai_4
X_1498_ _0775_ _0795_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout23 net27 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_2
Xfanout67 net68 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_52_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout45 _0394_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_2
Xfanout56 _0713_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
Xfanout78 _0700_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_4
Xfanout89 net91 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
Xfanout34 net35 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_2
XFILLER_0_51_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2470_ net195 _0177_ _0491_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1421_ net102 _0642_ net83 net92 _0641_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_66_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1352_ top8227.demux.state_machine.currentInstruction\[4\] top8227.demux.state_machine.currentInstruction\[5\]
+ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__and2b_1
XFILLER_0_58_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2737_ clknet_4_7_0_clk _0043_ net138 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2806_ clknet_4_4_0_clk _0110_ net129 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_2668_ _0270_ _0291_ _0635_ _0634_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__a31o_1
Xclkload9 clknet_4_10_0_clk VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__inv_8
X_1619_ _0744_ net40 _0898_ net44 _0894_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2599_ _1060_ _1247_ _0573_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__or3_1
XFILLER_0_66_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1970_ net66 _0809_ _1031_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2522_ net19 _0517_ _0518_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__o21a_1
X_2453_ _0476_ _0478_ net46 VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__o21ai_1
X_2384_ _0197_ _0394_ _0413_ _0414_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__o211ai_4
X_1404_ net102 net92 net95 net98 VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__or4b_2
Xinput2 dataBusIn[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_4
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_2_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1953_ net55 _1222_ _1225_ VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1884_ _1150_ _1153_ _1156_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2505_ _0465_ gpio[13] _0506_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2436_ _0459_ _0462_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__xnor2_1
X_2367_ _0214_ _0396_ _0398_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2298_ _1308_ net161 _0331_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2152_ top8227.internalDataflow.addressLowBusModule.busInputs\[25\] _1284_ _0204_
+ _1280_ _0206_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__a221o_2
X_2221_ _0255_ _0257_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2083_ top8227.internalDataflow.addressLowBusModule.busInputs\[36\] _1277_ _1282_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[20\] VGND VGND VPWR VPWR
+ _0138_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1867_ net115 _0724_ _0735_ net70 VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__a31o_1
X_1936_ _0664_ _0678_ _0747_ _1064_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1798_ _1058_ _1067_ _1070_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__o21a_1
X_2419_ _0444_ _0446_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2770_ clknet_4_7_0_clk _0076_ net138 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1721_ _0949_ _0993_ _0994_ _0996_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1583_ top8227.demux.state_machine.currentAddress\[2\] net41 net21 _0860_ _0867_
+ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1652_ net147 _0826_ _0850_ _0931_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__a31o_1
X_2135_ top8227.internalDataflow.addressLowBusModule.busInputs\[17\] _1129_ _0188_
+ _0189_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__a211oi_1
X_2204_ net28 _0157_ _0165_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_44_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2066_ top8227.internalDataflow.stackBusModule.busInputs\[36\] _1182_ _1183_ VGND
+ VGND VPWR VPWR _0121_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1919_ top8227.internalDataflow.addressLowBusModule.busInputs\[39\] _1188_ _1191_
+ _1183_ VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2753_ clknet_4_4_0_clk _0059_ net135 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2684_ top8227.PSRCurrentValue\[7\] _1255_ _0640_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__mux2_1
X_1704_ _0969_ _0972_ _0977_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__or3_1
X_1566_ net50 _0851_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__nor2_1
X_1635_ _0803_ _0914_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1497_ _0741_ _0749_ _0754_ _0788_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__or4_1
XFILLER_0_68_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2049_ top8227.internalDataflow.addressHighBusModule.busInputs\[21\] _1120_ _1130_
+ top8227.internalDataflow.accRegToDB\[5\] VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__a22o_1
X_2118_ top8227.internalDataflow.stackBusModule.busInputs\[42\] _1186_ _1188_ top8227.internalDataflow.addressLowBusModule.busInputs\[34\]
+ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout24 net27 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
Xfanout46 net47 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
Xfanout68 net69 VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_52_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout57 net58 VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_4
Xfanout79 net82 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_2
Xfanout35 net38 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_2
XFILLER_0_32_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1351_ _0653_ VGND VGND VPWR VPWR top8227.pulse_slower.nextEnableState\[0\] sky130_fd_sc_hd__inv_2
X_1420_ net97 _0660_ net85 VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_66_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2805_ clknet_4_4_0_clk _0109_ net129 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2736_ clknet_4_7_0_clk _0042_ net138 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_1618_ net54 _0895_ _0896_ _0897_ _0835_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__a32o_1
XFILLER_0_41_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2667_ _0586_ _0624_ _0289_ _0291_ _0293_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_14_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1549_ _0838_ _0839_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2598_ _1010_ _1038_ _1063_ _0572_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__or4_1
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2521_ net47 _0515_ net20 top8227.internalDataflow.addressLowBusModule.busInputs\[18\]
+ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2452_ _1300_ _0395_ _0477_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__a21bo_1
X_2383_ _0192_ _0394_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__nand2b_1
X_1403_ net104 net94 top8227.demux.state_machine.currentInstruction\[2\] net101 VGND
+ VGND VPWR VPWR _0705_ sky130_fd_sc_hd__nor4b_2
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 dataBusIn[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2719_ clknet_4_2_0_clk _0029_ net132 VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1952_ net67 _0815_ _0818_ _1223_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__or4_1
XFILLER_0_43_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1883_ _0749_ _1029_ _1154_ _1155_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__or4_1
X_2504_ _0456_ gpio[12] _0506_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__mux2_1
X_2435_ _0460_ _0461_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2366_ _0218_ net45 _0397_ _0223_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_39_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2297_ _1329_ net175 _0331_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2151_ top8227.internalDataflow.addressLowBusModule.busInputs\[33\] _1277_ _1281_
+ net2 _0205_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__a221o_1
X_2082_ _1253_ _1256_ _0135_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__mux2_1
X_2220_ net33 _0267_ _0274_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_44_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1797_ net67 _1068_ _1069_ net53 _1057_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__o311a_1
X_1866_ net50 _1138_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__or2_1
X_1935_ _1200_ _1202_ _1203_ _1207_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2418_ top8227.internalDataflow.addressHighBusModule.busInputs\[20\] net26 VGND VGND
+ VPWR VPWR _0446_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2349_ _0378_ _0380_ _0377_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_35_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_44_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1720_ _0902_ _0929_ _0935_ _0995_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__or4_1
X_1651_ net85 _0674_ net35 VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__and3_1
X_1582_ net54 gpio[21] _0828_ _0844_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__and4_1
XFILLER_0_21_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_53_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2134_ top8227.PSRCurrentValue\[1\] _1132_ _1133_ net2 VGND VGND VPWR VPWR _0189_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2065_ _0118_ _0119_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__nand2_1
X_2203_ _0255_ _0257_ _0187_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1849_ net50 _1119_ _1121_ _1106_ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__o211a_2
X_1918_ top8227.internalDataflow.stackBusModule.busInputs\[47\] _1186_ _1187_ top8227.internalDataflow.accRegToDB\[7\]
+ _1190_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1634_ net51 _0883_ _0903_ _0913_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2752_ clknet_4_9_0_clk _0058_ net133 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1703_ _0721_ net37 _0973_ _0974_ _0980_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_26_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2683_ _0745_ _1062_ _1108_ _0303_ net57 VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_69_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1565_ _0829_ _0853_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__or2_1
X_1496_ _0662_ _0696_ _0673_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__a21oi_1
X_2048_ net147 _1133_ _1122_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__a21oi_1
X_2117_ top8227.internalDataflow.accRegToDB\[2\] _1187_ _1189_ top8227.internalDataflow.addressLowBusModule.busInputs\[26\]
+ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout25 net27 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_4
Xfanout47 _0335_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_2
Xfanout69 _0652_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_52_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout36 net38 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_2
Xfanout58 net60 VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1350_ top8227.pulse_slower.currentEnableState\[1\] top8227.pulse_slower.currentEnableState\[0\]
+ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__or2_4
XFILLER_0_58_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2804_ clknet_4_4_0_clk _0108_ net130 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1617_ net51 _0892_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__nor2_2
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2735_ clknet_4_3_0_clk _0041_ net131 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfrtp_1
X_2666_ top8227.internalDataflow.addressLowBusModule.busInputs\[31\] _0576_ _0633_
+ _0271_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2597_ _0684_ _0690_ _0694_ _0750_ net117 VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__o41a_1
XFILLER_0_66_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1548_ net3 net61 net4 VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__and3b_1
X_1479_ _0700_ net74 VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2520_ _0381_ _0516_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__nor2_1
X_2451_ _1301_ _1296_ net45 VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1402_ _0701_ _0703_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__nor2_1
X_2382_ _0196_ _0395_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__nand2_1
Xinput4 dataBusIn[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_62_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2718_ clknet_4_11_0_clk _0028_ net142 VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.resetDetected
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2649_ _0265_ _0617_ net32 VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1951_ _0815_ _1223_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1882_ net109 _0694_ _0759_ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2503_ _0441_ gpio[11] _0506_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__mux2_1
X_2434_ top8227.internalDataflow.addressHighBusModule.busInputs\[21\] net25 VGND VGND
+ VPWR VPWR _0461_ sky130_fd_sc_hd__nand2_1
X_2365_ net30 net45 VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2296_ _0136_ net162 _0331_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2150_ top8227.internalDataflow.addressLowBusModule.busInputs\[17\] _1271_ _1278_
+ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__and3_1
X_2081_ _0135_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1934_ net65 _1206_ _1205_ _1204_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1796_ top8227.demux.state_machine.currentAddress\[12\] _0816_ net124 VGND VGND VPWR
+ VPWR _1069_ sky130_fd_sc_hd__o21a_1
X_1865_ _1031_ _1058_ _1123_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__nor3_1
XFILLER_0_24_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2417_ top8227.internalDataflow.addressHighBusModule.busInputs\[20\] net26 VGND VGND
+ VPWR VPWR _0445_ sky130_fd_sc_hd__nand2_1
X_2348_ top8227.internalDataflow.addressLowBusModule.busInputs\[16\] _0379_ VGND VGND
+ VPWR VPWR _0380_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2279_ top8227.demux.setInterruptFlag top8227.PSRCurrentValue\[2\] VGND VGND VPWR
+ VPWR _0324_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1581_ _0831_ _0843_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_41_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1650_ net91 _0674_ net38 _0881_ _0893_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__a32o_1
X_2202_ _0187_ _0256_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2133_ top8227.internalDataflow.addressHighBusModule.busInputs\[17\] _1120_ _1130_
+ top8227.internalDataflow.accRegToDB\[1\] _1122_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2064_ _1331_ _1335_ _1328_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1917_ top8227.internalDataflow.stackBusModule.busInputs\[39\] _1182_ _1189_ top8227.internalDataflow.addressLowBusModule.busInputs\[31\]
+ VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1779_ _0677_ _1051_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__or2_1
X_1848_ _1096_ _1115_ _1116_ net59 VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2751_ clknet_4_9_0_clk _0057_ net135 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2682_ net199 net41 _0639_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__o21ai_1
X_1564_ net7 _0852_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__nor2_2
X_1633_ _0826_ _0876_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1702_ _0796_ net37 _0884_ _0979_ _0978_ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1495_ _0662_ _0673_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__nor2_1
Xfanout26 net27 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_52_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2047_ top8227.internalDataflow.addressLowBusModule.busInputs\[21\] _1129_ VGND VGND
+ VPWR VPWR _1320_ sky130_fd_sc_hd__nand2_1
Xfanout37 net38 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
X_2116_ top8227.internalDataflow.stackBusModule.busInputs\[34\] _1182_ _1183_ VGND
+ VGND VPWR VPWR _0171_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_1_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout59 net60 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_4
Xfanout48 _0716_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_4
XFILLER_0_17_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2803_ clknet_4_1_0_clk _0107_ net133 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2734_ clknet_4_0_0_clk _0040_ net130 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1547_ net148 net4 _0832_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__a21oi_2
X_1616_ net146 net7 net62 VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2665_ net33 _0628_ _0629_ _0632_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__a31o_1
X_2596_ net33 _0568_ _0570_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_65_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1478_ _0688_ _0701_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__nor2_2
XFILLER_0_64_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2381_ _0410_ _0411_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__xnor2_1
X_2450_ _0465_ _0466_ _0475_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_23_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1401_ net98 net102 net92 net95 VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__or4_2
Xinput5 dataBusIn[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
XFILLER_0_36_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2717_ clknet_4_12_0_clk _0027_ net138 VGND VGND VPWR VPWR top8227.freeCarry sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2579_ _0207_ gpio[1] _0560_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__mux2_1
X_2648_ _1314_ _0118_ _0264_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1950_ net113 net106 _0807_ _0814_ top8227.demux.state_machine.currentAddress\[6\]
+ VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__o221a_1
X_2502_ _0430_ gpio[10] _0506_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1881_ top8227.demux.state_machine.timeState\[1\] net65 _0786_ net109 VGND VGND VPWR
+ VPWR _1154_ sky130_fd_sc_hd__a22o_1
X_2433_ top8227.internalDataflow.addressHighBusModule.busInputs\[21\] net25 VGND VGND
+ VPWR VPWR _0460_ sky130_fd_sc_hd__or2_1
X_2364_ _1077_ net45 VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__nand2_2
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2295_ _0159_ net183 _0331_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_9_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
X_2080_ _1091_ _0124_ _0131_ _1128_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_17_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1933_ net105 top8227.demux.state_machine.timeState\[5\] VGND VGND VPWR VPWR _1206_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_71_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1795_ net124 _0811_ _0814_ net128 VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__a22o_1
X_1864_ _1077_ _1128_ _1135_ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2416_ top8227.internalDataflow.addressHighBusModule.busInputs\[20\] net26 VGND VGND
+ VPWR VPWR _0444_ sky130_fd_sc_hd__and2_1
X_2347_ top8227.internalDataflow.addressLowBusModule.busInputs\[17\] net22 VGND VGND
+ VPWR VPWR _0379_ sky130_fd_sc_hd__xor2_1
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2278_ top8227.instructionLoader.interruptInjector.resetDetected net52 VGND VGND
+ VPWR VPWR _0028_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1580_ _0648_ _0804_ _0865_ _0864_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2132_ _0178_ _0182_ _0186_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__nor3_1
X_2201_ _0182_ _0186_ _0178_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2063_ _1328_ _1331_ _1335_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__or3_2
XFILLER_0_71_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1847_ _1096_ _1117_ net59 VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__and3b_2
XFILLER_0_44_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1916_ _1160_ _1170_ _1180_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__and3_2
XFILLER_0_29_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1778_ net125 top8227.demux.state_machine.currentAddress\[12\] VGND VGND VPWR VPWR
+ _1051_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2681_ top8227.demux.isAddressing net51 _0819_ net68 VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1701_ _0835_ _0866_ _0895_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__or3_1
X_2750_ clknet_4_5_0_clk _0056_ net134 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1563_ net146 net61 VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__nand2_1
X_1632_ _0695_ _0907_ _0911_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1494_ _0693_ _0706_ _0669_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__a21oi_1
X_2115_ _1077_ _1128_ _0169_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__or3_1
Xfanout27 _0357_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
X_2046_ top8227.internalDataflow.addressHighBusModule.busInputs\[21\] _1227_ _1228_
+ net147 _1234_ VGND VGND VPWR VPWR _1319_ sky130_fd_sc_hd__a221oi_2
Xfanout38 net43 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout49 net52 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_17_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2802_ clknet_4_8_0_clk net158 net141 VGND VGND VPWR VPWR top8227.pulse_slower.currentEnableState\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2733_ clknet_4_2_0_clk _0039_ net131 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2664_ _1289_ _0567_ _0630_ _0631_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_51 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1615_ _0831_ _0851_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__nor2_1
X_1546_ _0822_ _0836_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__and2_1
X_2595_ _0200_ _0273_ _0566_ _0241_ _0569_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__o221a_1
X_1477_ _0658_ _0701_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Left_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2029_ _1143_ _1300_ _1301_ _1142_ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_37_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_68_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2380_ top8227.internalDataflow.addressHighBusModule.busInputs\[17\] net24 VGND VGND
+ VPWR VPWR _0411_ sky130_fd_sc_hd__xor2_1
X_1400_ net100 net103 net94 net97 VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__nor4_2
Xinput6 dataBusIn[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_62_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2647_ _0616_ top8227.internalDataflow.addressLowBusModule.busInputs\[29\] _0576_
+ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__mux2_1
X_2716_ clknet_4_0_0_clk top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[6\]
+ net131 VGND VGND VPWR VPWR top8227.PSRCurrentValue\[6\] sky130_fd_sc_hd__dfrtp_2
X_2578_ _0236_ gpio[0] _0560_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__mux2_1
X_1529_ top8227.demux.state_machine.timeState\[5\] net49 _0820_ top8227.demux.state_machine.timeState\[1\]
+ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1880_ _1112_ _1151_ _1152_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__or3_1
X_2501_ _0415_ gpio[9] _0506_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2432_ _0446_ _0450_ _0445_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__o21ai_1
X_2363_ _1077_ net45 VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2294_ _0180_ net180 _0331_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1863_ _1077_ _1091_ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__nor2_1
X_1932_ net91 _0671_ _0682_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2415_ top8227.internalDataflow.addressHighBusModule.busInputs\[19\] _0408_ _0435_
+ net19 _0443_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__o221a_1
XFILLER_0_58_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1794_ _0665_ _1061_ _1064_ _1066_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__or4_1
X_2346_ top8227.internalDataflow.addressLowBusModule.busInputs\[17\] net22 VGND VGND
+ VPWR VPWR _0378_ sky130_fd_sc_hd__and2_1
X_2277_ net152 _0295_ _0323_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2131_ _1245_ _0185_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__nor2_1
X_2062_ _1245_ _1334_ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__nor2_1
X_2200_ _0253_ _0254_ _0210_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1777_ net128 top8227.demux.state_machine.currentAddress\[6\] VGND VGND VPWR VPWR
+ _1050_ sky130_fd_sc_hd__or2_1
X_1846_ _1115_ _1116_ _1105_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1915_ _1160_ _1171_ _1180_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__and3_2
XFILLER_0_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_31_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2329_ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] net23 VGND VGND
+ VPWR VPWR _0361_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_40_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_8_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2680_ _0295_ _0638_ net192 _1242_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_53_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1631_ net44 _0838_ _0848_ _0887_ _0910_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__a41o_1
XFILLER_0_41_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1700_ _0782_ net36 _0863_ _0878_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1562_ net148 net4 _0832_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__or3_1
X_1493_ _0669_ _0706_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2114_ top8227.internalDataflow.addressLowBusModule.busInputs\[18\] _1129_ _0168_
+ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__a21oi_1
X_2045_ _1315_ _1316_ _1317_ _1185_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__o31a_1
XFILLER_0_71_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout39 net43 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
Xfanout28 _1071_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_17_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1829_ net70 _1101_ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_68_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2801_ clknet_4_8_0_clk top8227.pulse_slower.nextEnableState\[0\] net141 VGND VGND
+ VPWR VPWR top8227.pulse_slower.currentEnableState\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1614_ _0786_ net39 _0889_ _0893_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2732_ clknet_4_2_0_clk _0038_ net131 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2663_ _0252_ _0272_ _0563_ _1291_ _0565_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__a221o_1
X_2594_ _0655_ _0696_ _1240_ _0240_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__or4b_1
XFILLER_0_66_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1545_ net2 net1 net61 VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__and3b_1
X_1476_ net82 _0702_ _0776_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2028_ top8227.internalDataflow.addressHighBusModule.busInputs\[22\] _1227_ _1228_
+ net7 _1234_ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 dataBusIn[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_19_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2577_ _0504_ _0559_ _0558_ net50 VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__a211o_4
X_2646_ _0270_ _0614_ _0615_ _0613_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__a31o_1
X_2715_ clknet_4_3_0_clk top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[3\]
+ net131 VGND VGND VPWR VPWR top8227.PSRCurrentValue\[3\] sky130_fd_sc_hd__dfrtp_2
X_1459_ net125 net81 net75 VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__and3_1
X_1528_ net108 net52 _0820_ net121 VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2431_ top8227.internalDataflow.addressHighBusModule.busInputs\[20\] net20 _0451_
+ net19 _0458_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__o221a_1
X_2500_ _0399_ gpio[8] _0506_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2362_ net70 _1138_ _1140_ _1141_ net53 VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__o2111a_2
X_2293_ _0201_ net172 _0331_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2629_ _0260_ _0565_ _0600_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1862_ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] _1129_ _1134_
+ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__a21oi_1
X_1931_ net80 _0755_ net73 VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__and3_1
X_1793_ _1016_ _1030_ _1063_ _1065_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__or4_1
X_2414_ _0438_ _0440_ _0442_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2345_ _0375_ _0376_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__nor2_1
X_2276_ net70 net53 _1068_ _1241_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_35_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2061_ _1280_ _1333_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__or2_2
X_2130_ _0647_ _1280_ _1284_ top8227.internalDataflow.addressLowBusModule.busInputs\[26\]
+ _0184_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__a221o_2
XFILLER_0_56_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1914_ _1172_ _1181_ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__nor2_2
XFILLER_0_29_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1776_ _0811_ _0814_ net67 VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__a21oi_1
X_1845_ _1115_ _1116_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2328_ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] net23 VGND VGND
+ VPWR VPWR _0360_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2259_ _0309_ _0310_ _0311_ VGND VGND VPWR VPWR top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[2\]
+ sky130_fd_sc_hd__or3_1
XFILLER_0_62_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1630_ net87 _0907_ _0908_ _0863_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1561_ net151 net41 _0850_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1492_ _0669_ _0693_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__nor2_2
XFILLER_0_55_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2113_ top8227.PSRCurrentValue\[2\] _1132_ _1133_ net3 _0167_ VGND VGND VPWR VPWR
+ _0168_ sky130_fd_sc_hd__a221o_1
X_2044_ top8227.internalDataflow.stackBusModule.busInputs\[37\] _1182_ _1189_ top8227.internalDataflow.addressLowBusModule.busInputs\[29\]
+ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout29 _0822_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_2
XFILLER_0_29_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1828_ _0813_ _0817_ _0818_ _0704_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_44_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1759_ net64 _0809_ _1031_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_68_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2731_ clknet_4_0_0_clk _0037_ net130 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfrtp_1
X_2800_ clknet_4_0_0_clk _0106_ net130 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_1544_ top8227.demux.state_machine.currentAddress\[6\] net42 _0827_ _0835_ VGND VGND
+ VPWR VPWR _0009_ sky130_fd_sc_hd__a22o_1
X_1613_ net39 _0892_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2662_ _1292_ _0566_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__or2_1
X_2593_ _0239_ _0567_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_7_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_1475_ net85 _0766_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_65_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2027_ _1297_ _1298_ _1299_ _1185_ VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__o31a_1
XFILLER_0_60_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 dataBusIn[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
X_2714_ clknet_4_2_0_clk top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[2\]
+ net132 VGND VGND VPWR VPWR top8227.PSRCurrentValue\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2576_ net128 _0809_ _0811_ net73 _0350_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__a221oi_2
X_1527_ top8227.demux.state_machine.timeState\[3\] net49 _0820_ top8227.demux.state_machine.timeState\[5\]
+ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__a22o_1
X_2645_ _0288_ _0291_ _0293_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__nand3_1
X_1458_ net112 net86 net81 VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__and3_1
X_1389_ _0683_ _0688_ _0655_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2430_ _0453_ _0455_ _0457_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__o21ai_1
X_2361_ _1286_ _1306_ _0358_ _0392_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2292_ _0229_ net177 _0331_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2559_ _0751_ _0771_ _0799_ net109 VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__o31a_1
XFILLER_0_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2628_ _0259_ _0563_ _0567_ _0166_ _0599_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_38_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1930_ _0671_ _0694_ _0790_ net73 _0770_ VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1861_ top8227.PSRCurrentValue\[7\] _1132_ _1133_ net146 _1131_ VGND VGND VPWR VPWR
+ _1134_ sky130_fd_sc_hd__a221o_1
X_1792_ net68 _1035_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__nand2_1
X_2413_ _0438_ _0440_ net46 VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__o21ai_1
X_2344_ top8227.internalDataflow.addressLowBusModule.busInputs\[18\] net27 VGND VGND
+ VPWR VPWR _0376_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2275_ top8227.branchForward _1242_ _0295_ _0322_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2060_ net147 _1281_ _1284_ top8227.internalDataflow.addressLowBusModule.busInputs\[29\]
+ _1332_ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1913_ _1172_ _1180_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__nor2_2
XFILLER_0_29_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1844_ _1115_ _1116_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__and2_1
X_1775_ _1024_ _1047_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2327_ top8227.internalDataflow.addressHighBusModule.busInputs\[16\] net23 VGND VGND
+ VPWR VPWR _0359_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2258_ top8227.demux.setInterruptFlag net57 _1219_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2189_ top8227.branchForward _1034_ _1054_ _0243_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__a211o_1
XFILLER_0_35_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1560_ net44 _0830_ _0849_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__and3_4
XFILLER_0_53_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2112_ top8227.internalDataflow.addressHighBusModule.busInputs\[18\] _1120_ _1130_
+ top8227.internalDataflow.accRegToDB\[2\] _1122_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__a221o_1
X_1491_ _0790_ _0791_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__or2_1
Xfanout19 _0356_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
XFILLER_0_55_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2043_ top8227.internalDataflow.accRegToDB\[5\] _1187_ _1188_ top8227.internalDataflow.addressLowBusModule.busInputs\[37\]
+ VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__a22o_1
X_1827_ net67 _1099_ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1758_ net122 net81 _0674_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__and3_2
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1689_ _0756_ net35 _0881_ _0956_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2730_ clknet_4_0_0_clk _0036_ net131 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfrtp_1
X_2661_ _1292_ _0315_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__or2_1
X_1543_ _0831_ _0833_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__nor2_1
X_1612_ _0648_ _0876_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2592_ net48 _1167_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__nor2_2
X_1474_ net87 _0682_ net77 net75 net78 VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__o41a_1
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2026_ top8227.internalDataflow.stackBusModule.busInputs\[46\] _1186_ _1187_ top8227.internalDataflow.accRegToDB\[6\]
+ VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_28_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 nrst VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2713_ clknet_4_0_0_clk top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[1\]
+ net131 VGND VGND VPWR VPWR top8227.PSRCurrentValue\[1\] sky130_fd_sc_hd__dfrtp_1
X_2644_ _0289_ _0291_ _0293_ _0288_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1526_ net71 net55 _0819_ net29 _0823_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__a311o_1
X_2575_ _1262_ _0557_ _0336_ _0497_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__and4bb_1
X_1457_ top8227.demux.state_machine.timeState\[3\] net86 net85 VGND VGND VPWR VPWR
+ _0758_ sky130_fd_sc_hd__and3_1
X_1388_ _0655_ _0683_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__nor2_1
X_2009_ _1271_ _1278_ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_6_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
X_2360_ _1334_ _0140_ _0391_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__or3_1
X_2291_ _1090_ _1102_ _0330_ net50 VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__a211o_4
XFILLER_0_47_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2627_ net28 _0133_ _0272_ net32 VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2558_ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] _0409_ _0546_
+ _0549_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__a211o_1
X_1509_ net114 net73 VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__or2_4
X_2489_ net112 _0787_ _1199_ _1210_ _1230_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__a2111oi_1
XTAP_TAPCELL_ROW_38_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1860_ net53 _1098_ _1105_ _1118_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_44_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1791_ net119 net89 _0695_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__and3_1
X_2412_ _0440_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2343_ top8227.internalDataflow.addressLowBusModule.busInputs\[18\] net22 VGND VGND
+ VPWR VPWR _0375_ sky130_fd_sc_hd__and2_1
X_2274_ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] _0648_ _1241_
+ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1989_ top8227.demux.state_machine.timeState\[1\] net63 _1084_ _0680_ VGND VGND VPWR
+ VPWR _1262_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1843_ net70 _1093_ _1100_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1912_ net48 _1035_ _1183_ VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1774_ _1033_ _1034_ _1046_ _1025_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__or4b_1
XFILLER_0_12_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2326_ net24 VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2257_ _0673_ _0703_ _1240_ _0298_ top8227.PSRCurrentValue\[2\] VGND VGND VPWR VPWR
+ _0310_ sky130_fd_sc_hd__o311a_1
XFILLER_0_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2188_ net64 net73 _0809_ net63 _1014_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1490_ net82 _0755_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2042_ top8227.internalDataflow.stackBusModule.busInputs\[45\] _1186_ _1183_ VGND
+ VGND VPWR VPWR _1315_ sky130_fd_sc_hd__a21o_1
X_2111_ _1072_ _0165_ _0157_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__nor3b_1
Xhold1 top8227.instructionLoader.interruptInjector.irqSync.nextQ2 VGND VGND VPWR VPWR
+ net149 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1826_ net111 net66 net65 net114 VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1757_ net120 _0742_ _1029_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__a21o_1
X_1688_ _0794_ net34 net21 _0897_ _0966_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _0744_ _0806_ _1201_ net64 VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_0_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1611_ net80 net74 net39 _0890_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__a31o_1
X_2660_ _1292_ _0315_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__nand2_1
X_1542_ net29 _0833_ _0834_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2591_ _0673_ _0688_ _1240_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__or3_2
X_1473_ net87 net75 net78 VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_65_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2025_ top8227.internalDataflow.addressLowBusModule.busInputs\[38\] _1188_ _1189_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[30\] VGND VGND VPWR VPWR
+ _1298_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2789_ clknet_4_7_0_clk _0095_ net136 VGND VGND VPWR VPWR gpio[4] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_32_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1809_ net87 net77 net73 net79 VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2574_ _0670_ _0553_ _0554_ _0556_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__a211o_1
XFILLER_0_22_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2712_ clknet_4_3_0_clk top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[0\]
+ net132 VGND VGND VPWR VPWR top8227.PSRCurrentValue\[0\] sky130_fd_sc_hd__dfrtp_4
X_2643_ _0270_ _0612_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__nor2_1
X_1525_ net125 top8227.demux.state_machine.timeState\[3\] net55 VGND VGND VPWR VPWR
+ _0823_ sky130_fd_sc_hd__mux2_1
X_1387_ _0655_ _0688_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__nor2_1
X_1456_ net88 _0674_ _0755_ net83 VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__a22o_1
X_2008_ _1272_ _1276_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_25_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2290_ _1243_ _1263_ _0329_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_56_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_65_Left_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2557_ _1286_ _0547_ _0548_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2626_ _0279_ net32 VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__nand2b_1
X_1439_ net65 net63 VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__or2_1
X_1508_ net120 net116 VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__or2_1
X_2488_ top8227.instructionLoader.interruptInjector.resetDetected net56 _0495_ top8227.demux.reset
+ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1790_ net117 _0751_ _1044_ _1062_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__a211o_1
X_2411_ _0151_ net45 _0396_ _0150_ _0439_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__o221a_2
XFILLER_0_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2342_ _0372_ _0373_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__nor2_1
X_2273_ gpio[18] net69 _0711_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__nand3_1
X_1988_ net125 _0644_ _0677_ _1049_ _1260_ VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__o311a_1
XFILLER_0_47_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2609_ net32 _0582_ _0578_ _0271_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__o211a_1
Xclkbuf_4_5_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_65_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1842_ _1022_ _1107_ _1114_ _1075_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1911_ net48 _1035_ _1183_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1773_ _1013_ _1043_ _1044_ _1045_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__or4_1
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2325_ _0803_ _0824_ _0352_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__o21ai_1
X_2187_ net123 net128 _1089_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__a21bo_1
X_2256_ _0179_ _0298_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2110_ _0160_ _0164_ _1246_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__mux2_1
Xhold2 top8227.instructionLoader.interruptInjector.nmiSync.nextQ2 VGND VGND VPWR VPWR
+ net150 sky130_fd_sc_hd__dlygate4sd3_1
X_2041_ _1312_ _1313_ VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_29_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1825_ net59 _1097_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1756_ net109 net105 net65 VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2308_ _0740_ _1201_ _0339_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__a21o_1
X_1687_ net89 _0705_ net34 _0863_ _0938_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_68_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2239_ _0270_ _0293_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1610_ net54 net44 _0887_ _0889_ _0888_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_14_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2590_ net117 net57 _0751_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__and3_1
X_1541_ top8227.demux.state_machine.currentAddress\[7\] net29 _0827_ _0830_ VGND VGND
+ VPWR VPWR _0834_ sky130_fd_sc_hd__a2bb2o_1
X_1472_ net110 _0769_ _0772_ _0768_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2024_ top8227.internalDataflow.stackBusModule.busInputs\[38\] _1182_ _1183_ VGND
+ VGND VPWR VPWR _1297_ sky130_fd_sc_hd__a21o_1
XFILLER_0_64_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2788_ clknet_4_6_0_clk _0094_ net136 VGND VGND VPWR VPWR gpio[3] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1808_ _0745_ _0746_ _0753_ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__or3_1
X_1739_ _1010_ _1011_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2711_ clknet_4_10_0_clk _0025_ net142 VGND VGND VPWR VPWR top8227.demux.state_machine.currentInstruction\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_1524_ net42 VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__inv_2
X_2573_ _0676_ _1205_ _0555_ _0341_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__or4b_1
X_2642_ net32 _0264_ _0611_ _0610_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_10_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1386_ net98 net102 net95 net92 VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__or4b_4
X_1455_ net89 _0755_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__and2_1
X_2007_ _1229_ _1279_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__nor2_2
XFILLER_0_26_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2556_ _1286_ _0547_ net47 VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__o21ai_1
X_1507_ net125 net114 VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__nor2_1
X_2487_ net56 _0324_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__nand2_1
X_2625_ _0166_ _0271_ _0278_ _0596_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__or4b_1
XFILLER_0_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1438_ net90 net77 VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__and2_1
X_1369_ net114 net105 VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__or2_2
XFILLER_0_65_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2341_ top8227.internalDataflow.addressLowBusModule.busInputs\[19\] net22 VGND VGND
+ VPWR VPWR _0373_ sky130_fd_sc_hd__nor2_1
X_2410_ net30 _0156_ net45 VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__nand3_1
X_2272_ clknet_4_8_0_clk top8227.pulse_slower.nextEnableState\[0\] VGND VGND VPWR
+ VPWR gpio[24] sky130_fd_sc_hd__and2_2
XFILLER_0_59_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1987_ _0814_ _0816_ _1051_ _0679_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_15_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2539_ _0526_ _0532_ _1334_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__o21a_1
X_2608_ _0580_ _0581_ _0210_ _0567_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1910_ _1159_ _1181_ _1179_ _1172_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__o211a_4
XFILLER_0_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1841_ _1109_ _1110_ _1111_ _1113_ VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__or4_2
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1772_ net117 _1039_ _1042_ _1038_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__a211o_1
X_2324_ net46 _0355_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__or2_1
X_2255_ _0179_ _0202_ _0308_ _0306_ VGND VGND VPWR VPWR top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[1\]
+ sky130_fd_sc_hd__a31o_1
X_2186_ _0239_ _0240_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3 top8227.demux.state_machine.currentAddress\[8\] VGND VGND VPWR VPWR net151
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2040_ _1304_ _1311_ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_71_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1824_ top8227.branchForward _1034_ _1094_ _1095_ _1031_ VGND VGND VPWR VPWR _1097_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_40_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_4_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
X_1686_ _0962_ _0963_ _0964_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__or3_1
XFILLER_0_25_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1755_ net119 _1027_ _1026_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__a21o_1
X_2307_ _0758_ _1199_ _1205_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2238_ _0266_ _0284_ _1290_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_68_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2169_ net30 _0223_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1540_ _0832_ net148 net4 VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__or3b_1
XFILLER_0_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1471_ net116 _0659_ _0771_ net109 _0770_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2023_ _1077_ _1128_ _1295_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__or3_2
XFILLER_0_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1807_ _0691_ _0771_ _0775_ net108 VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__o31a_1
X_2787_ clknet_4_6_0_clk _0093_ net136 VGND VGND VPWR VPWR gpio[2] sky130_fd_sc_hd__dfrtp_4
X_1669_ _0765_ net37 _0881_ _0943_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1738_ net118 net88 net75 VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__and3_2
XFILLER_0_31_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2710_ clknet_4_10_0_clk _0024_ net144 VGND VGND VPWR VPWR top8227.demux.state_machine.currentInstruction\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1523_ top8227.instructionLoader.interruptInjector.resetDetected net54 gpio[21] VGND
+ VGND VPWR VPWR _0821_ sky130_fd_sc_hd__a21oi_1
X_2572_ net127 _1201_ _0675_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__o21a_1
X_1454_ net104 net93 net96 net99 VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__and4b_2
X_2641_ _0120_ _0263_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1385_ net98 net102 net95 net92 VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__nor4b_2
XFILLER_0_45_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2006_ _1272_ _1277_ _1278_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2624_ _0276_ _0277_ _0586_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__or3_1
X_2555_ net24 _0402_ _0541_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__o21ba_1
X_1506_ net125 net113 VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__or2_2
X_1437_ net90 net86 VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__and2_1
X_2486_ net168 _1237_ _0494_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1368_ net86 net85 VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2340_ top8227.internalDataflow.addressLowBusModule.busInputs\[19\] net22 VGND VGND
+ VPWR VPWR _0372_ sky130_fd_sc_hd__and2_1
X_2271_ _1308_ _0318_ _0321_ _0317_ VGND VGND VPWR VPWR top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[6\]
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_43_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1986_ _1231_ _1258_ net59 VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_35_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2607_ _0254_ _0566_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__nor2_1
X_2538_ net23 _0401_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__nor2_1
X_2469_ net189 _0199_ _0491_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1840_ net119 _0684_ _1073_ _1112_ net72 VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_69_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1771_ net117 net79 net74 VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__and3_1
X_2323_ _0352_ _0354_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__nor2_1
X_2254_ _1255_ _0307_ _0228_ _0304_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_47_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2185_ _1071_ _0225_ _0238_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1969_ net48 _1025_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold4 top8227.freeCarry VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1823_ top8227.branchForward _1034_ _1095_ _1031_ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1685_ net90 net76 net37 _0827_ _0889_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__a32o_1
X_1754_ _0689_ _0786_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_68_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ _0735_ _0337_ _0336_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2237_ _0289_ _0291_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2168_ _0220_ _0221_ _0222_ _1127_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2099_ top8227.PSRCurrentValue\[3\] _1132_ _1133_ net4 _0153_ VGND VGND VPWR VPWR
+ _0154_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1470_ net89 net75 VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2022_ top8227.internalDataflow.addressLowBusModule.busInputs\[22\] _1129_ _1294_
+ VGND VGND VPWR VPWR _1295_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2786_ clknet_4_6_0_clk _0092_ net136 VGND VGND VPWR VPWR gpio[1] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_25_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1806_ _0769_ _0795_ _0797_ _1078_ net108 VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__o41a_1
XPHY_EDGE_ROW_17_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1599_ net81 _0766_ net39 VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1668_ _0694_ net35 _0875_ _0908_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1737_ net118 _0775_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_62_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2640_ _0118_ _0567_ _0608_ _0609_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__o2bb2a_1
X_2571_ top8227.demux.state_machine.timeState\[5\] _0739_ _0758_ net71 VGND VGND VPWR
+ VPWR _0554_ sky130_fd_sc_hd__a211o_1
XFILLER_0_22_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1522_ net116 net49 _0820_ net110 VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__a22o_1
X_1453_ _0687_ net77 net74 net79 net108 VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__o311a_1
X_2005_ _1217_ _1259_ _1275_ VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__nor3_1
X_1384_ _0658_ _0683_ _0673_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2769_ clknet_4_7_0_clk _0075_ net138 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2554_ _0362_ _0363_ _0385_ _0545_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__o31a_1
XFILLER_0_42_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2623_ top8227.internalDataflow.addressLowBusModule.busInputs\[26\] _0576_ _0595_
+ _0270_ _0594_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1505_ net126 net112 VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__nor2_2
X_1436_ _0734_ _0736_ _0724_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__o21a_1
X_2485_ net178 _1303_ _0494_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_34_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1367_ top8227.demux.state_machine.currentInstruction\[5\] top8227.demux.state_machine.currentInstruction\[4\]
+ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__or2_4
XPHY_EDGE_ROW_43_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Left_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2270_ _0268_ _0319_ _0320_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_35_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1985_ net123 top8227.demux.state_machine.timeState\[1\] net65 VGND VGND VPWR VPWR
+ _1258_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2537_ _0409_ _0525_ _0530_ _0531_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__o31a_1
XFILLER_0_2_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2606_ _0178_ _0273_ _0566_ _0579_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2399_ _0175_ _0170_ net45 VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__mux2_1
X_2468_ net191 _0225_ _0491_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__mux2_1
X_1419_ net100 net103 net94 net97 VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1770_ net120 net89 net76 _0665_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__a31o_1
XFILLER_0_69_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2322_ net124 net90 _0656_ net60 _0353_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__a41o_1
X_2184_ _0238_ _0225_ net28 VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__and3b_1
X_2253_ _1308_ _1329_ _0136_ _0159_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1968_ net48 _1025_ VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1899_ net53 _1158_ _1166_ _1170_ _1148_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold5 top8227.negEdgeDetector.q1 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1822_ net123 net86 net84 VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__and3_1
X_1753_ net123 net86 net81 net72 VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__a31o_1
XFILLER_0_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1684_ net85 _0755_ net36 _0881_ _0904_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__a32o_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2167_ top8227.PSRCurrentValue\[0\] _1132_ _1133_ net1 VGND VGND VPWR VPWR _0222_
+ sky130_fd_sc_hd__a22oi_1
X_2305_ _0732_ _0733_ _1273_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__a21oi_1
X_2236_ _1292_ _0290_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2098_ top8227.internalDataflow.addressHighBusModule.busInputs\[19\] _1120_ _1130_
+ top8227.internalDataflow.accRegToDB\[3\] _1122_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2021_ top8227.PSRCurrentValue\[6\] _1132_ _1133_ net7 _1293_ VGND VGND VPWR VPWR
+ _1294_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_8_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2785_ clknet_4_6_0_clk _0091_ net136 VGND VGND VPWR VPWR gpio[0] sky130_fd_sc_hd__dfrtp_4
X_1736_ top8227.pulse_slower.currentEnableState\[1\] net157 VGND VGND VPWR VPWR top8227.pulse_slower.nextEnableState\[1\]
+ sky130_fd_sc_hd__and2b_1
X_1805_ _0657_ net79 _0695_ net83 VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__a22o_1
X_1598_ net51 _0877_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1667_ net6 _0850_ _0853_ _0945_ _0946_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__a311o_1
X_2219_ _1071_ _0225_ _0272_ _0270_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2570_ _0808_ _0499_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1521_ top8227.demux.state_machine.timeState\[1\] net49 _0820_ net107 VGND VGND VPWR
+ VPWR _0014_ sky130_fd_sc_hd__a22o_1
X_1452_ net110 _0751_ _0752_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__a21o_1
X_1383_ _0658_ _0673_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__nor2_1
X_2004_ _1217_ _1275_ _1268_ _1259_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__o211a_2
XFILLER_0_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2768_ clknet_4_12_0_clk _0074_ net143 VGND VGND VPWR VPWR gpio[15] sky130_fd_sc_hd__dfrtp_4
X_1719_ _0791_ net36 net21 _0878_ _0944_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__a221o_1
X_2699_ clknet_4_8_0_clk _0014_ net141 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2553_ net19 _0386_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__nor2_1
X_1504_ top8227.instructionLoader.interruptInjector.resetDetected gpio[21] VGND VGND
+ VPWR VPWR _0804_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_30_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2622_ _0276_ _0589_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1435_ _0643_ _0735_ net105 VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__o21bai_1
X_2484_ net165 _1327_ _0494_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__mux2_1
X_1366_ top8227.demux.state_machine.currentInstruction\[5\] top8227.demux.state_machine.currentInstruction\[4\]
+ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_21_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1984_ _1253_ _1256_ _1254_ VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2536_ top8227.internalDataflow.addressLowBusModule.busInputs\[20\] net20 VGND VGND
+ VPWR VPWR _0531_ sky130_fd_sc_hd__or2_1
X_2467_ _1153_ _1154_ _0490_ net60 VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__o31a_4
XFILLER_0_23_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2605_ _0200_ _0209_ _0655_ _0696_ _1240_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__a2111o_1
X_2398_ _0405_ _0415_ _0427_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__o21ba_1
X_1349_ top8227.demux.state_machine.currentAddress\[2\] top8227.demux.state_machine.currentAddress\[9\]
+ _0650_ top8227.demux.isAddressing VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__or4b_1
XFILLER_0_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1418_ _0657_ _0717_ _0718_ net83 VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__o31a_1
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2321_ _0803_ _0824_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__nor2_1
X_2183_ _1246_ _0230_ _0231_ _0237_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__o31a_1
X_2252_ _0201_ _0298_ _0305_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1898_ _1166_ _1170_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__nand2_1
X_1967_ net117 net57 VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__nand2_2
X_2519_ _0377_ _0378_ _0380_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__nor3_1
XFILLER_0_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold6 top8227.instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ
+ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1821_ _1093_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__inv_2
X_1752_ net123 _0724_ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__nand2_2
XFILLER_0_37_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1683_ _0769_ net37 _0863_ _0883_ _0961_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2304_ _0724_ _1037_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2097_ _1144_ _0150_ _0151_ _1142_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__o22ai_1
X_2166_ top8227.internalDataflow.addressHighBusModule.busInputs\[16\] _1120_ _1130_
+ top8227.internalDataflow.accRegToDB\[0\] _1122_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_0_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2235_ _1312_ _0284_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__and2b_1
XFILLER_0_63_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2020_ top8227.internalDataflow.addressHighBusModule.busInputs\[22\] _1120_ _1130_
+ top8227.internalDataflow.accRegToDB\[6\] _1122_ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2784_ clknet_4_6_0_clk _0090_ net135 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1804_ net59 _1076_ VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__nand2_2
XFILLER_0_40_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1735_ _1005_ _1007_ _1009_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1666_ _0657_ net85 net35 _0942_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__a31o_1
X_1597_ net146 _0876_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__nand2_1
X_2149_ top8227.demux.reset _0647_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__nand2_1
X_2218_ _0272_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1520_ net71 _0819_ net44 net51 VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__a211oi_4
XTAP_TAPCELL_ROW_10_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1451_ net110 net79 net74 VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__and3_1
X_1382_ _0673_ _0683_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__nor2_2
X_2003_ _1217_ _1275_ _1268_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2767_ clknet_4_13_0_clk _0073_ net145 VGND VGND VPWR VPWR gpio[14] sky130_fd_sc_hd__dfrtp_4
X_2698_ clknet_4_15_0_clk _0013_ net145 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_1649_ _0927_ _0928_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__or2_1
X_1718_ _0962_ _0977_ _0980_ _0985_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__or4_1
XFILLER_0_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2552_ top8227.internalDataflow.addressLowBusModule.busInputs\[22\] net20 _0538_
+ _0544_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__o211a_1
X_1503_ top8227.instructionLoader.interruptInjector.resetDetected gpio[21] VGND VGND
+ VPWR VPWR _0803_ sky130_fd_sc_hd__nor2_4
X_2483_ net169 _0133_ _0494_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__mux2_1
X_2621_ _0270_ _0593_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1434_ top8227.branchBackward top8227.branchForward VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__or2_2
X_1365_ top8227.demux.state_machine.currentInstruction\[4\] net86 VGND VGND VPWR VPWR
+ _0667_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_38_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2604_ net32 _0277_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__nand2_1
X_1983_ _1011_ _1014_ net57 VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__o21ai_4
X_2535_ net22 _0529_ _0527_ net47 VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2466_ net120 _0779_ _1031_ _0748_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__a211o_1
XFILLER_0_23_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1417_ net103 net94 net97 net100 VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2397_ _0415_ _0416_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__and2_1
X_1348_ top8227.demux.state_machine.currentAddress\[2\] top8227.demux.state_machine.currentAddress\[9\]
+ _0650_ top8227.demux.isAddressing VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout140 net9 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2320_ net70 net53 _0351_ _0348_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__a31o_1
X_2251_ _0645_ _0304_ _0298_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2182_ _1245_ _0235_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__or2_1
Xclkbuf_4_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1966_ _1238_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1897_ _1147_ _1169_ net59 VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2449_ _0467_ _0465_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__and2b_1
X_2518_ _0185_ _0514_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_Left_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold7 _0328_ VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1820_ net123 _0659_ net66 net114 VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_52_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1751_ net53 _1023_ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__and2_2
XFILLER_0_37_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1682_ _0783_ net39 _0871_ _0917_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2303_ net67 _0333_ _0334_ net55 VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_74 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2234_ _0284_ _0285_ _0288_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__a21o_1
X_2096_ top8227.internalDataflow.addressHighBusModule.busInputs\[19\] _1227_ _1228_
+ net4 _1234_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_48_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2165_ top8227.internalDataflow.addressLowBusModule.busInputs\[16\] _1129_ VGND VGND
+ VPWR VPWR _0220_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1949_ net71 _1031_ _1123_ _1221_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2783_ clknet_4_6_0_clk _0089_ net135 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1803_ _1074_ _1075_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1596_ net7 net61 net147 VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__and3b_1
X_1665_ _0659_ net36 _0889_ _0904_ _0944_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1734_ _0923_ _0935_ _0959_ _1008_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2217_ _0690_ _0694_ _0774_ net57 net118 VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__o311a_2
XFILLER_0_48_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2148_ _1256_ _1253_ _0201_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__mux2_1
X_2079_ net28 _0133_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1450_ _0673_ _0688_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__nor2_2
X_1381_ net98 net95 net92 net102 VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__or4bb_2
XTAP_TAPCELL_ROW_61_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2002_ _1195_ _1211_ _1274_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__nor3b_1
X_2766_ clknet_4_13_0_clk _0072_ net143 VGND VGND VPWR VPWR gpio[13] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_60_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2697_ clknet_4_14_0_clk _0003_ net145 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_1579_ net51 _0829_ _0851_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__nor3_1
X_1648_ net65 net36 _0866_ _0893_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__a22o_1
X_1717_ _0942_ _0957_ _0958_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2620_ _0591_ _0592_ net32 _0276_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_15_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2551_ net47 _0543_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__nand2_1
X_1433_ net111 _0732_ _0733_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__and3_1
X_2482_ net184 _0157_ _0494_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__mux2_1
X_1502_ _0801_ _0802_ net60 VGND VGND VPWR VPWR gpio[21] sky130_fd_sc_hd__o21a_4
XFILLER_0_10_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1364_ net97 net94 net103 net100 VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__and4b_1
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2749_ clknet_4_5_0_clk _0055_ net134 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1982_ _1254_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2534_ _0401_ _0528_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__nor2_1
X_2603_ _0261_ _0280_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__nor2_1
X_2396_ top8227.internalDataflow.addressHighBusModule.busInputs\[18\] net20 VGND VGND
+ VPWR VPWR _0426_ sky130_fd_sc_hd__or2_1
X_1347_ top8227.demux.state_machine.currentAddress\[8\] top8227.demux.state_machine.currentAddress\[0\]
+ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__or2_1
X_2465_ top8227.internalDataflow.addressHighBusModule.busInputs\[23\] net20 _0483_
+ _0356_ _0489_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__o221a_1
X_1416_ net103 net97 net94 net100 VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout141 net142 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_4
Xfanout130 net140 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2250_ _0745_ _0746_ _0303_ net58 VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__o31a_1
XFILLER_0_20_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2181_ _0235_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1965_ _1071_ _1237_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2517_ _0508_ _0509_ _0208_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__mux2_1
X_1896_ _1010_ _1111_ _1168_ _1167_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__or4b_1
X_2379_ top8227.internalDataflow.addressHighBusModule.busInputs\[16\] net24 _0387_
+ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__a21oi_1
X_2448_ _0471_ _0473_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold8 _0033_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dlygate4sd3_1
X_1750_ top8227.demux.state_machine.currentAddress\[12\] _0809_ _1019_ _1022_ VGND
+ VGND VPWR VPWR _1023_ sky130_fd_sc_hd__a211o_1
X_1681_ _0957_ _0959_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__or2_1
X_2164_ _1142_ _0218_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__nor2_1
X_2302_ _0760_ _1034_ _1140_ _1221_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__or4_1
XFILLER_0_29_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2233_ _0283_ _0287_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2095_ _1183_ _0149_ _1185_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_0_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1948_ top8227.demux.state_machine.timeState\[1\] _0740_ _1220_ VGND VGND VPWR VPWR
+ _1221_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_31_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1879_ net107 net66 net64 net116 VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2782_ clknet_4_5_0_clk _0088_ net135 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1802_ _0694_ _0724_ _0792_ net119 VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__o31a_1
X_1733_ _0933_ _0945_ _0968_ _0972_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_13_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1595_ _0840_ _0845_ _0874_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__a21o_2
XFILLER_0_40_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1664_ _0778_ net36 _0889_ _0943_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2147_ _0201_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2216_ net48 _0245_ _0269_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__or3_2
X_2078_ net31 _0126_ _0132_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_8_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1380_ net100 net97 top8227.demux.state_machine.currentInstruction\[3\] net103 VGND
+ VGND VPWR VPWR _0682_ sky130_fd_sc_hd__and4bb_2
X_2001_ _0734_ _1273_ _1213_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_61_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2765_ clknet_4_13_0_clk _0071_ net143 VGND VGND VPWR VPWR gpio[12] sky130_fd_sc_hd__dfrtp_4
X_2696_ clknet_4_15_0_clk _0002_ net143 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1716_ net29 _0836_ _0887_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1578_ top8227.demux.state_machine.currentAddress\[0\] net41 _0863_ VGND VGND VPWR
+ VPWR _0864_ sky130_fd_sc_hd__a21o_1
X_1647_ _0781_ net36 _0926_ net44 VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2550_ _0540_ _0541_ _0542_ _0358_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2481_ net173 _0177_ _0494_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__mux2_1
X_1501_ _0737_ _0764_ _0773_ _0798_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1432_ _0726_ _0728_ _0729_ _0731_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__and4_2
X_1363_ _0641_ net109 net88 _0656_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_38_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2679_ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] _0648_ _1242_
+ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__or3_1
X_2748_ clknet_4_5_0_clk _0054_ net134 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1981_ _1128_ _1135_ _1193_ _1092_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__o22a_1
XFILLER_0_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2533_ _0163_ _0400_ _0140_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2602_ _0562_ _0571_ _0576_ net201 VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__a22o_1
X_2395_ _0423_ _0424_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__nor2_1
X_2464_ _0485_ _0487_ _0488_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1346_ gpio[16] VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.nmiSync.in
+ sky130_fd_sc_hd__inv_2
X_1415_ net69 net56 VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout120 net122 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_2
Xfanout131 net132 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout142 net9 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__buf_2
XFILLER_0_56_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2180_ _1279_ _0234_ _0233_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__o21a_2
XFILLER_0_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_25_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1964_ net30 _1236_ _1137_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_43_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1895_ _0742_ _0778_ _0782_ _0793_ net121 VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__o41a_1
X_2447_ _0460_ _0472_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__nand2_1
X_2516_ top8227.internalDataflow.addressLowBusModule.busInputs\[17\] _0409_ _0511_
+ net47 _0513_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2378_ net19 _0389_ _0408_ top8227.internalDataflow.addressHighBusModule.busInputs\[16\]
+ _0407_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__o221a_1
XFILLER_0_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold9 top8227.pulse_slower.currentEnableState\[0\] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2301_ top8227.demux.state_machine.currentAddress\[6\] top8227.demux.state_machine.currentAddress\[7\]
+ _1223_ _0332_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__o22a_1
X_1680_ net63 net37 _0866_ _0909_ _0958_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__a221o_1
X_2163_ _1227_ _1228_ _0216_ _0217_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__o31a_1
XFILLER_0_29_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2232_ _0120_ _0263_ _0281_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_51_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2094_ top8227.internalDataflow.addressLowBusModule.busInputs\[35\] _1188_ _0147_
+ _0148_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_16_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1947_ net105 net64 _1219_ VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1878_ net109 net89 net76 _0659_ net116 VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_8_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2781_ clknet_4_6_0_clk _0087_ net135 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1663_ net39 _0877_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1801_ net119 _0697_ _1015_ _1073_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__a211o_1
X_1732_ _0940_ _0948_ _0988_ _1006_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_13_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1594_ gpio[21] _0828_ _0838_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2077_ _1127_ _0131_ net30 VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__or3b_2
X_2146_ _0191_ _0196_ _1091_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__mux2_2
X_2215_ top8227.PSRCurrentValue\[3\] net33 _0268_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__and3_4
XFILLER_0_48_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2000_ net105 _0808_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_61_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2764_ clknet_4_13_0_clk _0070_ net143 VGND VGND VPWR VPWR gpio[11] sky130_fd_sc_hd__dfrtp_4
X_2695_ clknet_4_14_0_clk _0001_ net144 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1646_ net56 _0881_ _0887_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__and3_1
X_1715_ _0941_ _0982_ _0990_ _0991_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__or4_1
XFILLER_0_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1577_ _0803_ _0861_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__nor2_4
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2129_ top8227.internalDataflow.addressLowBusModule.busInputs\[34\] _1277_ _1282_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[18\] _0183_ VGND VGND VPWR
+ VPWR _0184_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2480_ net163 _0199_ _0494_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__mux2_1
X_1500_ _0777_ _0799_ _0800_ net109 VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__o31a_1
XFILLER_0_2_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1431_ _0645_ _0723_ _0725_ _0727_ _0730_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__a2111oi_4
X_1362_ _0641_ net88 _0656_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_38_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2747_ clknet_4_5_0_clk _0053_ net134 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_1629_ net44 _0908_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__and2_1
X_2678_ net164 _1237_ _0637_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1980_ _1024_ _1252_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__nand2_2
X_2532_ _0140_ _0391_ _0526_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__a21bo_1
X_2463_ _0485_ _0487_ net46 VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_23_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2601_ _1034_ _0575_ _1024_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__o21ai_4
X_2394_ _0420_ _0421_ _0422_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__nor3_1
XFILLER_0_64_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1414_ gpio[19] _0711_ top8227.pulse_slower.nextEnableState\[0\] net69 VGND VGND
+ VPWR VPWR _0715_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1345_ gpio[17] VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.interruptRequest
+ sky130_fd_sc_hd__inv_2
XFILLER_0_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout143 net145 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_4
Xfanout121 net122 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_4
Xfanout132 net133 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_4
Xfanout110 top8227.demux.state_machine.timeState\[4\] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_69_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1963_ _1144_ _1193_ _1235_ _1142_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1894_ net117 _0794_ _1062_ VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__a21oi_1
X_2446_ _0459_ _0461_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__nand2b_1
X_2515_ top8227.internalDataflow.addressLowBusModule.busInputs\[16\] _0379_ _0512_
+ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2377_ net20 VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2300_ net125 net113 net81 net75 VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__and4b_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2231_ _0284_ _0285_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__nand2_1
X_2162_ top8227.internalDataflow.addressHighBusModule.busInputs\[16\] _1227_ _1228_
+ net1 VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__a22oi_1
X_2093_ top8227.internalDataflow.stackBusModule.busInputs\[43\] _1186_ _1187_ top8227.internalDataflow.accRegToDB\[3\]
+ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1946_ top8227.demux.state_machine.timeState\[5\] net87 net83 VGND VGND VPWR VPWR
+ _1219_ sky130_fd_sc_hd__and3_1
X_1877_ _1079_ _1080_ _1149_ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__or3_1
X_2429_ _0453_ _0455_ net47 VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_66_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1800_ net116 net88 net76 VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__and3_1
X_2780_ clknet_4_5_0_clk _0086_ net134 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1731_ _0973_ _0975_ _0978_ _0984_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1662_ _0685_ net34 _0875_ _0883_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__a22o_1
X_1593_ net186 net41 _0870_ _0873_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2214_ top8227.PSRCurrentValue\[3\] net33 VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_64_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2076_ top8227.internalDataflow.addressLowBusModule.busInputs\[20\] _1129_ _0127_
+ _0130_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__a211oi_1
X_2145_ net28 _0199_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__nand2_2
X_1929_ top8227.demux.state_machine.timeState\[5\] net63 _1201_ net64 net71 VGND VGND
+ VPWR VPWR _1202_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2763_ clknet_4_13_0_clk _0069_ net143 VGND VGND VPWR VPWR gpio[10] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_61_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2694_ clknet_4_15_0_clk _0012_ net144 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1576_ _0861_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__inv_2
X_1645_ _0900_ _0906_ _0921_ _0924_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__or4_1
XFILLER_0_13_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1714_ _0910_ _0952_ _0985_ _0986_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2128_ net3 _1272_ _1276_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__and3_1
X_2059_ top8227.internalDataflow.addressLowBusModule.busInputs\[37\] _1277_ _1282_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[21\] VGND VGND VPWR VPWR
+ _1332_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_24_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1430_ top8227.PSRCurrentValue\[6\] _0669_ net75 VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__or3b_1
XFILLER_0_37_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1361_ _0655_ _0662_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__nor2_1
X_2746_ clknet_4_5_0_clk _0052_ net134 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1559_ net4 net62 _0832_ net148 VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__and4b_1
XFILLER_0_41_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1628_ net147 net54 _0826_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__and3b_2
X_2677_ net185 _1303_ _0637_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2600_ _1033_ _0574_ _1025_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__or3b_1
XFILLER_0_2_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2393_ _0421_ _0422_ _0420_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__o21a_1
X_2531_ _0140_ _0391_ net22 VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__o21a_1
X_2462_ _1193_ _0396_ _0486_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__o21ai_2
X_1413_ _0653_ _0712_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1344_ top8227.instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning VGND
+ VGND VPWR VPWR _0649_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2729_ clknet_4_2_0_clk _0035_ net131 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout144 net145 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_4
Xfanout122 top8227.demux.state_machine.timeState\[0\] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout111 net112 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_2
Xfanout133 net140 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__buf_2
Xfanout100 net101 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_57_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1962_ top8227.internalDataflow.addressHighBusModule.busInputs\[23\] _1227_ _1228_
+ net146 _1234_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_34_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1893_ _0653_ _0712_ _1162_ _1165_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__or4_2
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2445_ top8227.internalDataflow.addressHighBusModule.busInputs\[22\] net25 VGND VGND
+ VPWR VPWR _0471_ sky130_fd_sc_hd__xor2_1
X_2514_ net19 _0380_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__nor2_1
X_2376_ net46 _0352_ _0354_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__or3_2
XFILLER_0_19_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2230_ _1314_ _0118_ _0283_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__nand3_1
X_2161_ net48 _1233_ _1229_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2092_ top8227.internalDataflow.stackBusModule.busInputs\[35\] _1182_ _1189_ top8227.internalDataflow.addressLowBusModule.busInputs\[27\]
+ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1945_ _1212_ _1214_ _1217_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1876_ net108 _0684_ _0754_ VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__a21o_1
X_2428_ _0455_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__inv_2
X_2359_ _0164_ _0390_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1592_ _0871_ _0872_ _0804_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__o21a_1
X_1730_ _0912_ _1000_ _1001_ _1004_ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1661_ _0934_ _0936_ _0939_ _0940_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__or4_1
X_2144_ net31 _0198_ _0192_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__o21ai_4
XPHY_EDGE_ROW_37_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2213_ net48 _0245_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_64_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2075_ net148 _1133_ _0129_ _1132_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1859_ _1098_ _1119_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__nor2_2
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1928_ top8227.demux.state_machine.timeState\[1\] top8227.demux.state_machine.timeState\[5\]
+ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_55_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_64_Left_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2762_ clknet_4_15_0_clk _0068_ net143 VGND VGND VPWR VPWR gpio[9] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1713_ _0886_ _0960_ _0989_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2693_ clknet_4_14_0_clk _0011_ net144 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1575_ _0829_ _0859_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1644_ _0697_ net35 _0875_ _0922_ _0923_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2127_ _1256_ _0180_ _0181_ _1245_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2058_ _1245_ _1330_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_24_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1360_ net99 net104 net93 net96 VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__or4b_2
XFILLER_0_58_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2745_ clknet_4_5_0_clk _0051_ net135 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_2676_ net182 _1327_ _0637_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__mux2_1
X_2814_ clknet_4_1_0_clk VGND VGND VPWR VPWR gpio[23] sky130_fd_sc_hd__buf_2
X_1558_ net54 net21 _0841_ _0847_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__a31o_1
X_1627_ _0701_ net29 VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__nor2_1
X_1489_ net89 _0702_ _0766_ net82 VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2530_ _0371_ _0372_ _0382_ _0524_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__o31a_1
X_2392_ _0387_ _0411_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__and2_1
X_2461_ _1235_ _1137_ net45 VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__mux2_1
X_1343_ net146 VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__inv_2
X_1412_ _0653_ _0712_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2728_ clknet_4_3_0_clk _0034_ net131 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2659_ top8227.internalDataflow.addressLowBusModule.busInputs\[30\] _0576_ _0622_
+ _0627_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__a22o_1
Xfanout123 top8227.demux.state_machine.timeState\[0\] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_4
Xfanout145 net9 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__buf_2
Xfanout134 net135 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_4
Xfanout112 top8227.demux.state_machine.timeState\[4\] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_4
Xfanout101 top8227.demux.state_machine.currentInstruction\[1\] VGND VGND VPWR VPWR
+ net101 sky130_fd_sc_hd__buf_2
XFILLER_0_69_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1961_ _1227_ _1228_ _1229_ _1233_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__nor4b_4
X_1892_ net127 _1163_ _1164_ net72 VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_7_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2513_ _0207_ _0510_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__xnor2_1
X_2375_ net46 _0406_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__nand2_1
X_2444_ top8227.internalDataflow.addressHighBusModule.busInputs\[21\] _0408_ _0463_
+ net19 _0470_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__o221a_1
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_48 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2160_ _1144_ _0214_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2091_ _0143_ _0144_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__or2_1
X_1944_ _0653_ _0712_ _1216_ VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__or3_2
X_1875_ net59 _1147_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2427_ _0124_ _0395_ _0454_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_24_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_15_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
X_2358_ _0185_ _0208_ _0235_ _0354_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__and4b_1
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2289_ net111 _0698_ _1230_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1591_ net146 net7 _0865_ _0848_ _0839_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__a32o_1
XFILLER_0_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1660_ net6 _0826_ _0875_ _0690_ net34 VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__a32o_1
X_2143_ _1143_ _0196_ _0197_ _1142_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__o2bb2a_1
X_2212_ _1290_ _0266_ _0265_ _1292_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_64_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2074_ net114 _0647_ net66 _0128_ _1230_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__a41o_1
X_1858_ top8227.internalDataflow.addressHighBusModule.busInputs\[23\] _1120_ _1130_
+ top8227.internalDataflow.accRegToDB\[7\] _1122_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__a221o_1
X_1927_ _0771_ net73 _1199_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1789_ net117 net83 net74 VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_27_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2761_ clknet_4_13_0_clk _0067_ net143 VGND VGND VPWR VPWR gpio[8] sky130_fd_sc_hd__dfrtp_4
X_2692_ clknet_4_14_0_clk _0010_ net144 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_1 _0648_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1712_ _0906_ _0963_ _0987_ _0988_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1643_ net91 _0695_ net34 net21 _0922_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__a32o_1
X_1574_ _0859_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2057_ _1256_ _1253_ _1329_ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__mux2_1
X_2126_ _1253_ _0179_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_16_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2813_ clknet_4_3_0_clk _0117_ net131 VGND VGND VPWR VPWR top8227.PSRCurrentValue\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_21_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2744_ clknet_4_9_0_clk _0050_ net139 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_2675_ net171 _0133_ _0637_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__mux2_1
X_1626_ _0901_ _0902_ _0905_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1557_ net50 _0831_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1488_ _0655_ _0703_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__nor2_1
X_2109_ _0163_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_37_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2460_ _0475_ _0478_ _0484_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__a21oi_1
X_2391_ top8227.internalDataflow.addressHighBusModule.busInputs\[17\] top8227.internalDataflow.addressHighBusModule.busInputs\[16\]
+ net25 VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1411_ net69 _0711_ gpio[19] VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__a21oi_4
X_1342_ top8227.demux.nmi VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout113 top8227.demux.state_machine.timeState\[4\] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_1
X_1609_ _0831_ _0859_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__nor2_2
X_2589_ net58 _1064_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__nand2_1
X_2727_ clknet_4_2_0_clk net150 net133 VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.nmiGeneratedFF.synchronizedNMI
+ sky130_fd_sc_hd__dfrtp_1
X_2658_ _0292_ _0293_ _0626_ _0623_ _0271_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__a311o_1
Xfanout102 net104 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__buf_2
XFILLER_0_14_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout124 top8227.demux.state_machine.timeState\[0\] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
Xfanout146 net8 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_4
Xfanout135 net140 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_19_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1960_ _1231_ _1232_ _1085_ VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__and3b_1
X_1891_ _0750_ _0769_ _0779_ net121 VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__o31a_1
XFILLER_0_28_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2443_ _0465_ _0466_ _0467_ _0469_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__a31o_1
XFILLER_0_59_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2512_ _0508_ _0509_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2374_ _0399_ _0404_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_19_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2090_ _0143_ _0144_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1943_ net67 _1215_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1874_ _1146_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2426_ _0125_ _0132_ net45 VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__mux2_1
X_2357_ _0387_ _0388_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_67_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2288_ top8227.instructionLoader.interruptInjector.irqGenerated _0311_ net155 VGND
+ VGND VPWR VPWR _0033_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1590_ net54 _0828_ _0869_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2142_ top8227.internalDataflow.addressHighBusModule.busInputs\[17\] _1227_ _1228_
+ net2 _1234_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__a221oi_4
X_2073_ top8227.demux.reset top8227.demux.setInterruptFlag VGND VGND VPWR VPWR _0128_
+ sky130_fd_sc_hd__nor2_1
X_2211_ _1289_ _1312_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1857_ net50 _1104_ _1118_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__nor3_2
X_1926_ _0687_ _0743_ net90 _0671_ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1788_ _1012_ _1060_ _1025_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__or3b_1
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2409_ _0427_ _0430_ _0436_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_27_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_14_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
X_2691_ clknet_4_14_0_clk _0009_ net144 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_2 _0720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1642_ net52 _0903_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__nor2_1
X_1711_ _0689_ net35 _0875_ _0897_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2760_ clknet_4_9_0_clk _0066_ net141 VGND VGND VPWR VPWR top8227.demux.reset sky130_fd_sc_hd__dfrtp_4
XFILLER_0_67_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1573_ net148 _0839_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__nand2b_1
X_2056_ _1318_ _1325_ _1092_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__mux2_1
X_2125_ _0179_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1909_ _1171_ _1179_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__nor2_2
XFILLER_0_29_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2812_ clknet_4_15_0_clk _0116_ net145 VGND VGND VPWR VPWR top8227.demux.isAddressing
+ sky130_fd_sc_hd__dfstp_1
X_2743_ clknet_4_12_0_clk _0049_ net139 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_46_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1556_ _0842_ _0846_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2674_ net181 _0157_ _0637_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__mux2_1
X_1625_ net66 net36 _0866_ _0904_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__a22o_1
X_1487_ _0698_ _0787_ net107 VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__o21a_1
XFILLER_0_68_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2108_ _1280_ _0162_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_37_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2039_ _1311_ _1304_ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1410_ net69 _0711_ VGND VGND VPWR VPWR gpio[22] sky130_fd_sc_hd__nand2_4
X_2390_ top8227.internalDataflow.addressHighBusModule.busInputs\[18\] net25 VGND VGND
+ VPWR VPWR _0420_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1341_ top8227.PSRCurrentValue\[6\] VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2726_ clknet_4_2_0_clk top8227.instructionLoader.interruptInjector.nmiSync.in net132
+ VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.nmiSync.nextQ2 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout136 net137 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_4
X_1539_ net3 net61 VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__nand2_1
Xfanout125 net127 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
X_1608_ _0780_ net39 _0863_ _0887_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__a22o_1
Xfanout147 net6 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_4
Xfanout114 top8227.demux.state_machine.timeState\[2\] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2657_ _0586_ _0625_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__xnor2_1
Xfanout103 net104 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_2
X_2588_ net58 _1064_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_48_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1890_ net80 _0695_ _0780_ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2373_ _0393_ _0399_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__or2_1
X_2442_ net46 _0468_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__nand2_1
X_2511_ _0235_ _0354_ net22 VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2709_ clknet_4_11_0_clk _0023_ net142 VGND VGND VPWR VPWR top8227.demux.state_machine.currentInstruction\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1942_ top8227.demux.state_machine.currentAddress\[6\] top8227.demux.state_machine.currentAddress\[7\]
+ _0811_ _1019_ net124 VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__o32a_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1873_ _1043_ _1145_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2356_ _0359_ _0360_ _0386_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__nor3_1
X_2425_ _0427_ _0430_ _0441_ _0452_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__a31o_1
XFILLER_0_66_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2287_ net154 _0324_ top8227.instructionLoader.interruptInjector.irqGenerated VGND
+ VGND VPWR VPWR _0328_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2210_ _0118_ _0264_ _1314_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_64_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2072_ top8227.internalDataflow.addressHighBusModule.busInputs\[20\] _1120_ _1130_
+ top8227.internalDataflow.accRegToDB\[4\] _1122_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__a221o_1
X_2141_ _0193_ _0194_ _0195_ _1185_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__o31a_1
XFILLER_0_71_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1925_ _0671_ _0686_ _0752_ _1196_ _1197_ VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_71_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1856_ _1106_ _1117_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__nor2_2
XFILLER_0_12_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1787_ net118 _1039_ _1059_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__a21o_1
X_2408_ _0403_ _0415_ _0430_ _0399_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__nand4b_1
X_2339_ _0369_ _0370_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_33_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold50 top8227.internalDataflow.addressLowBusModule.busInputs\[35\] VGND VGND VPWR
+ VPWR net198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1572_ top8227.demux.state_machine.currentAddress\[1\] net42 net21 _0849_ VGND VGND
+ VPWR VPWR _0004_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2690_ clknet_4_15_0_clk _0008_ net143 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1641_ _0912_ _0916_ _0920_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__or3_1
X_1710_ _0897_ _0908_ _0850_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_3 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Left_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2124_ _1128_ _0169_ _0174_ _1092_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__o22a_2
X_2055_ net28 _1327_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__nand2_1
X_1908_ _1166_ _1178_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1839_ net107 net89 net77 VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2742_ clknet_4_12_0_clk _0048_ net139 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[22\]
+ sky130_fd_sc_hd__dfrtp_4
X_2811_ clknet_4_12_0_clk _0115_ net139 VGND VGND VPWR VPWR top8227.branchBackward
+ sky130_fd_sc_hd__dfrtp_1
X_1555_ net54 _0840_ _0845_ net42 top8227.demux.state_machine.currentAddress\[4\]
+ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__a32o_1
X_2673_ net167 _0177_ _0637_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__mux2_1
X_1624_ net36 _0903_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__nor2_1
X_2107_ net4 _1281_ _1284_ top8227.internalDataflow.addressLowBusModule.busInputs\[27\]
+ _0161_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_37_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1486_ net98 net88 _0656_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__and3_2
XFILLER_0_64_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2038_ _1245_ _1309_ _1310_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_13_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1340_ top8227.PSRCurrentValue\[1\] VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2725_ clknet_4_2_0_clk net149 net141 VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2656_ _0289_ _0624_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout137 net140 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
Xfanout148 net5 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_4
X_1538_ net2 net1 net62 VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__o21a_1
Xfanout126 net127 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
Xfanout115 top8227.demux.state_machine.timeState\[2\] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__buf_2
X_1607_ net147 _0853_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__and2b_4
X_1469_ net108 net89 _0705_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__and3_1
Xfanout104 top8227.demux.state_machine.currentInstruction\[0\] VGND VGND VPWR VPWR
+ net104 sky130_fd_sc_hd__clkbuf_2
X_2587_ net33 _0561_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2510_ _0235_ net22 VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2372_ net24 _0403_ _0393_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__o21ai_1
X_2441_ _0466_ _0467_ _0465_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2708_ clknet_4_10_0_clk _0022_ net142 VGND VGND VPWR VPWR top8227.demux.state_machine.currentInstruction\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2639_ _1304_ _0272_ _0563_ _0119_ _0567_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1941_ _0736_ _0806_ _1213_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__o21ai_1
X_1872_ _0783_ _0786_ _1084_ net123 VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__o31a_1
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2355_ _0360_ _0386_ _0359_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__o21a_1
X_2424_ _0436_ _0440_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__and2_1
X_2286_ top8227.demux.nmi _0311_ _0327_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2140_ top8227.internalDataflow.stackBusModule.busInputs\[41\] _1186_ _1189_ top8227.internalDataflow.addressLowBusModule.busInputs\[25\]
+ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2071_ _1143_ _0124_ _0125_ _1142_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_48_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1855_ _1091_ _1127_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__or2_2
X_1924_ _0750_ _0769_ net111 VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1786_ net98 net102 net83 _0692_ net121 VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_21_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2407_ _0405_ _0415_ _0430_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__nor3_1
X_2338_ top8227.internalDataflow.addressLowBusModule.busInputs\[20\] net22 VGND VGND
+ VPWR VPWR _0370_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2269_ net49 gpio[20] top8227.negEdgeDetector.q1 VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__or3b_1
XFILLER_0_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold40 top8227.internalDataflow.addressLowBusModule.busInputs\[36\] VGND VGND VPWR
+ VPWR net188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold51 top8227.demux.isAddressing VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1571_ net2 _0853_ _0857_ net41 net179 VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__a32o_1
X_1640_ _0883_ _0917_ _0919_ net54 VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__and4b_1
XANTENNA_4 dataBusIn[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2123_ net28 _0177_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__nand2_1
X_2054_ _1326_ _1325_ net30 VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__mux2_2
X_1907_ _1166_ _1178_ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_32_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1838_ net120 _0751_ _1011_ _1064_ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__a211o_1
X_1769_ _1040_ _1041_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2741_ clknet_4_12_0_clk _0047_ net138 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[21\]
+ sky130_fd_sc_hd__dfrtp_2
X_2810_ clknet_4_4_0_clk _0114_ net130 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_2672_ net166 _0199_ _0637_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1554_ gpio[21] _0828_ _0843_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__and3_1
X_1623_ net8 net147 net7 net61 VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__o31a_1
X_1485_ net90 net74 VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__and2_1
.ends

